module bp_fe_top (clk_i,
    reset_i,
    freeze_i,
    icache_id_i,
    cfg_w_v_i,
    fe_cmd_v_i,
    fe_cmd_ready_o,
    fe_queue_v_o,
    fe_queue_ready_i,
    lce_req_v_o,
    lce_req_ready_i,
    lce_resp_v_o,
    lce_resp_ready_i,
    lce_data_resp_v_o,
    lce_data_resp_ready_i,
    lce_cmd_v_i,
    lce_cmd_ready_o,
    lce_data_cmd_v_i,
    lce_data_cmd_ready_o,
    lce_data_cmd_v_o,
    lce_data_cmd_ready_i,
    cfg_addr_i,
    cfg_data_i,
    fe_cmd_i,
    fe_queue_o,
    lce_cmd_i,
    lce_data_cmd_i,
    lce_data_cmd_o,
    lce_data_resp_o,
    lce_req_o,
    lce_resp_o);
 input clk_i;
 input reset_i;
 input freeze_i;
 input icache_id_i;
 input cfg_w_v_i;
 input fe_cmd_v_i;
 output fe_cmd_ready_o;
 output fe_queue_v_o;
 input fe_queue_ready_i;
 output lce_req_v_o;
 input lce_req_ready_i;
 output lce_resp_v_o;
 input lce_resp_ready_i;
 output lce_data_resp_v_o;
 input lce_data_resp_ready_i;
 input lce_cmd_v_i;
 output lce_cmd_ready_o;
 input lce_data_cmd_v_i;
 output lce_data_cmd_ready_o;
 output lce_data_cmd_v_o;
 input lce_data_cmd_ready_i;
 input [15:0] cfg_addr_i;
 input [31:0] cfg_data_i;
 input [75:0] fe_cmd_i;
 output [99:0] fe_queue_o;
 input [52:0] lce_cmd_i;
 input [517:0] lce_data_cmd_i;
 output [517:0] lce_data_cmd_o;
 output [553:0] lce_data_resp_o;
 output [113:0] lce_req_o;
 output [42:0] lce_resp_o;

 FILLCELL_X1 PHY_1 ();
 FILLCELL_X1 PHY_10 ();
 FILLCELL_X1 PHY_100 ();
 FILLCELL_X1 PHY_1000 ();
 FILLCELL_X1 PHY_1001 ();
 FILLCELL_X1 PHY_1002 ();
 FILLCELL_X1 PHY_1003 ();
 FILLCELL_X1 PHY_1004 ();
 FILLCELL_X1 PHY_1005 ();
 FILLCELL_X1 PHY_1006 ();
 FILLCELL_X1 PHY_1007 ();
 FILLCELL_X1 PHY_1008 ();
 FILLCELL_X1 PHY_1009 ();
 FILLCELL_X1 PHY_101 ();
 FILLCELL_X1 PHY_1010 ();
 FILLCELL_X1 PHY_1011 ();
 FILLCELL_X1 PHY_1012 ();
 FILLCELL_X1 PHY_1013 ();
 FILLCELL_X1 PHY_1014 ();
 FILLCELL_X1 PHY_1015 ();
 FILLCELL_X1 PHY_1016 ();
 FILLCELL_X1 PHY_1017 ();
 FILLCELL_X1 PHY_1018 ();
 FILLCELL_X1 PHY_1019 ();
 FILLCELL_X1 PHY_102 ();
 FILLCELL_X1 PHY_1020 ();
 FILLCELL_X1 PHY_1021 ();
 FILLCELL_X1 PHY_1022 ();
 FILLCELL_X1 PHY_1023 ();
 FILLCELL_X1 PHY_1024 ();
 FILLCELL_X1 PHY_1025 ();
 FILLCELL_X1 PHY_1026 ();
 FILLCELL_X1 PHY_1027 ();
 FILLCELL_X1 PHY_1028 ();
 FILLCELL_X1 PHY_1029 ();
 FILLCELL_X1 PHY_103 ();
 FILLCELL_X1 PHY_1030 ();
 FILLCELL_X1 PHY_1031 ();
 FILLCELL_X1 PHY_1032 ();
 FILLCELL_X1 PHY_1033 ();
 FILLCELL_X1 PHY_1034 ();
 FILLCELL_X1 PHY_1035 ();
 FILLCELL_X1 PHY_1036 ();
 FILLCELL_X1 PHY_1037 ();
 FILLCELL_X1 PHY_1038 ();
 FILLCELL_X1 PHY_1039 ();
 FILLCELL_X1 PHY_104 ();
 FILLCELL_X1 PHY_1040 ();
 FILLCELL_X1 PHY_1041 ();
 FILLCELL_X1 PHY_1042 ();
 FILLCELL_X1 PHY_1043 ();
 FILLCELL_X1 PHY_1044 ();
 FILLCELL_X1 PHY_1045 ();
 FILLCELL_X1 PHY_1046 ();
 FILLCELL_X1 PHY_1047 ();
 FILLCELL_X1 PHY_1048 ();
 FILLCELL_X1 PHY_1049 ();
 FILLCELL_X1 PHY_105 ();
 FILLCELL_X1 PHY_1050 ();
 FILLCELL_X1 PHY_1051 ();
 FILLCELL_X1 PHY_1052 ();
 FILLCELL_X1 PHY_1053 ();
 FILLCELL_X1 PHY_1054 ();
 FILLCELL_X1 PHY_1055 ();
 FILLCELL_X1 PHY_1056 ();
 FILLCELL_X1 PHY_1057 ();
 FILLCELL_X1 PHY_1058 ();
 FILLCELL_X1 PHY_1059 ();
 FILLCELL_X1 PHY_106 ();
 FILLCELL_X1 PHY_1060 ();
 FILLCELL_X1 PHY_1061 ();
 FILLCELL_X1 PHY_1062 ();
 FILLCELL_X1 PHY_1063 ();
 FILLCELL_X1 PHY_1064 ();
 FILLCELL_X1 PHY_1065 ();
 FILLCELL_X1 PHY_1066 ();
 FILLCELL_X1 PHY_1067 ();
 FILLCELL_X1 PHY_1068 ();
 FILLCELL_X1 PHY_1069 ();
 FILLCELL_X1 PHY_107 ();
 FILLCELL_X1 PHY_1070 ();
 FILLCELL_X1 PHY_1071 ();
 FILLCELL_X1 PHY_1072 ();
 FILLCELL_X1 PHY_1073 ();
 FILLCELL_X1 PHY_1074 ();
 FILLCELL_X1 PHY_1075 ();
 FILLCELL_X1 PHY_1076 ();
 FILLCELL_X1 PHY_1077 ();
 FILLCELL_X1 PHY_1078 ();
 FILLCELL_X1 PHY_1079 ();
 FILLCELL_X1 PHY_108 ();
 FILLCELL_X1 PHY_1080 ();
 FILLCELL_X1 PHY_1081 ();
 FILLCELL_X1 PHY_1082 ();
 FILLCELL_X1 PHY_1083 ();
 FILLCELL_X1 PHY_1084 ();
 FILLCELL_X1 PHY_1085 ();
 FILLCELL_X1 PHY_1086 ();
 FILLCELL_X1 PHY_1087 ();
 FILLCELL_X1 PHY_1088 ();
 FILLCELL_X1 PHY_1089 ();
 FILLCELL_X1 PHY_109 ();
 FILLCELL_X1 PHY_1090 ();
 FILLCELL_X1 PHY_1091 ();
 FILLCELL_X1 PHY_1092 ();
 FILLCELL_X1 PHY_1093 ();
 FILLCELL_X1 PHY_1094 ();
 FILLCELL_X1 PHY_1095 ();
 FILLCELL_X1 PHY_1096 ();
 FILLCELL_X1 PHY_1097 ();
 FILLCELL_X1 PHY_1098 ();
 FILLCELL_X1 PHY_1099 ();
 FILLCELL_X1 PHY_11 ();
 FILLCELL_X1 PHY_110 ();
 FILLCELL_X1 PHY_1100 ();
 FILLCELL_X1 PHY_1101 ();
 FILLCELL_X1 PHY_1102 ();
 FILLCELL_X1 PHY_1103 ();
 FILLCELL_X1 PHY_1104 ();
 FILLCELL_X1 PHY_1105 ();
 FILLCELL_X1 PHY_1106 ();
 FILLCELL_X1 PHY_1107 ();
 FILLCELL_X1 PHY_1108 ();
 FILLCELL_X1 PHY_1109 ();
 FILLCELL_X1 PHY_111 ();
 FILLCELL_X1 PHY_1110 ();
 FILLCELL_X1 PHY_1111 ();
 FILLCELL_X1 PHY_1112 ();
 FILLCELL_X1 PHY_1113 ();
 FILLCELL_X1 PHY_1114 ();
 FILLCELL_X1 PHY_1115 ();
 FILLCELL_X1 PHY_1116 ();
 FILLCELL_X1 PHY_1117 ();
 FILLCELL_X1 PHY_1118 ();
 FILLCELL_X1 PHY_1119 ();
 FILLCELL_X1 PHY_112 ();
 FILLCELL_X1 PHY_1120 ();
 FILLCELL_X1 PHY_1121 ();
 FILLCELL_X1 PHY_1122 ();
 FILLCELL_X1 PHY_1123 ();
 FILLCELL_X1 PHY_1124 ();
 FILLCELL_X1 PHY_1125 ();
 FILLCELL_X1 PHY_1126 ();
 FILLCELL_X1 PHY_1127 ();
 FILLCELL_X1 PHY_1128 ();
 FILLCELL_X1 PHY_1129 ();
 FILLCELL_X1 PHY_113 ();
 FILLCELL_X1 PHY_1130 ();
 FILLCELL_X1 PHY_1131 ();
 FILLCELL_X1 PHY_1132 ();
 FILLCELL_X1 PHY_1133 ();
 FILLCELL_X1 PHY_1134 ();
 FILLCELL_X1 PHY_1135 ();
 FILLCELL_X1 PHY_1136 ();
 FILLCELL_X1 PHY_1137 ();
 FILLCELL_X1 PHY_1138 ();
 FILLCELL_X1 PHY_1139 ();
 FILLCELL_X1 PHY_114 ();
 FILLCELL_X1 PHY_1140 ();
 FILLCELL_X1 PHY_1141 ();
 FILLCELL_X1 PHY_1142 ();
 FILLCELL_X1 PHY_1143 ();
 FILLCELL_X1 PHY_1144 ();
 FILLCELL_X1 PHY_1145 ();
 FILLCELL_X1 PHY_1146 ();
 FILLCELL_X1 PHY_1147 ();
 FILLCELL_X1 PHY_1148 ();
 FILLCELL_X1 PHY_1149 ();
 FILLCELL_X1 PHY_115 ();
 FILLCELL_X1 PHY_1150 ();
 FILLCELL_X1 PHY_1151 ();
 FILLCELL_X1 PHY_1152 ();
 FILLCELL_X1 PHY_1153 ();
 FILLCELL_X1 PHY_1154 ();
 FILLCELL_X1 PHY_1155 ();
 FILLCELL_X1 PHY_1156 ();
 FILLCELL_X1 PHY_1157 ();
 FILLCELL_X1 PHY_1158 ();
 FILLCELL_X1 PHY_1159 ();
 FILLCELL_X1 PHY_116 ();
 FILLCELL_X1 PHY_1160 ();
 FILLCELL_X1 PHY_1161 ();
 FILLCELL_X1 PHY_1162 ();
 FILLCELL_X1 PHY_1163 ();
 FILLCELL_X1 PHY_1164 ();
 FILLCELL_X1 PHY_1165 ();
 FILLCELL_X1 PHY_1166 ();
 FILLCELL_X1 PHY_1167 ();
 FILLCELL_X1 PHY_1168 ();
 FILLCELL_X1 PHY_1169 ();
 FILLCELL_X1 PHY_117 ();
 FILLCELL_X1 PHY_1170 ();
 FILLCELL_X1 PHY_1171 ();
 FILLCELL_X1 PHY_1172 ();
 FILLCELL_X1 PHY_1173 ();
 FILLCELL_X1 PHY_1174 ();
 FILLCELL_X1 PHY_1175 ();
 FILLCELL_X1 PHY_1176 ();
 FILLCELL_X1 PHY_1177 ();
 FILLCELL_X1 PHY_1178 ();
 FILLCELL_X1 PHY_1179 ();
 FILLCELL_X1 PHY_118 ();
 FILLCELL_X1 PHY_1180 ();
 FILLCELL_X1 PHY_1181 ();
 FILLCELL_X1 PHY_1182 ();
 FILLCELL_X1 PHY_1183 ();
 FILLCELL_X1 PHY_1184 ();
 FILLCELL_X1 PHY_1185 ();
 FILLCELL_X1 PHY_1186 ();
 FILLCELL_X1 PHY_1187 ();
 FILLCELL_X1 PHY_1188 ();
 FILLCELL_X1 PHY_1189 ();
 FILLCELL_X1 PHY_119 ();
 FILLCELL_X1 PHY_1190 ();
 FILLCELL_X1 PHY_1191 ();
 FILLCELL_X1 PHY_1192 ();
 FILLCELL_X1 PHY_1193 ();
 FILLCELL_X1 PHY_1194 ();
 FILLCELL_X1 PHY_1195 ();
 FILLCELL_X1 PHY_1196 ();
 FILLCELL_X1 PHY_1197 ();
 FILLCELL_X1 PHY_1198 ();
 FILLCELL_X1 PHY_1199 ();
 FILLCELL_X1 PHY_12 ();
 FILLCELL_X1 PHY_120 ();
 FILLCELL_X1 PHY_1200 ();
 FILLCELL_X1 PHY_1201 ();
 FILLCELL_X1 PHY_1202 ();
 FILLCELL_X1 PHY_1203 ();
 FILLCELL_X1 PHY_1204 ();
 FILLCELL_X1 PHY_1205 ();
 FILLCELL_X1 PHY_1206 ();
 FILLCELL_X1 PHY_1207 ();
 FILLCELL_X1 PHY_1208 ();
 FILLCELL_X1 PHY_1209 ();
 FILLCELL_X1 PHY_121 ();
 FILLCELL_X1 PHY_1210 ();
 FILLCELL_X1 PHY_1211 ();
 FILLCELL_X1 PHY_1212 ();
 FILLCELL_X1 PHY_1213 ();
 FILLCELL_X1 PHY_1214 ();
 FILLCELL_X1 PHY_1215 ();
 FILLCELL_X1 PHY_1216 ();
 FILLCELL_X1 PHY_1217 ();
 FILLCELL_X1 PHY_1218 ();
 FILLCELL_X1 PHY_1219 ();
 FILLCELL_X1 PHY_122 ();
 FILLCELL_X1 PHY_1220 ();
 FILLCELL_X1 PHY_1221 ();
 FILLCELL_X1 PHY_1222 ();
 FILLCELL_X1 PHY_1223 ();
 FILLCELL_X1 PHY_1224 ();
 FILLCELL_X1 PHY_1225 ();
 FILLCELL_X1 PHY_1226 ();
 FILLCELL_X1 PHY_1227 ();
 FILLCELL_X1 PHY_1228 ();
 FILLCELL_X1 PHY_1229 ();
 FILLCELL_X1 PHY_123 ();
 FILLCELL_X1 PHY_1230 ();
 FILLCELL_X1 PHY_1231 ();
 FILLCELL_X1 PHY_1232 ();
 FILLCELL_X1 PHY_1233 ();
 FILLCELL_X1 PHY_1234 ();
 FILLCELL_X1 PHY_1235 ();
 FILLCELL_X1 PHY_1236 ();
 FILLCELL_X1 PHY_1237 ();
 FILLCELL_X1 PHY_1238 ();
 FILLCELL_X1 PHY_1239 ();
 FILLCELL_X1 PHY_124 ();
 FILLCELL_X1 PHY_1240 ();
 FILLCELL_X1 PHY_1241 ();
 FILLCELL_X1 PHY_1242 ();
 FILLCELL_X1 PHY_1243 ();
 FILLCELL_X1 PHY_1244 ();
 FILLCELL_X1 PHY_1245 ();
 FILLCELL_X1 PHY_1246 ();
 FILLCELL_X1 PHY_1247 ();
 FILLCELL_X1 PHY_1248 ();
 FILLCELL_X1 PHY_1249 ();
 FILLCELL_X1 PHY_125 ();
 FILLCELL_X1 PHY_1250 ();
 FILLCELL_X1 PHY_1251 ();
 FILLCELL_X1 PHY_1252 ();
 FILLCELL_X1 PHY_1253 ();
 FILLCELL_X1 PHY_1254 ();
 FILLCELL_X1 PHY_1255 ();
 FILLCELL_X1 PHY_1256 ();
 FILLCELL_X1 PHY_1257 ();
 FILLCELL_X1 PHY_1258 ();
 FILLCELL_X1 PHY_1259 ();
 FILLCELL_X1 PHY_126 ();
 FILLCELL_X1 PHY_1260 ();
 FILLCELL_X1 PHY_1261 ();
 FILLCELL_X1 PHY_1262 ();
 FILLCELL_X1 PHY_1263 ();
 FILLCELL_X1 PHY_1264 ();
 FILLCELL_X1 PHY_1265 ();
 FILLCELL_X1 PHY_1266 ();
 FILLCELL_X1 PHY_1267 ();
 FILLCELL_X1 PHY_1268 ();
 FILLCELL_X1 PHY_1269 ();
 FILLCELL_X1 PHY_127 ();
 FILLCELL_X1 PHY_1270 ();
 FILLCELL_X1 PHY_1271 ();
 FILLCELL_X1 PHY_1272 ();
 FILLCELL_X1 PHY_1273 ();
 FILLCELL_X1 PHY_1274 ();
 FILLCELL_X1 PHY_1275 ();
 FILLCELL_X1 PHY_1276 ();
 FILLCELL_X1 PHY_1277 ();
 FILLCELL_X1 PHY_1278 ();
 FILLCELL_X1 PHY_1279 ();
 FILLCELL_X1 PHY_128 ();
 FILLCELL_X1 PHY_1280 ();
 FILLCELL_X1 PHY_1281 ();
 FILLCELL_X1 PHY_1282 ();
 FILLCELL_X1 PHY_1283 ();
 FILLCELL_X1 PHY_1284 ();
 FILLCELL_X1 PHY_1285 ();
 FILLCELL_X1 PHY_1286 ();
 FILLCELL_X1 PHY_1287 ();
 FILLCELL_X1 PHY_1288 ();
 FILLCELL_X1 PHY_1289 ();
 FILLCELL_X1 PHY_129 ();
 FILLCELL_X1 PHY_1290 ();
 FILLCELL_X1 PHY_1291 ();
 FILLCELL_X1 PHY_1292 ();
 FILLCELL_X1 PHY_1293 ();
 FILLCELL_X1 PHY_1294 ();
 FILLCELL_X1 PHY_1295 ();
 FILLCELL_X1 PHY_1296 ();
 FILLCELL_X1 PHY_1297 ();
 FILLCELL_X1 PHY_1298 ();
 FILLCELL_X1 PHY_1299 ();
 FILLCELL_X1 PHY_13 ();
 FILLCELL_X1 PHY_130 ();
 FILLCELL_X1 PHY_1300 ();
 FILLCELL_X1 PHY_1301 ();
 FILLCELL_X1 PHY_1302 ();
 FILLCELL_X1 PHY_1303 ();
 FILLCELL_X1 PHY_1304 ();
 FILLCELL_X1 PHY_1305 ();
 FILLCELL_X1 PHY_1306 ();
 FILLCELL_X1 PHY_1307 ();
 FILLCELL_X1 PHY_1308 ();
 FILLCELL_X1 PHY_1309 ();
 FILLCELL_X1 PHY_131 ();
 FILLCELL_X1 PHY_1310 ();
 FILLCELL_X1 PHY_1311 ();
 FILLCELL_X1 PHY_1312 ();
 FILLCELL_X1 PHY_1313 ();
 FILLCELL_X1 PHY_1314 ();
 FILLCELL_X1 PHY_1315 ();
 FILLCELL_X1 PHY_1316 ();
 FILLCELL_X1 PHY_1317 ();
 FILLCELL_X1 PHY_1318 ();
 FILLCELL_X1 PHY_1319 ();
 FILLCELL_X1 PHY_132 ();
 FILLCELL_X1 PHY_1320 ();
 FILLCELL_X1 PHY_1321 ();
 FILLCELL_X1 PHY_1322 ();
 FILLCELL_X1 PHY_1323 ();
 FILLCELL_X1 PHY_1324 ();
 FILLCELL_X1 PHY_1325 ();
 FILLCELL_X1 PHY_1326 ();
 FILLCELL_X1 PHY_1327 ();
 FILLCELL_X1 PHY_1328 ();
 FILLCELL_X1 PHY_1329 ();
 FILLCELL_X1 PHY_133 ();
 FILLCELL_X1 PHY_1330 ();
 FILLCELL_X1 PHY_1331 ();
 FILLCELL_X1 PHY_1332 ();
 FILLCELL_X1 PHY_1333 ();
 FILLCELL_X1 PHY_1334 ();
 FILLCELL_X1 PHY_1335 ();
 FILLCELL_X1 PHY_1336 ();
 FILLCELL_X1 PHY_1337 ();
 FILLCELL_X1 PHY_1338 ();
 FILLCELL_X1 PHY_1339 ();
 FILLCELL_X1 PHY_134 ();
 FILLCELL_X1 PHY_1340 ();
 FILLCELL_X1 PHY_1341 ();
 FILLCELL_X1 PHY_1342 ();
 FILLCELL_X1 PHY_1343 ();
 FILLCELL_X1 PHY_1344 ();
 FILLCELL_X1 PHY_1345 ();
 FILLCELL_X1 PHY_1346 ();
 FILLCELL_X1 PHY_1347 ();
 FILLCELL_X1 PHY_1348 ();
 FILLCELL_X1 PHY_1349 ();
 FILLCELL_X1 PHY_135 ();
 FILLCELL_X1 PHY_1350 ();
 FILLCELL_X1 PHY_1351 ();
 FILLCELL_X1 PHY_1352 ();
 FILLCELL_X1 PHY_1353 ();
 FILLCELL_X1 PHY_1354 ();
 FILLCELL_X1 PHY_1355 ();
 FILLCELL_X1 PHY_1356 ();
 FILLCELL_X1 PHY_1357 ();
 FILLCELL_X1 PHY_1358 ();
 FILLCELL_X1 PHY_1359 ();
 FILLCELL_X1 PHY_136 ();
 FILLCELL_X1 PHY_1360 ();
 FILLCELL_X1 PHY_1361 ();
 FILLCELL_X1 PHY_1362 ();
 FILLCELL_X1 PHY_1363 ();
 FILLCELL_X1 PHY_1364 ();
 FILLCELL_X1 PHY_1365 ();
 FILLCELL_X1 PHY_1366 ();
 FILLCELL_X1 PHY_1367 ();
 FILLCELL_X1 PHY_1368 ();
 FILLCELL_X1 PHY_1369 ();
 FILLCELL_X1 PHY_137 ();
 FILLCELL_X1 PHY_1370 ();
 FILLCELL_X1 PHY_1371 ();
 FILLCELL_X1 PHY_1372 ();
 FILLCELL_X1 PHY_1373 ();
 FILLCELL_X1 PHY_1374 ();
 FILLCELL_X1 PHY_1375 ();
 FILLCELL_X1 PHY_1376 ();
 FILLCELL_X1 PHY_1377 ();
 FILLCELL_X1 PHY_1378 ();
 FILLCELL_X1 PHY_1379 ();
 FILLCELL_X1 PHY_138 ();
 FILLCELL_X1 PHY_1380 ();
 FILLCELL_X1 PHY_1381 ();
 FILLCELL_X1 PHY_1382 ();
 FILLCELL_X1 PHY_1383 ();
 FILLCELL_X1 PHY_1384 ();
 FILLCELL_X1 PHY_1385 ();
 FILLCELL_X1 PHY_1386 ();
 FILLCELL_X1 PHY_1387 ();
 FILLCELL_X1 PHY_1388 ();
 FILLCELL_X1 PHY_1389 ();
 FILLCELL_X1 PHY_139 ();
 FILLCELL_X1 PHY_1390 ();
 FILLCELL_X1 PHY_1391 ();
 FILLCELL_X1 PHY_1392 ();
 FILLCELL_X1 PHY_1393 ();
 FILLCELL_X1 PHY_1394 ();
 FILLCELL_X1 PHY_1395 ();
 FILLCELL_X1 PHY_1396 ();
 FILLCELL_X1 PHY_1397 ();
 FILLCELL_X1 PHY_1398 ();
 FILLCELL_X1 PHY_1399 ();
 FILLCELL_X1 PHY_14 ();
 FILLCELL_X1 PHY_140 ();
 FILLCELL_X1 PHY_1400 ();
 FILLCELL_X1 PHY_1401 ();
 FILLCELL_X1 PHY_1402 ();
 FILLCELL_X1 PHY_1403 ();
 FILLCELL_X1 PHY_1404 ();
 FILLCELL_X1 PHY_1405 ();
 FILLCELL_X1 PHY_1406 ();
 FILLCELL_X1 PHY_1407 ();
 FILLCELL_X1 PHY_1408 ();
 FILLCELL_X1 PHY_1409 ();
 FILLCELL_X1 PHY_141 ();
 FILLCELL_X1 PHY_1410 ();
 FILLCELL_X1 PHY_1411 ();
 FILLCELL_X1 PHY_1412 ();
 FILLCELL_X1 PHY_1413 ();
 FILLCELL_X1 PHY_1414 ();
 FILLCELL_X1 PHY_1415 ();
 FILLCELL_X1 PHY_1416 ();
 FILLCELL_X1 PHY_1417 ();
 FILLCELL_X1 PHY_1418 ();
 FILLCELL_X1 PHY_1419 ();
 FILLCELL_X1 PHY_142 ();
 FILLCELL_X1 PHY_1420 ();
 FILLCELL_X1 PHY_1421 ();
 FILLCELL_X1 PHY_1422 ();
 FILLCELL_X1 PHY_1423 ();
 FILLCELL_X1 PHY_1424 ();
 FILLCELL_X1 PHY_1425 ();
 FILLCELL_X1 PHY_1426 ();
 FILLCELL_X1 PHY_1427 ();
 FILLCELL_X1 PHY_1428 ();
 FILLCELL_X1 PHY_1429 ();
 FILLCELL_X1 PHY_143 ();
 FILLCELL_X1 PHY_1430 ();
 FILLCELL_X1 PHY_1431 ();
 FILLCELL_X1 PHY_1432 ();
 FILLCELL_X1 PHY_1433 ();
 FILLCELL_X1 PHY_1434 ();
 FILLCELL_X1 PHY_1435 ();
 FILLCELL_X1 PHY_1436 ();
 FILLCELL_X1 PHY_1437 ();
 FILLCELL_X1 PHY_1438 ();
 FILLCELL_X1 PHY_1439 ();
 FILLCELL_X1 PHY_144 ();
 FILLCELL_X1 PHY_1440 ();
 FILLCELL_X1 PHY_1441 ();
 FILLCELL_X1 PHY_1442 ();
 FILLCELL_X1 PHY_1443 ();
 FILLCELL_X1 PHY_1444 ();
 FILLCELL_X1 PHY_1445 ();
 FILLCELL_X1 PHY_1446 ();
 FILLCELL_X1 PHY_1447 ();
 FILLCELL_X1 PHY_1448 ();
 FILLCELL_X1 PHY_1449 ();
 FILLCELL_X1 PHY_145 ();
 FILLCELL_X1 PHY_1450 ();
 FILLCELL_X1 PHY_1451 ();
 FILLCELL_X1 PHY_1452 ();
 FILLCELL_X1 PHY_1453 ();
 FILLCELL_X1 PHY_1454 ();
 FILLCELL_X1 PHY_1455 ();
 FILLCELL_X1 PHY_1456 ();
 FILLCELL_X1 PHY_1457 ();
 FILLCELL_X1 PHY_1458 ();
 FILLCELL_X1 PHY_1459 ();
 FILLCELL_X1 PHY_146 ();
 FILLCELL_X1 PHY_1460 ();
 FILLCELL_X1 PHY_1461 ();
 FILLCELL_X1 PHY_1462 ();
 FILLCELL_X1 PHY_1463 ();
 FILLCELL_X1 PHY_1464 ();
 FILLCELL_X1 PHY_1465 ();
 FILLCELL_X1 PHY_1466 ();
 FILLCELL_X1 PHY_1467 ();
 FILLCELL_X1 PHY_1468 ();
 FILLCELL_X1 PHY_1469 ();
 FILLCELL_X1 PHY_147 ();
 FILLCELL_X1 PHY_1470 ();
 FILLCELL_X1 PHY_1471 ();
 FILLCELL_X1 PHY_1472 ();
 FILLCELL_X1 PHY_1473 ();
 FILLCELL_X1 PHY_1474 ();
 FILLCELL_X1 PHY_1475 ();
 FILLCELL_X1 PHY_1476 ();
 FILLCELL_X1 PHY_1477 ();
 FILLCELL_X1 PHY_1478 ();
 FILLCELL_X1 PHY_1479 ();
 FILLCELL_X1 PHY_148 ();
 FILLCELL_X1 PHY_1480 ();
 FILLCELL_X1 PHY_1481 ();
 FILLCELL_X1 PHY_1482 ();
 FILLCELL_X1 PHY_1483 ();
 FILLCELL_X1 PHY_1484 ();
 FILLCELL_X1 PHY_1485 ();
 FILLCELL_X1 PHY_1486 ();
 FILLCELL_X1 PHY_1487 ();
 FILLCELL_X1 PHY_1488 ();
 FILLCELL_X1 PHY_1489 ();
 FILLCELL_X1 PHY_149 ();
 FILLCELL_X1 PHY_1490 ();
 FILLCELL_X1 PHY_1491 ();
 FILLCELL_X1 PHY_1492 ();
 FILLCELL_X1 PHY_1493 ();
 FILLCELL_X1 PHY_1494 ();
 FILLCELL_X1 PHY_1495 ();
 FILLCELL_X1 PHY_1496 ();
 FILLCELL_X1 PHY_1497 ();
 FILLCELL_X1 PHY_1498 ();
 FILLCELL_X1 PHY_1499 ();
 FILLCELL_X1 PHY_15 ();
 FILLCELL_X1 PHY_150 ();
 FILLCELL_X1 PHY_1500 ();
 FILLCELL_X1 PHY_1501 ();
 FILLCELL_X1 PHY_1502 ();
 FILLCELL_X1 PHY_1503 ();
 FILLCELL_X1 PHY_1504 ();
 FILLCELL_X1 PHY_1505 ();
 FILLCELL_X1 PHY_1506 ();
 FILLCELL_X1 PHY_1507 ();
 FILLCELL_X1 PHY_1508 ();
 FILLCELL_X1 PHY_1509 ();
 FILLCELL_X1 PHY_151 ();
 FILLCELL_X1 PHY_1510 ();
 FILLCELL_X1 PHY_1511 ();
 FILLCELL_X1 PHY_1512 ();
 FILLCELL_X1 PHY_1513 ();
 FILLCELL_X1 PHY_1514 ();
 FILLCELL_X1 PHY_1515 ();
 FILLCELL_X1 PHY_1516 ();
 FILLCELL_X1 PHY_1517 ();
 FILLCELL_X1 PHY_1518 ();
 FILLCELL_X1 PHY_1519 ();
 FILLCELL_X1 PHY_152 ();
 FILLCELL_X1 PHY_1520 ();
 FILLCELL_X1 PHY_1521 ();
 FILLCELL_X1 PHY_1522 ();
 FILLCELL_X1 PHY_1523 ();
 FILLCELL_X1 PHY_1524 ();
 FILLCELL_X1 PHY_1525 ();
 FILLCELL_X1 PHY_1526 ();
 FILLCELL_X1 PHY_1527 ();
 FILLCELL_X1 PHY_1528 ();
 FILLCELL_X1 PHY_1529 ();
 FILLCELL_X1 PHY_153 ();
 FILLCELL_X1 PHY_1530 ();
 FILLCELL_X1 PHY_1531 ();
 FILLCELL_X1 PHY_1532 ();
 FILLCELL_X1 PHY_1533 ();
 FILLCELL_X1 PHY_1534 ();
 FILLCELL_X1 PHY_1535 ();
 FILLCELL_X1 PHY_1536 ();
 FILLCELL_X1 PHY_1537 ();
 FILLCELL_X1 PHY_1538 ();
 FILLCELL_X1 PHY_1539 ();
 FILLCELL_X1 PHY_154 ();
 FILLCELL_X1 PHY_1540 ();
 FILLCELL_X1 PHY_1541 ();
 FILLCELL_X1 PHY_1542 ();
 FILLCELL_X1 PHY_1543 ();
 FILLCELL_X1 PHY_1544 ();
 FILLCELL_X1 PHY_1545 ();
 FILLCELL_X1 PHY_1546 ();
 FILLCELL_X1 PHY_1547 ();
 FILLCELL_X1 PHY_1548 ();
 FILLCELL_X1 PHY_1549 ();
 FILLCELL_X1 PHY_155 ();
 FILLCELL_X1 PHY_1550 ();
 FILLCELL_X1 PHY_1551 ();
 FILLCELL_X1 PHY_1552 ();
 FILLCELL_X1 PHY_1553 ();
 FILLCELL_X1 PHY_1554 ();
 FILLCELL_X1 PHY_1555 ();
 FILLCELL_X1 PHY_1556 ();
 FILLCELL_X1 PHY_1557 ();
 FILLCELL_X1 PHY_1558 ();
 FILLCELL_X1 PHY_1559 ();
 FILLCELL_X1 PHY_156 ();
 FILLCELL_X1 PHY_1560 ();
 FILLCELL_X1 PHY_1561 ();
 FILLCELL_X1 PHY_1562 ();
 FILLCELL_X1 PHY_1563 ();
 FILLCELL_X1 PHY_1564 ();
 FILLCELL_X1 PHY_1565 ();
 FILLCELL_X1 PHY_1566 ();
 FILLCELL_X1 PHY_1567 ();
 FILLCELL_X1 PHY_1568 ();
 FILLCELL_X1 PHY_1569 ();
 FILLCELL_X1 PHY_157 ();
 FILLCELL_X1 PHY_1570 ();
 FILLCELL_X1 PHY_1571 ();
 FILLCELL_X1 PHY_1572 ();
 FILLCELL_X1 PHY_1573 ();
 FILLCELL_X1 PHY_1574 ();
 FILLCELL_X1 PHY_1575 ();
 FILLCELL_X1 PHY_1576 ();
 FILLCELL_X1 PHY_1577 ();
 FILLCELL_X1 PHY_1578 ();
 FILLCELL_X1 PHY_1579 ();
 FILLCELL_X1 PHY_158 ();
 FILLCELL_X1 PHY_1580 ();
 FILLCELL_X1 PHY_1581 ();
 FILLCELL_X1 PHY_1582 ();
 FILLCELL_X1 PHY_1583 ();
 FILLCELL_X1 PHY_1584 ();
 FILLCELL_X1 PHY_1585 ();
 FILLCELL_X1 PHY_1586 ();
 FILLCELL_X1 PHY_1587 ();
 FILLCELL_X1 PHY_1588 ();
 FILLCELL_X1 PHY_1589 ();
 FILLCELL_X1 PHY_159 ();
 FILLCELL_X1 PHY_1590 ();
 FILLCELL_X1 PHY_1591 ();
 FILLCELL_X1 PHY_1592 ();
 FILLCELL_X1 PHY_1593 ();
 FILLCELL_X1 PHY_1594 ();
 FILLCELL_X1 PHY_1595 ();
 FILLCELL_X1 PHY_1596 ();
 FILLCELL_X1 PHY_1597 ();
 FILLCELL_X1 PHY_1598 ();
 FILLCELL_X1 PHY_1599 ();
 FILLCELL_X1 PHY_16 ();
 FILLCELL_X1 PHY_160 ();
 FILLCELL_X1 PHY_1600 ();
 FILLCELL_X1 PHY_1601 ();
 FILLCELL_X1 PHY_1602 ();
 FILLCELL_X1 PHY_1603 ();
 FILLCELL_X1 PHY_1604 ();
 FILLCELL_X1 PHY_1605 ();
 FILLCELL_X1 PHY_1606 ();
 FILLCELL_X1 PHY_1607 ();
 FILLCELL_X1 PHY_1608 ();
 FILLCELL_X1 PHY_1609 ();
 FILLCELL_X1 PHY_161 ();
 FILLCELL_X1 PHY_1610 ();
 FILLCELL_X1 PHY_1611 ();
 FILLCELL_X1 PHY_1612 ();
 FILLCELL_X1 PHY_1613 ();
 FILLCELL_X1 PHY_1614 ();
 FILLCELL_X1 PHY_1615 ();
 FILLCELL_X1 PHY_1616 ();
 FILLCELL_X1 PHY_1617 ();
 FILLCELL_X1 PHY_1618 ();
 FILLCELL_X1 PHY_1619 ();
 FILLCELL_X1 PHY_162 ();
 FILLCELL_X1 PHY_1620 ();
 FILLCELL_X1 PHY_1621 ();
 FILLCELL_X1 PHY_1622 ();
 FILLCELL_X1 PHY_1623 ();
 FILLCELL_X1 PHY_1624 ();
 FILLCELL_X1 PHY_1625 ();
 FILLCELL_X1 PHY_1626 ();
 FILLCELL_X1 PHY_1627 ();
 FILLCELL_X1 PHY_1628 ();
 FILLCELL_X1 PHY_1629 ();
 FILLCELL_X1 PHY_163 ();
 FILLCELL_X1 PHY_1630 ();
 FILLCELL_X1 PHY_1631 ();
 FILLCELL_X1 PHY_1632 ();
 FILLCELL_X1 PHY_1633 ();
 FILLCELL_X1 PHY_1634 ();
 FILLCELL_X1 PHY_1635 ();
 FILLCELL_X1 PHY_1636 ();
 FILLCELL_X1 PHY_1637 ();
 FILLCELL_X1 PHY_1638 ();
 FILLCELL_X1 PHY_1639 ();
 FILLCELL_X1 PHY_164 ();
 FILLCELL_X1 PHY_1640 ();
 FILLCELL_X1 PHY_1641 ();
 FILLCELL_X1 PHY_1642 ();
 FILLCELL_X1 PHY_1643 ();
 FILLCELL_X1 PHY_1644 ();
 FILLCELL_X1 PHY_1645 ();
 FILLCELL_X1 PHY_1646 ();
 FILLCELL_X1 PHY_1647 ();
 FILLCELL_X1 PHY_1648 ();
 FILLCELL_X1 PHY_1649 ();
 FILLCELL_X1 PHY_165 ();
 FILLCELL_X1 PHY_1650 ();
 FILLCELL_X1 PHY_1651 ();
 FILLCELL_X1 PHY_1652 ();
 FILLCELL_X1 PHY_1653 ();
 FILLCELL_X1 PHY_1654 ();
 FILLCELL_X1 PHY_1655 ();
 FILLCELL_X1 PHY_1656 ();
 FILLCELL_X1 PHY_1657 ();
 FILLCELL_X1 PHY_1658 ();
 FILLCELL_X1 PHY_1659 ();
 FILLCELL_X1 PHY_166 ();
 FILLCELL_X1 PHY_1660 ();
 FILLCELL_X1 PHY_1661 ();
 FILLCELL_X1 PHY_1662 ();
 FILLCELL_X1 PHY_1663 ();
 FILLCELL_X1 PHY_1664 ();
 FILLCELL_X1 PHY_1665 ();
 FILLCELL_X1 PHY_1666 ();
 FILLCELL_X1 PHY_1667 ();
 FILLCELL_X1 PHY_1668 ();
 FILLCELL_X1 PHY_1669 ();
 FILLCELL_X1 PHY_167 ();
 FILLCELL_X1 PHY_1670 ();
 FILLCELL_X1 PHY_1671 ();
 FILLCELL_X1 PHY_1672 ();
 FILLCELL_X1 PHY_1673 ();
 FILLCELL_X1 PHY_1674 ();
 FILLCELL_X1 PHY_1675 ();
 FILLCELL_X1 PHY_1676 ();
 FILLCELL_X1 PHY_1677 ();
 FILLCELL_X1 PHY_1678 ();
 FILLCELL_X1 PHY_1679 ();
 FILLCELL_X1 PHY_168 ();
 FILLCELL_X1 PHY_1680 ();
 FILLCELL_X1 PHY_1681 ();
 FILLCELL_X1 PHY_1682 ();
 FILLCELL_X1 PHY_1683 ();
 FILLCELL_X1 PHY_1684 ();
 FILLCELL_X1 PHY_1685 ();
 FILLCELL_X1 PHY_1686 ();
 FILLCELL_X1 PHY_1687 ();
 FILLCELL_X1 PHY_1688 ();
 FILLCELL_X1 PHY_1689 ();
 FILLCELL_X1 PHY_169 ();
 FILLCELL_X1 PHY_1690 ();
 FILLCELL_X1 PHY_1691 ();
 FILLCELL_X1 PHY_1692 ();
 FILLCELL_X1 PHY_1693 ();
 FILLCELL_X1 PHY_1694 ();
 FILLCELL_X1 PHY_1695 ();
 FILLCELL_X1 PHY_1696 ();
 FILLCELL_X1 PHY_1697 ();
 FILLCELL_X1 PHY_1698 ();
 FILLCELL_X1 PHY_1699 ();
 FILLCELL_X1 PHY_17 ();
 FILLCELL_X1 PHY_170 ();
 FILLCELL_X1 PHY_1700 ();
 FILLCELL_X1 PHY_1701 ();
 FILLCELL_X1 PHY_1702 ();
 FILLCELL_X1 PHY_1703 ();
 FILLCELL_X1 PHY_1704 ();
 FILLCELL_X1 PHY_1705 ();
 FILLCELL_X1 PHY_1706 ();
 FILLCELL_X1 PHY_1707 ();
 FILLCELL_X1 PHY_1708 ();
 FILLCELL_X1 PHY_1709 ();
 FILLCELL_X1 PHY_171 ();
 FILLCELL_X1 PHY_1710 ();
 FILLCELL_X1 PHY_1711 ();
 FILLCELL_X1 PHY_1712 ();
 FILLCELL_X1 PHY_1713 ();
 FILLCELL_X1 PHY_1714 ();
 FILLCELL_X1 PHY_1715 ();
 FILLCELL_X1 PHY_1716 ();
 FILLCELL_X1 PHY_1717 ();
 FILLCELL_X1 PHY_1718 ();
 FILLCELL_X1 PHY_1719 ();
 FILLCELL_X1 PHY_172 ();
 FILLCELL_X1 PHY_1720 ();
 FILLCELL_X1 PHY_1721 ();
 FILLCELL_X1 PHY_1722 ();
 FILLCELL_X1 PHY_1723 ();
 FILLCELL_X1 PHY_1724 ();
 FILLCELL_X1 PHY_1725 ();
 FILLCELL_X1 PHY_1726 ();
 FILLCELL_X1 PHY_1727 ();
 FILLCELL_X1 PHY_1728 ();
 FILLCELL_X1 PHY_1729 ();
 FILLCELL_X1 PHY_173 ();
 FILLCELL_X1 PHY_1730 ();
 FILLCELL_X1 PHY_1731 ();
 FILLCELL_X1 PHY_1732 ();
 FILLCELL_X1 PHY_1733 ();
 FILLCELL_X1 PHY_1734 ();
 FILLCELL_X1 PHY_1735 ();
 FILLCELL_X1 PHY_1736 ();
 FILLCELL_X1 PHY_1737 ();
 FILLCELL_X1 PHY_1738 ();
 FILLCELL_X1 PHY_1739 ();
 FILLCELL_X1 PHY_174 ();
 FILLCELL_X1 PHY_1740 ();
 FILLCELL_X1 PHY_1741 ();
 FILLCELL_X1 PHY_1742 ();
 FILLCELL_X1 PHY_1743 ();
 FILLCELL_X1 PHY_1744 ();
 FILLCELL_X1 PHY_1745 ();
 FILLCELL_X1 PHY_1746 ();
 FILLCELL_X1 PHY_1747 ();
 FILLCELL_X1 PHY_1748 ();
 FILLCELL_X1 PHY_1749 ();
 FILLCELL_X1 PHY_175 ();
 FILLCELL_X1 PHY_1750 ();
 FILLCELL_X1 PHY_1751 ();
 FILLCELL_X1 PHY_1752 ();
 FILLCELL_X1 PHY_1753 ();
 FILLCELL_X1 PHY_1754 ();
 FILLCELL_X1 PHY_1755 ();
 FILLCELL_X1 PHY_1756 ();
 FILLCELL_X1 PHY_1757 ();
 FILLCELL_X1 PHY_1758 ();
 FILLCELL_X1 PHY_1759 ();
 FILLCELL_X1 PHY_176 ();
 FILLCELL_X1 PHY_1760 ();
 FILLCELL_X1 PHY_1761 ();
 FILLCELL_X1 PHY_1762 ();
 FILLCELL_X1 PHY_1763 ();
 FILLCELL_X1 PHY_1764 ();
 FILLCELL_X1 PHY_1765 ();
 FILLCELL_X1 PHY_1766 ();
 FILLCELL_X1 PHY_1767 ();
 FILLCELL_X1 PHY_1768 ();
 FILLCELL_X1 PHY_1769 ();
 FILLCELL_X1 PHY_177 ();
 FILLCELL_X1 PHY_1770 ();
 FILLCELL_X1 PHY_1771 ();
 FILLCELL_X1 PHY_1772 ();
 FILLCELL_X1 PHY_1773 ();
 FILLCELL_X1 PHY_1774 ();
 FILLCELL_X1 PHY_1775 ();
 FILLCELL_X1 PHY_1776 ();
 FILLCELL_X1 PHY_1777 ();
 FILLCELL_X1 PHY_1778 ();
 FILLCELL_X1 PHY_1779 ();
 FILLCELL_X1 PHY_178 ();
 FILLCELL_X1 PHY_1780 ();
 FILLCELL_X1 PHY_1781 ();
 FILLCELL_X1 PHY_1782 ();
 FILLCELL_X1 PHY_1783 ();
 FILLCELL_X1 PHY_1784 ();
 FILLCELL_X1 PHY_1785 ();
 FILLCELL_X1 PHY_1786 ();
 FILLCELL_X1 PHY_1787 ();
 FILLCELL_X1 PHY_1788 ();
 FILLCELL_X1 PHY_1789 ();
 FILLCELL_X1 PHY_179 ();
 FILLCELL_X1 PHY_1790 ();
 FILLCELL_X1 PHY_1791 ();
 FILLCELL_X1 PHY_1792 ();
 FILLCELL_X1 PHY_1793 ();
 FILLCELL_X1 PHY_1794 ();
 FILLCELL_X1 PHY_1795 ();
 FILLCELL_X1 PHY_1796 ();
 FILLCELL_X1 PHY_1797 ();
 FILLCELL_X1 PHY_1798 ();
 FILLCELL_X1 PHY_1799 ();
 FILLCELL_X1 PHY_18 ();
 FILLCELL_X1 PHY_180 ();
 FILLCELL_X1 PHY_1800 ();
 FILLCELL_X1 PHY_1801 ();
 FILLCELL_X1 PHY_1802 ();
 FILLCELL_X1 PHY_1803 ();
 FILLCELL_X1 PHY_1804 ();
 FILLCELL_X1 PHY_1805 ();
 FILLCELL_X1 PHY_1806 ();
 FILLCELL_X1 PHY_1807 ();
 FILLCELL_X1 PHY_1808 ();
 FILLCELL_X1 PHY_1809 ();
 FILLCELL_X1 PHY_181 ();
 FILLCELL_X1 PHY_1810 ();
 FILLCELL_X1 PHY_1811 ();
 FILLCELL_X1 PHY_1812 ();
 FILLCELL_X1 PHY_1813 ();
 FILLCELL_X1 PHY_1814 ();
 FILLCELL_X1 PHY_1815 ();
 FILLCELL_X1 PHY_1816 ();
 FILLCELL_X1 PHY_1817 ();
 FILLCELL_X1 PHY_1818 ();
 FILLCELL_X1 PHY_1819 ();
 FILLCELL_X1 PHY_182 ();
 FILLCELL_X1 PHY_1820 ();
 FILLCELL_X1 PHY_1821 ();
 FILLCELL_X1 PHY_1822 ();
 FILLCELL_X1 PHY_1823 ();
 FILLCELL_X1 PHY_1824 ();
 FILLCELL_X1 PHY_1825 ();
 FILLCELL_X1 PHY_1826 ();
 FILLCELL_X1 PHY_1827 ();
 FILLCELL_X1 PHY_1828 ();
 FILLCELL_X1 PHY_1829 ();
 FILLCELL_X1 PHY_183 ();
 FILLCELL_X1 PHY_1830 ();
 FILLCELL_X1 PHY_1831 ();
 FILLCELL_X1 PHY_1832 ();
 FILLCELL_X1 PHY_1833 ();
 FILLCELL_X1 PHY_1834 ();
 FILLCELL_X1 PHY_1835 ();
 FILLCELL_X1 PHY_1836 ();
 FILLCELL_X1 PHY_1837 ();
 FILLCELL_X1 PHY_1838 ();
 FILLCELL_X1 PHY_1839 ();
 FILLCELL_X1 PHY_184 ();
 FILLCELL_X1 PHY_1840 ();
 FILLCELL_X1 PHY_1841 ();
 FILLCELL_X1 PHY_1842 ();
 FILLCELL_X1 PHY_1843 ();
 FILLCELL_X1 PHY_1844 ();
 FILLCELL_X1 PHY_1845 ();
 FILLCELL_X1 PHY_1846 ();
 FILLCELL_X1 PHY_1847 ();
 FILLCELL_X1 PHY_1848 ();
 FILLCELL_X1 PHY_1849 ();
 FILLCELL_X1 PHY_185 ();
 FILLCELL_X1 PHY_1850 ();
 FILLCELL_X1 PHY_1851 ();
 FILLCELL_X1 PHY_1852 ();
 FILLCELL_X1 PHY_1853 ();
 FILLCELL_X1 PHY_1854 ();
 FILLCELL_X1 PHY_1855 ();
 FILLCELL_X1 PHY_1856 ();
 FILLCELL_X1 PHY_1857 ();
 FILLCELL_X1 PHY_1858 ();
 FILLCELL_X1 PHY_1859 ();
 FILLCELL_X1 PHY_186 ();
 FILLCELL_X1 PHY_1860 ();
 FILLCELL_X1 PHY_1861 ();
 FILLCELL_X1 PHY_1862 ();
 FILLCELL_X1 PHY_1863 ();
 FILLCELL_X1 PHY_1864 ();
 FILLCELL_X1 PHY_1865 ();
 FILLCELL_X1 PHY_1866 ();
 FILLCELL_X1 PHY_1867 ();
 FILLCELL_X1 PHY_1868 ();
 FILLCELL_X1 PHY_1869 ();
 FILLCELL_X1 PHY_187 ();
 FILLCELL_X1 PHY_1870 ();
 FILLCELL_X1 PHY_1871 ();
 FILLCELL_X1 PHY_1872 ();
 FILLCELL_X1 PHY_1873 ();
 FILLCELL_X1 PHY_1874 ();
 FILLCELL_X1 PHY_1875 ();
 FILLCELL_X1 PHY_1876 ();
 FILLCELL_X1 PHY_1877 ();
 FILLCELL_X1 PHY_1878 ();
 FILLCELL_X1 PHY_1879 ();
 FILLCELL_X1 PHY_188 ();
 FILLCELL_X1 PHY_1880 ();
 FILLCELL_X1 PHY_1881 ();
 FILLCELL_X1 PHY_1882 ();
 FILLCELL_X1 PHY_1883 ();
 FILLCELL_X1 PHY_1884 ();
 FILLCELL_X1 PHY_1885 ();
 FILLCELL_X1 PHY_1886 ();
 FILLCELL_X1 PHY_1887 ();
 FILLCELL_X1 PHY_1888 ();
 FILLCELL_X1 PHY_1889 ();
 FILLCELL_X1 PHY_189 ();
 FILLCELL_X1 PHY_1890 ();
 FILLCELL_X1 PHY_1891 ();
 FILLCELL_X1 PHY_1892 ();
 FILLCELL_X1 PHY_1893 ();
 FILLCELL_X1 PHY_1894 ();
 FILLCELL_X1 PHY_1895 ();
 FILLCELL_X1 PHY_1896 ();
 FILLCELL_X1 PHY_1897 ();
 FILLCELL_X1 PHY_1898 ();
 FILLCELL_X1 PHY_1899 ();
 FILLCELL_X1 PHY_19 ();
 FILLCELL_X1 PHY_190 ();
 FILLCELL_X1 PHY_1900 ();
 FILLCELL_X1 PHY_1901 ();
 FILLCELL_X1 PHY_1902 ();
 FILLCELL_X1 PHY_1903 ();
 FILLCELL_X1 PHY_1904 ();
 FILLCELL_X1 PHY_1905 ();
 FILLCELL_X1 PHY_1906 ();
 FILLCELL_X1 PHY_1907 ();
 FILLCELL_X1 PHY_1908 ();
 FILLCELL_X1 PHY_1909 ();
 FILLCELL_X1 PHY_191 ();
 FILLCELL_X1 PHY_1910 ();
 FILLCELL_X1 PHY_1911 ();
 FILLCELL_X1 PHY_1912 ();
 FILLCELL_X1 PHY_1913 ();
 FILLCELL_X1 PHY_1914 ();
 FILLCELL_X1 PHY_1915 ();
 FILLCELL_X1 PHY_1916 ();
 FILLCELL_X1 PHY_1917 ();
 FILLCELL_X1 PHY_1918 ();
 FILLCELL_X1 PHY_1919 ();
 FILLCELL_X1 PHY_192 ();
 FILLCELL_X1 PHY_1920 ();
 FILLCELL_X1 PHY_1921 ();
 FILLCELL_X1 PHY_1922 ();
 FILLCELL_X1 PHY_1923 ();
 FILLCELL_X1 PHY_1924 ();
 FILLCELL_X1 PHY_1925 ();
 FILLCELL_X1 PHY_1926 ();
 FILLCELL_X1 PHY_1927 ();
 FILLCELL_X1 PHY_1928 ();
 FILLCELL_X1 PHY_1929 ();
 FILLCELL_X1 PHY_193 ();
 FILLCELL_X1 PHY_1930 ();
 FILLCELL_X1 PHY_1931 ();
 FILLCELL_X1 PHY_1932 ();
 FILLCELL_X1 PHY_1933 ();
 FILLCELL_X1 PHY_1934 ();
 FILLCELL_X1 PHY_1935 ();
 FILLCELL_X1 PHY_1936 ();
 FILLCELL_X1 PHY_1937 ();
 FILLCELL_X1 PHY_1938 ();
 FILLCELL_X1 PHY_1939 ();
 FILLCELL_X1 PHY_194 ();
 FILLCELL_X1 PHY_1940 ();
 FILLCELL_X1 PHY_1941 ();
 FILLCELL_X1 PHY_1942 ();
 FILLCELL_X1 PHY_1943 ();
 FILLCELL_X1 PHY_1944 ();
 FILLCELL_X1 PHY_1945 ();
 FILLCELL_X1 PHY_1946 ();
 FILLCELL_X1 PHY_1947 ();
 FILLCELL_X1 PHY_1948 ();
 FILLCELL_X1 PHY_1949 ();
 FILLCELL_X1 PHY_195 ();
 FILLCELL_X1 PHY_1950 ();
 FILLCELL_X1 PHY_1951 ();
 FILLCELL_X1 PHY_1952 ();
 FILLCELL_X1 PHY_1953 ();
 FILLCELL_X1 PHY_1954 ();
 FILLCELL_X1 PHY_1955 ();
 FILLCELL_X1 PHY_1956 ();
 FILLCELL_X1 PHY_1957 ();
 FILLCELL_X1 PHY_1958 ();
 FILLCELL_X1 PHY_1959 ();
 FILLCELL_X1 PHY_196 ();
 FILLCELL_X1 PHY_1960 ();
 FILLCELL_X1 PHY_1961 ();
 FILLCELL_X1 PHY_1962 ();
 FILLCELL_X1 PHY_1963 ();
 FILLCELL_X1 PHY_1964 ();
 FILLCELL_X1 PHY_1965 ();
 FILLCELL_X1 PHY_1966 ();
 FILLCELL_X1 PHY_1967 ();
 FILLCELL_X1 PHY_1968 ();
 FILLCELL_X1 PHY_1969 ();
 FILLCELL_X1 PHY_197 ();
 FILLCELL_X1 PHY_1970 ();
 FILLCELL_X1 PHY_1971 ();
 FILLCELL_X1 PHY_1972 ();
 FILLCELL_X1 PHY_1973 ();
 FILLCELL_X1 PHY_1974 ();
 FILLCELL_X1 PHY_1975 ();
 FILLCELL_X1 PHY_1976 ();
 FILLCELL_X1 PHY_1977 ();
 FILLCELL_X1 PHY_1978 ();
 FILLCELL_X1 PHY_1979 ();
 FILLCELL_X1 PHY_198 ();
 FILLCELL_X1 PHY_1980 ();
 FILLCELL_X1 PHY_1981 ();
 FILLCELL_X1 PHY_1982 ();
 FILLCELL_X1 PHY_1983 ();
 FILLCELL_X1 PHY_1984 ();
 FILLCELL_X1 PHY_1985 ();
 FILLCELL_X1 PHY_1986 ();
 FILLCELL_X1 PHY_1987 ();
 FILLCELL_X1 PHY_1988 ();
 FILLCELL_X1 PHY_1989 ();
 FILLCELL_X1 PHY_199 ();
 FILLCELL_X1 PHY_1990 ();
 FILLCELL_X1 PHY_1991 ();
 FILLCELL_X1 PHY_1992 ();
 FILLCELL_X1 PHY_1993 ();
 FILLCELL_X1 PHY_1994 ();
 FILLCELL_X1 PHY_1995 ();
 FILLCELL_X1 PHY_1996 ();
 FILLCELL_X1 PHY_1997 ();
 FILLCELL_X1 PHY_1998 ();
 FILLCELL_X1 PHY_1999 ();
 FILLCELL_X1 PHY_2 ();
 FILLCELL_X1 PHY_20 ();
 FILLCELL_X1 PHY_200 ();
 FILLCELL_X1 PHY_2000 ();
 FILLCELL_X1 PHY_2001 ();
 FILLCELL_X1 PHY_2002 ();
 FILLCELL_X1 PHY_2003 ();
 FILLCELL_X1 PHY_2004 ();
 FILLCELL_X1 PHY_2005 ();
 FILLCELL_X1 PHY_2006 ();
 FILLCELL_X1 PHY_2007 ();
 FILLCELL_X1 PHY_2008 ();
 FILLCELL_X1 PHY_2009 ();
 FILLCELL_X1 PHY_201 ();
 FILLCELL_X1 PHY_2010 ();
 FILLCELL_X1 PHY_2011 ();
 FILLCELL_X1 PHY_2012 ();
 FILLCELL_X1 PHY_2013 ();
 FILLCELL_X1 PHY_2014 ();
 FILLCELL_X1 PHY_2015 ();
 FILLCELL_X1 PHY_2016 ();
 FILLCELL_X1 PHY_2017 ();
 FILLCELL_X1 PHY_2018 ();
 FILLCELL_X1 PHY_2019 ();
 FILLCELL_X1 PHY_202 ();
 FILLCELL_X1 PHY_2020 ();
 FILLCELL_X1 PHY_2021 ();
 FILLCELL_X1 PHY_2022 ();
 FILLCELL_X1 PHY_2023 ();
 FILLCELL_X1 PHY_2024 ();
 FILLCELL_X1 PHY_2025 ();
 FILLCELL_X1 PHY_2026 ();
 FILLCELL_X1 PHY_2027 ();
 FILLCELL_X1 PHY_2028 ();
 FILLCELL_X1 PHY_2029 ();
 FILLCELL_X1 PHY_203 ();
 FILLCELL_X1 PHY_2030 ();
 FILLCELL_X1 PHY_2031 ();
 FILLCELL_X1 PHY_2032 ();
 FILLCELL_X1 PHY_2033 ();
 FILLCELL_X1 PHY_2034 ();
 FILLCELL_X1 PHY_2035 ();
 FILLCELL_X1 PHY_2036 ();
 FILLCELL_X1 PHY_2037 ();
 FILLCELL_X1 PHY_2038 ();
 FILLCELL_X1 PHY_2039 ();
 FILLCELL_X1 PHY_204 ();
 FILLCELL_X1 PHY_2040 ();
 FILLCELL_X1 PHY_2041 ();
 FILLCELL_X1 PHY_2042 ();
 FILLCELL_X1 PHY_2043 ();
 FILLCELL_X1 PHY_2044 ();
 FILLCELL_X1 PHY_2045 ();
 FILLCELL_X1 PHY_2046 ();
 FILLCELL_X1 PHY_2047 ();
 FILLCELL_X1 PHY_2048 ();
 FILLCELL_X1 PHY_2049 ();
 FILLCELL_X1 PHY_205 ();
 FILLCELL_X1 PHY_2050 ();
 FILLCELL_X1 PHY_2051 ();
 FILLCELL_X1 PHY_2052 ();
 FILLCELL_X1 PHY_2053 ();
 FILLCELL_X1 PHY_2054 ();
 FILLCELL_X1 PHY_2055 ();
 FILLCELL_X1 PHY_2056 ();
 FILLCELL_X1 PHY_2057 ();
 FILLCELL_X1 PHY_2058 ();
 FILLCELL_X1 PHY_2059 ();
 FILLCELL_X1 PHY_206 ();
 FILLCELL_X1 PHY_2060 ();
 FILLCELL_X1 PHY_2061 ();
 FILLCELL_X1 PHY_2062 ();
 FILLCELL_X1 PHY_2063 ();
 FILLCELL_X1 PHY_2064 ();
 FILLCELL_X1 PHY_2065 ();
 FILLCELL_X1 PHY_2066 ();
 FILLCELL_X1 PHY_2067 ();
 FILLCELL_X1 PHY_2068 ();
 FILLCELL_X1 PHY_2069 ();
 FILLCELL_X1 PHY_207 ();
 FILLCELL_X1 PHY_2070 ();
 FILLCELL_X1 PHY_2071 ();
 FILLCELL_X1 PHY_2072 ();
 FILLCELL_X1 PHY_2073 ();
 FILLCELL_X1 PHY_2074 ();
 FILLCELL_X1 PHY_2075 ();
 FILLCELL_X1 PHY_2076 ();
 FILLCELL_X1 PHY_2077 ();
 FILLCELL_X1 PHY_2078 ();
 FILLCELL_X1 PHY_2079 ();
 FILLCELL_X1 PHY_208 ();
 FILLCELL_X1 PHY_2080 ();
 FILLCELL_X1 PHY_2081 ();
 FILLCELL_X1 PHY_2082 ();
 FILLCELL_X1 PHY_2083 ();
 FILLCELL_X1 PHY_2084 ();
 FILLCELL_X1 PHY_2085 ();
 FILLCELL_X1 PHY_2086 ();
 FILLCELL_X1 PHY_2087 ();
 FILLCELL_X1 PHY_2088 ();
 FILLCELL_X1 PHY_2089 ();
 FILLCELL_X1 PHY_209 ();
 FILLCELL_X1 PHY_2090 ();
 FILLCELL_X1 PHY_2091 ();
 FILLCELL_X1 PHY_2092 ();
 FILLCELL_X1 PHY_2093 ();
 FILLCELL_X1 PHY_2094 ();
 FILLCELL_X1 PHY_2095 ();
 FILLCELL_X1 PHY_2096 ();
 FILLCELL_X1 PHY_2097 ();
 FILLCELL_X1 PHY_2098 ();
 FILLCELL_X1 PHY_2099 ();
 FILLCELL_X1 PHY_21 ();
 FILLCELL_X1 PHY_210 ();
 FILLCELL_X1 PHY_2100 ();
 FILLCELL_X1 PHY_2101 ();
 FILLCELL_X1 PHY_2102 ();
 FILLCELL_X1 PHY_2103 ();
 FILLCELL_X1 PHY_2104 ();
 FILLCELL_X1 PHY_2105 ();
 FILLCELL_X1 PHY_2106 ();
 FILLCELL_X1 PHY_2107 ();
 FILLCELL_X1 PHY_2108 ();
 FILLCELL_X1 PHY_2109 ();
 FILLCELL_X1 PHY_211 ();
 FILLCELL_X1 PHY_2110 ();
 FILLCELL_X1 PHY_2111 ();
 FILLCELL_X1 PHY_2112 ();
 FILLCELL_X1 PHY_2113 ();
 FILLCELL_X1 PHY_2114 ();
 FILLCELL_X1 PHY_2115 ();
 FILLCELL_X1 PHY_2116 ();
 FILLCELL_X1 PHY_2117 ();
 FILLCELL_X1 PHY_2118 ();
 FILLCELL_X1 PHY_2119 ();
 FILLCELL_X1 PHY_212 ();
 FILLCELL_X1 PHY_2120 ();
 FILLCELL_X1 PHY_2121 ();
 FILLCELL_X1 PHY_2122 ();
 FILLCELL_X1 PHY_2123 ();
 FILLCELL_X1 PHY_2124 ();
 FILLCELL_X1 PHY_2125 ();
 FILLCELL_X1 PHY_2126 ();
 FILLCELL_X1 PHY_2127 ();
 FILLCELL_X1 PHY_2128 ();
 FILLCELL_X1 PHY_2129 ();
 FILLCELL_X1 PHY_213 ();
 FILLCELL_X1 PHY_2130 ();
 FILLCELL_X1 PHY_2131 ();
 FILLCELL_X1 PHY_2132 ();
 FILLCELL_X1 PHY_2133 ();
 FILLCELL_X1 PHY_2134 ();
 FILLCELL_X1 PHY_2135 ();
 FILLCELL_X1 PHY_2136 ();
 FILLCELL_X1 PHY_2137 ();
 FILLCELL_X1 PHY_2138 ();
 FILLCELL_X1 PHY_2139 ();
 FILLCELL_X1 PHY_214 ();
 FILLCELL_X1 PHY_2140 ();
 FILLCELL_X1 PHY_2141 ();
 FILLCELL_X1 PHY_2142 ();
 FILLCELL_X1 PHY_2143 ();
 FILLCELL_X1 PHY_2144 ();
 FILLCELL_X1 PHY_2145 ();
 FILLCELL_X1 PHY_2146 ();
 FILLCELL_X1 PHY_2147 ();
 FILLCELL_X1 PHY_2148 ();
 FILLCELL_X1 PHY_2149 ();
 FILLCELL_X1 PHY_215 ();
 FILLCELL_X1 PHY_2150 ();
 FILLCELL_X1 PHY_2151 ();
 FILLCELL_X1 PHY_2152 ();
 FILLCELL_X1 PHY_2153 ();
 FILLCELL_X1 PHY_2154 ();
 FILLCELL_X1 PHY_2155 ();
 FILLCELL_X1 PHY_2156 ();
 FILLCELL_X1 PHY_2157 ();
 FILLCELL_X1 PHY_2158 ();
 FILLCELL_X1 PHY_2159 ();
 FILLCELL_X1 PHY_216 ();
 FILLCELL_X1 PHY_2160 ();
 FILLCELL_X1 PHY_2161 ();
 FILLCELL_X1 PHY_2162 ();
 FILLCELL_X1 PHY_2163 ();
 FILLCELL_X1 PHY_2164 ();
 FILLCELL_X1 PHY_2165 ();
 FILLCELL_X1 PHY_2166 ();
 FILLCELL_X1 PHY_2167 ();
 FILLCELL_X1 PHY_2168 ();
 FILLCELL_X1 PHY_2169 ();
 FILLCELL_X1 PHY_217 ();
 FILLCELL_X1 PHY_2170 ();
 FILLCELL_X1 PHY_2171 ();
 FILLCELL_X1 PHY_2172 ();
 FILLCELL_X1 PHY_2173 ();
 FILLCELL_X1 PHY_2174 ();
 FILLCELL_X1 PHY_2175 ();
 FILLCELL_X1 PHY_2176 ();
 FILLCELL_X1 PHY_2177 ();
 FILLCELL_X1 PHY_2178 ();
 FILLCELL_X1 PHY_2179 ();
 FILLCELL_X1 PHY_218 ();
 FILLCELL_X1 PHY_2180 ();
 FILLCELL_X1 PHY_2181 ();
 FILLCELL_X1 PHY_2182 ();
 FILLCELL_X1 PHY_2183 ();
 FILLCELL_X1 PHY_2184 ();
 FILLCELL_X1 PHY_2185 ();
 FILLCELL_X1 PHY_2186 ();
 FILLCELL_X1 PHY_2187 ();
 FILLCELL_X1 PHY_2188 ();
 FILLCELL_X1 PHY_2189 ();
 FILLCELL_X1 PHY_219 ();
 FILLCELL_X1 PHY_2190 ();
 FILLCELL_X1 PHY_2191 ();
 FILLCELL_X1 PHY_2192 ();
 FILLCELL_X1 PHY_2193 ();
 FILLCELL_X1 PHY_2194 ();
 FILLCELL_X1 PHY_2195 ();
 FILLCELL_X1 PHY_2196 ();
 FILLCELL_X1 PHY_2197 ();
 FILLCELL_X1 PHY_2198 ();
 FILLCELL_X1 PHY_2199 ();
 FILLCELL_X1 PHY_22 ();
 FILLCELL_X1 PHY_220 ();
 FILLCELL_X1 PHY_2200 ();
 FILLCELL_X1 PHY_2201 ();
 FILLCELL_X1 PHY_2202 ();
 FILLCELL_X1 PHY_2203 ();
 FILLCELL_X1 PHY_2204 ();
 FILLCELL_X1 PHY_2205 ();
 FILLCELL_X1 PHY_2206 ();
 FILLCELL_X1 PHY_2207 ();
 FILLCELL_X1 PHY_2208 ();
 FILLCELL_X1 PHY_2209 ();
 FILLCELL_X1 PHY_221 ();
 FILLCELL_X1 PHY_2210 ();
 FILLCELL_X1 PHY_2211 ();
 FILLCELL_X1 PHY_2212 ();
 FILLCELL_X1 PHY_2213 ();
 FILLCELL_X1 PHY_2214 ();
 FILLCELL_X1 PHY_2215 ();
 FILLCELL_X1 PHY_2216 ();
 FILLCELL_X1 PHY_2217 ();
 FILLCELL_X1 PHY_2218 ();
 FILLCELL_X1 PHY_2219 ();
 FILLCELL_X1 PHY_222 ();
 FILLCELL_X1 PHY_2220 ();
 FILLCELL_X1 PHY_2221 ();
 FILLCELL_X1 PHY_2222 ();
 FILLCELL_X1 PHY_2223 ();
 FILLCELL_X1 PHY_2224 ();
 FILLCELL_X1 PHY_2225 ();
 FILLCELL_X1 PHY_2226 ();
 FILLCELL_X1 PHY_2227 ();
 FILLCELL_X1 PHY_2228 ();
 FILLCELL_X1 PHY_2229 ();
 FILLCELL_X1 PHY_223 ();
 FILLCELL_X1 PHY_2230 ();
 FILLCELL_X1 PHY_2231 ();
 FILLCELL_X1 PHY_2232 ();
 FILLCELL_X1 PHY_2233 ();
 FILLCELL_X1 PHY_2234 ();
 FILLCELL_X1 PHY_2235 ();
 FILLCELL_X1 PHY_2236 ();
 FILLCELL_X1 PHY_2237 ();
 FILLCELL_X1 PHY_2238 ();
 FILLCELL_X1 PHY_2239 ();
 FILLCELL_X1 PHY_224 ();
 FILLCELL_X1 PHY_2240 ();
 FILLCELL_X1 PHY_2241 ();
 FILLCELL_X1 PHY_2242 ();
 FILLCELL_X1 PHY_2243 ();
 FILLCELL_X1 PHY_2244 ();
 FILLCELL_X1 PHY_2245 ();
 FILLCELL_X1 PHY_2246 ();
 FILLCELL_X1 PHY_2247 ();
 FILLCELL_X1 PHY_2248 ();
 FILLCELL_X1 PHY_2249 ();
 FILLCELL_X1 PHY_225 ();
 FILLCELL_X1 PHY_2250 ();
 FILLCELL_X1 PHY_2251 ();
 FILLCELL_X1 PHY_2252 ();
 FILLCELL_X1 PHY_2253 ();
 FILLCELL_X1 PHY_2254 ();
 FILLCELL_X1 PHY_2255 ();
 FILLCELL_X1 PHY_2256 ();
 FILLCELL_X1 PHY_2257 ();
 FILLCELL_X1 PHY_2258 ();
 FILLCELL_X1 PHY_2259 ();
 FILLCELL_X1 PHY_226 ();
 FILLCELL_X1 PHY_2260 ();
 FILLCELL_X1 PHY_2261 ();
 FILLCELL_X1 PHY_2262 ();
 FILLCELL_X1 PHY_2263 ();
 FILLCELL_X1 PHY_2264 ();
 FILLCELL_X1 PHY_2265 ();
 FILLCELL_X1 PHY_2266 ();
 FILLCELL_X1 PHY_2267 ();
 FILLCELL_X1 PHY_2268 ();
 FILLCELL_X1 PHY_2269 ();
 FILLCELL_X1 PHY_227 ();
 FILLCELL_X1 PHY_2270 ();
 FILLCELL_X1 PHY_2271 ();
 FILLCELL_X1 PHY_2272 ();
 FILLCELL_X1 PHY_2273 ();
 FILLCELL_X1 PHY_2274 ();
 FILLCELL_X1 PHY_2275 ();
 FILLCELL_X1 PHY_2276 ();
 FILLCELL_X1 PHY_2277 ();
 FILLCELL_X1 PHY_2278 ();
 FILLCELL_X1 PHY_2279 ();
 FILLCELL_X1 PHY_228 ();
 FILLCELL_X1 PHY_2280 ();
 FILLCELL_X1 PHY_2281 ();
 FILLCELL_X1 PHY_2282 ();
 FILLCELL_X1 PHY_2283 ();
 FILLCELL_X1 PHY_2284 ();
 FILLCELL_X1 PHY_2285 ();
 FILLCELL_X1 PHY_2286 ();
 FILLCELL_X1 PHY_2287 ();
 FILLCELL_X1 PHY_2288 ();
 FILLCELL_X1 PHY_2289 ();
 FILLCELL_X1 PHY_229 ();
 FILLCELL_X1 PHY_2290 ();
 FILLCELL_X1 PHY_2291 ();
 FILLCELL_X1 PHY_2292 ();
 FILLCELL_X1 PHY_2293 ();
 FILLCELL_X1 PHY_2294 ();
 FILLCELL_X1 PHY_2295 ();
 FILLCELL_X1 PHY_2296 ();
 FILLCELL_X1 PHY_2297 ();
 FILLCELL_X1 PHY_2298 ();
 FILLCELL_X1 PHY_2299 ();
 FILLCELL_X1 PHY_23 ();
 FILLCELL_X1 PHY_230 ();
 FILLCELL_X1 PHY_2300 ();
 FILLCELL_X1 PHY_2301 ();
 FILLCELL_X1 PHY_2302 ();
 FILLCELL_X1 PHY_2303 ();
 FILLCELL_X1 PHY_2304 ();
 FILLCELL_X1 PHY_2305 ();
 FILLCELL_X1 PHY_2306 ();
 FILLCELL_X1 PHY_2307 ();
 FILLCELL_X1 PHY_2308 ();
 FILLCELL_X1 PHY_2309 ();
 FILLCELL_X1 PHY_231 ();
 FILLCELL_X1 PHY_2310 ();
 FILLCELL_X1 PHY_2311 ();
 FILLCELL_X1 PHY_2312 ();
 FILLCELL_X1 PHY_2313 ();
 FILLCELL_X1 PHY_2314 ();
 FILLCELL_X1 PHY_2315 ();
 FILLCELL_X1 PHY_2316 ();
 FILLCELL_X1 PHY_2317 ();
 FILLCELL_X1 PHY_2318 ();
 FILLCELL_X1 PHY_2319 ();
 FILLCELL_X1 PHY_232 ();
 FILLCELL_X1 PHY_2320 ();
 FILLCELL_X1 PHY_2321 ();
 FILLCELL_X1 PHY_2322 ();
 FILLCELL_X1 PHY_2323 ();
 FILLCELL_X1 PHY_2324 ();
 FILLCELL_X1 PHY_2325 ();
 FILLCELL_X1 PHY_2326 ();
 FILLCELL_X1 PHY_2327 ();
 FILLCELL_X1 PHY_2328 ();
 FILLCELL_X1 PHY_2329 ();
 FILLCELL_X1 PHY_233 ();
 FILLCELL_X1 PHY_2330 ();
 FILLCELL_X1 PHY_2331 ();
 FILLCELL_X1 PHY_2332 ();
 FILLCELL_X1 PHY_2333 ();
 FILLCELL_X1 PHY_2334 ();
 FILLCELL_X1 PHY_2335 ();
 FILLCELL_X1 PHY_2336 ();
 FILLCELL_X1 PHY_2337 ();
 FILLCELL_X1 PHY_2338 ();
 FILLCELL_X1 PHY_2339 ();
 FILLCELL_X1 PHY_234 ();
 FILLCELL_X1 PHY_2340 ();
 FILLCELL_X1 PHY_2341 ();
 FILLCELL_X1 PHY_2342 ();
 FILLCELL_X1 PHY_2343 ();
 FILLCELL_X1 PHY_2344 ();
 FILLCELL_X1 PHY_2345 ();
 FILLCELL_X1 PHY_2346 ();
 FILLCELL_X1 PHY_2347 ();
 FILLCELL_X1 PHY_2348 ();
 FILLCELL_X1 PHY_2349 ();
 FILLCELL_X1 PHY_235 ();
 FILLCELL_X1 PHY_2350 ();
 FILLCELL_X1 PHY_2351 ();
 FILLCELL_X1 PHY_2352 ();
 FILLCELL_X1 PHY_2353 ();
 FILLCELL_X1 PHY_2354 ();
 FILLCELL_X1 PHY_2355 ();
 FILLCELL_X1 PHY_2356 ();
 FILLCELL_X1 PHY_2357 ();
 FILLCELL_X1 PHY_2358 ();
 FILLCELL_X1 PHY_2359 ();
 FILLCELL_X1 PHY_236 ();
 FILLCELL_X1 PHY_2360 ();
 FILLCELL_X1 PHY_2361 ();
 FILLCELL_X1 PHY_2362 ();
 FILLCELL_X1 PHY_2363 ();
 FILLCELL_X1 PHY_2364 ();
 FILLCELL_X1 PHY_2365 ();
 FILLCELL_X1 PHY_2366 ();
 FILLCELL_X1 PHY_2367 ();
 FILLCELL_X1 PHY_2368 ();
 FILLCELL_X1 PHY_2369 ();
 FILLCELL_X1 PHY_237 ();
 FILLCELL_X1 PHY_2370 ();
 FILLCELL_X1 PHY_2371 ();
 FILLCELL_X1 PHY_2372 ();
 FILLCELL_X1 PHY_2373 ();
 FILLCELL_X1 PHY_2374 ();
 FILLCELL_X1 PHY_2375 ();
 FILLCELL_X1 PHY_2376 ();
 FILLCELL_X1 PHY_2377 ();
 FILLCELL_X1 PHY_2378 ();
 FILLCELL_X1 PHY_2379 ();
 FILLCELL_X1 PHY_238 ();
 FILLCELL_X1 PHY_2380 ();
 FILLCELL_X1 PHY_2381 ();
 FILLCELL_X1 PHY_2382 ();
 FILLCELL_X1 PHY_2383 ();
 FILLCELL_X1 PHY_2384 ();
 FILLCELL_X1 PHY_2385 ();
 FILLCELL_X1 PHY_2386 ();
 FILLCELL_X1 PHY_2387 ();
 FILLCELL_X1 PHY_2388 ();
 FILLCELL_X1 PHY_2389 ();
 FILLCELL_X1 PHY_239 ();
 FILLCELL_X1 PHY_2390 ();
 FILLCELL_X1 PHY_2391 ();
 FILLCELL_X1 PHY_2392 ();
 FILLCELL_X1 PHY_2393 ();
 FILLCELL_X1 PHY_2394 ();
 FILLCELL_X1 PHY_2395 ();
 FILLCELL_X1 PHY_2396 ();
 FILLCELL_X1 PHY_2397 ();
 FILLCELL_X1 PHY_2398 ();
 FILLCELL_X1 PHY_2399 ();
 FILLCELL_X1 PHY_24 ();
 FILLCELL_X1 PHY_240 ();
 FILLCELL_X1 PHY_2400 ();
 FILLCELL_X1 PHY_2401 ();
 FILLCELL_X1 PHY_2402 ();
 FILLCELL_X1 PHY_2403 ();
 FILLCELL_X1 PHY_2404 ();
 FILLCELL_X1 PHY_2405 ();
 FILLCELL_X1 PHY_2406 ();
 FILLCELL_X1 PHY_2407 ();
 FILLCELL_X1 PHY_2408 ();
 FILLCELL_X1 PHY_2409 ();
 FILLCELL_X1 PHY_241 ();
 FILLCELL_X1 PHY_2410 ();
 FILLCELL_X1 PHY_2411 ();
 FILLCELL_X1 PHY_2412 ();
 FILLCELL_X1 PHY_2413 ();
 FILLCELL_X1 PHY_2414 ();
 FILLCELL_X1 PHY_2415 ();
 FILLCELL_X1 PHY_2416 ();
 FILLCELL_X1 PHY_2417 ();
 FILLCELL_X1 PHY_2418 ();
 FILLCELL_X1 PHY_2419 ();
 FILLCELL_X1 PHY_242 ();
 FILLCELL_X1 PHY_2420 ();
 FILLCELL_X1 PHY_2421 ();
 FILLCELL_X1 PHY_2422 ();
 FILLCELL_X1 PHY_2423 ();
 FILLCELL_X1 PHY_2424 ();
 FILLCELL_X1 PHY_2425 ();
 FILLCELL_X1 PHY_2426 ();
 FILLCELL_X1 PHY_2427 ();
 FILLCELL_X1 PHY_2428 ();
 FILLCELL_X1 PHY_2429 ();
 FILLCELL_X1 PHY_243 ();
 FILLCELL_X1 PHY_2430 ();
 FILLCELL_X1 PHY_2431 ();
 FILLCELL_X1 PHY_2432 ();
 FILLCELL_X1 PHY_2433 ();
 FILLCELL_X1 PHY_2434 ();
 FILLCELL_X1 PHY_2435 ();
 FILLCELL_X1 PHY_2436 ();
 FILLCELL_X1 PHY_2437 ();
 FILLCELL_X1 PHY_2438 ();
 FILLCELL_X1 PHY_2439 ();
 FILLCELL_X1 PHY_244 ();
 FILLCELL_X1 PHY_2440 ();
 FILLCELL_X1 PHY_2441 ();
 FILLCELL_X1 PHY_2442 ();
 FILLCELL_X1 PHY_2443 ();
 FILLCELL_X1 PHY_2444 ();
 FILLCELL_X1 PHY_2445 ();
 FILLCELL_X1 PHY_2446 ();
 FILLCELL_X1 PHY_2447 ();
 FILLCELL_X1 PHY_2448 ();
 FILLCELL_X1 PHY_2449 ();
 FILLCELL_X1 PHY_245 ();
 FILLCELL_X1 PHY_2450 ();
 FILLCELL_X1 PHY_2451 ();
 FILLCELL_X1 PHY_2452 ();
 FILLCELL_X1 PHY_2453 ();
 FILLCELL_X1 PHY_2454 ();
 FILLCELL_X1 PHY_2455 ();
 FILLCELL_X1 PHY_2456 ();
 FILLCELL_X1 PHY_2457 ();
 FILLCELL_X1 PHY_2458 ();
 FILLCELL_X1 PHY_2459 ();
 FILLCELL_X1 PHY_246 ();
 FILLCELL_X1 PHY_2460 ();
 FILLCELL_X1 PHY_2461 ();
 FILLCELL_X1 PHY_2462 ();
 FILLCELL_X1 PHY_2463 ();
 FILLCELL_X1 PHY_2464 ();
 FILLCELL_X1 PHY_2465 ();
 FILLCELL_X1 PHY_2466 ();
 FILLCELL_X1 PHY_2467 ();
 FILLCELL_X1 PHY_2468 ();
 FILLCELL_X1 PHY_2469 ();
 FILLCELL_X1 PHY_247 ();
 FILLCELL_X1 PHY_2470 ();
 FILLCELL_X1 PHY_2471 ();
 FILLCELL_X1 PHY_2472 ();
 FILLCELL_X1 PHY_2473 ();
 FILLCELL_X1 PHY_2474 ();
 FILLCELL_X1 PHY_2475 ();
 FILLCELL_X1 PHY_2476 ();
 FILLCELL_X1 PHY_2477 ();
 FILLCELL_X1 PHY_2478 ();
 FILLCELL_X1 PHY_2479 ();
 FILLCELL_X1 PHY_248 ();
 FILLCELL_X1 PHY_2480 ();
 FILLCELL_X1 PHY_2481 ();
 FILLCELL_X1 PHY_2482 ();
 FILLCELL_X1 PHY_2483 ();
 FILLCELL_X1 PHY_2484 ();
 FILLCELL_X1 PHY_2485 ();
 FILLCELL_X1 PHY_2486 ();
 FILLCELL_X1 PHY_2487 ();
 FILLCELL_X1 PHY_2488 ();
 FILLCELL_X1 PHY_2489 ();
 FILLCELL_X1 PHY_249 ();
 FILLCELL_X1 PHY_2490 ();
 FILLCELL_X1 PHY_2491 ();
 FILLCELL_X1 PHY_2492 ();
 FILLCELL_X1 PHY_2493 ();
 FILLCELL_X1 PHY_2494 ();
 FILLCELL_X1 PHY_2495 ();
 FILLCELL_X1 PHY_2496 ();
 FILLCELL_X1 PHY_2497 ();
 FILLCELL_X1 PHY_2498 ();
 FILLCELL_X1 PHY_2499 ();
 FILLCELL_X1 PHY_25 ();
 FILLCELL_X1 PHY_250 ();
 FILLCELL_X1 PHY_2500 ();
 FILLCELL_X1 PHY_2501 ();
 FILLCELL_X1 PHY_2502 ();
 FILLCELL_X1 PHY_2503 ();
 FILLCELL_X1 PHY_2504 ();
 FILLCELL_X1 PHY_2505 ();
 FILLCELL_X1 PHY_2506 ();
 FILLCELL_X1 PHY_2507 ();
 FILLCELL_X1 PHY_2508 ();
 FILLCELL_X1 PHY_2509 ();
 FILLCELL_X1 PHY_251 ();
 FILLCELL_X1 PHY_2510 ();
 FILLCELL_X1 PHY_2511 ();
 FILLCELL_X1 PHY_2512 ();
 FILLCELL_X1 PHY_2513 ();
 FILLCELL_X1 PHY_2514 ();
 FILLCELL_X1 PHY_2515 ();
 FILLCELL_X1 PHY_2516 ();
 FILLCELL_X1 PHY_2517 ();
 FILLCELL_X1 PHY_2518 ();
 FILLCELL_X1 PHY_2519 ();
 FILLCELL_X1 PHY_252 ();
 FILLCELL_X1 PHY_2520 ();
 FILLCELL_X1 PHY_2521 ();
 FILLCELL_X1 PHY_2522 ();
 FILLCELL_X1 PHY_2523 ();
 FILLCELL_X1 PHY_2524 ();
 FILLCELL_X1 PHY_2525 ();
 FILLCELL_X1 PHY_2526 ();
 FILLCELL_X1 PHY_2527 ();
 FILLCELL_X1 PHY_2528 ();
 FILLCELL_X1 PHY_2529 ();
 FILLCELL_X1 PHY_253 ();
 FILLCELL_X1 PHY_2530 ();
 FILLCELL_X1 PHY_2531 ();
 FILLCELL_X1 PHY_2532 ();
 FILLCELL_X1 PHY_2533 ();
 FILLCELL_X1 PHY_2534 ();
 FILLCELL_X1 PHY_2535 ();
 FILLCELL_X1 PHY_2536 ();
 FILLCELL_X1 PHY_2537 ();
 FILLCELL_X1 PHY_2538 ();
 FILLCELL_X1 PHY_2539 ();
 FILLCELL_X1 PHY_254 ();
 FILLCELL_X1 PHY_2540 ();
 FILLCELL_X1 PHY_2541 ();
 FILLCELL_X1 PHY_2542 ();
 FILLCELL_X1 PHY_2543 ();
 FILLCELL_X1 PHY_2544 ();
 FILLCELL_X1 PHY_2545 ();
 FILLCELL_X1 PHY_2546 ();
 FILLCELL_X1 PHY_2547 ();
 FILLCELL_X1 PHY_2548 ();
 FILLCELL_X1 PHY_2549 ();
 FILLCELL_X1 PHY_255 ();
 FILLCELL_X1 PHY_2550 ();
 FILLCELL_X1 PHY_2551 ();
 FILLCELL_X1 PHY_2552 ();
 FILLCELL_X1 PHY_2553 ();
 FILLCELL_X1 PHY_2554 ();
 FILLCELL_X1 PHY_2555 ();
 FILLCELL_X1 PHY_2556 ();
 FILLCELL_X1 PHY_2557 ();
 FILLCELL_X1 PHY_2558 ();
 FILLCELL_X1 PHY_2559 ();
 FILLCELL_X1 PHY_256 ();
 FILLCELL_X1 PHY_2560 ();
 FILLCELL_X1 PHY_2561 ();
 FILLCELL_X1 PHY_2562 ();
 FILLCELL_X1 PHY_2563 ();
 FILLCELL_X1 PHY_2564 ();
 FILLCELL_X1 PHY_2565 ();
 FILLCELL_X1 PHY_2566 ();
 FILLCELL_X1 PHY_2567 ();
 FILLCELL_X1 PHY_2568 ();
 FILLCELL_X1 PHY_2569 ();
 FILLCELL_X1 PHY_257 ();
 FILLCELL_X1 PHY_2570 ();
 FILLCELL_X1 PHY_2571 ();
 FILLCELL_X1 PHY_2572 ();
 FILLCELL_X1 PHY_2573 ();
 FILLCELL_X1 PHY_2574 ();
 FILLCELL_X1 PHY_2575 ();
 FILLCELL_X1 PHY_2576 ();
 FILLCELL_X1 PHY_2577 ();
 FILLCELL_X1 PHY_2578 ();
 FILLCELL_X1 PHY_2579 ();
 FILLCELL_X1 PHY_258 ();
 FILLCELL_X1 PHY_2580 ();
 FILLCELL_X1 PHY_2581 ();
 FILLCELL_X1 PHY_2582 ();
 FILLCELL_X1 PHY_2583 ();
 FILLCELL_X1 PHY_2584 ();
 FILLCELL_X1 PHY_2585 ();
 FILLCELL_X1 PHY_2586 ();
 FILLCELL_X1 PHY_2587 ();
 FILLCELL_X1 PHY_2588 ();
 FILLCELL_X1 PHY_2589 ();
 FILLCELL_X1 PHY_259 ();
 FILLCELL_X1 PHY_2590 ();
 FILLCELL_X1 PHY_2591 ();
 FILLCELL_X1 PHY_2592 ();
 FILLCELL_X1 PHY_2593 ();
 FILLCELL_X1 PHY_2594 ();
 FILLCELL_X1 PHY_2595 ();
 FILLCELL_X1 PHY_2596 ();
 FILLCELL_X1 PHY_2597 ();
 FILLCELL_X1 PHY_2598 ();
 FILLCELL_X1 PHY_2599 ();
 FILLCELL_X1 PHY_26 ();
 FILLCELL_X1 PHY_260 ();
 FILLCELL_X1 PHY_2600 ();
 FILLCELL_X1 PHY_2601 ();
 FILLCELL_X1 PHY_2602 ();
 FILLCELL_X1 PHY_2603 ();
 FILLCELL_X1 PHY_2604 ();
 FILLCELL_X1 PHY_2605 ();
 FILLCELL_X1 PHY_2606 ();
 FILLCELL_X1 PHY_2607 ();
 FILLCELL_X1 PHY_2608 ();
 FILLCELL_X1 PHY_2609 ();
 FILLCELL_X1 PHY_261 ();
 FILLCELL_X1 PHY_2610 ();
 FILLCELL_X1 PHY_2611 ();
 FILLCELL_X1 PHY_2612 ();
 FILLCELL_X1 PHY_2613 ();
 FILLCELL_X1 PHY_2614 ();
 FILLCELL_X1 PHY_2615 ();
 FILLCELL_X1 PHY_2616 ();
 FILLCELL_X1 PHY_2617 ();
 FILLCELL_X1 PHY_2618 ();
 FILLCELL_X1 PHY_2619 ();
 FILLCELL_X1 PHY_262 ();
 FILLCELL_X1 PHY_2620 ();
 FILLCELL_X1 PHY_2621 ();
 FILLCELL_X1 PHY_2622 ();
 FILLCELL_X1 PHY_2623 ();
 FILLCELL_X1 PHY_2624 ();
 FILLCELL_X1 PHY_2625 ();
 FILLCELL_X1 PHY_2626 ();
 FILLCELL_X1 PHY_2627 ();
 FILLCELL_X1 PHY_2628 ();
 FILLCELL_X1 PHY_2629 ();
 FILLCELL_X1 PHY_263 ();
 FILLCELL_X1 PHY_2630 ();
 FILLCELL_X1 PHY_2631 ();
 FILLCELL_X1 PHY_2632 ();
 FILLCELL_X1 PHY_2633 ();
 FILLCELL_X1 PHY_2634 ();
 FILLCELL_X1 PHY_2635 ();
 FILLCELL_X1 PHY_2636 ();
 FILLCELL_X1 PHY_2637 ();
 FILLCELL_X1 PHY_2638 ();
 FILLCELL_X1 PHY_2639 ();
 FILLCELL_X1 PHY_264 ();
 FILLCELL_X1 PHY_2640 ();
 FILLCELL_X1 PHY_2641 ();
 FILLCELL_X1 PHY_2642 ();
 FILLCELL_X1 PHY_2643 ();
 FILLCELL_X1 PHY_2644 ();
 FILLCELL_X1 PHY_2645 ();
 FILLCELL_X1 PHY_2646 ();
 FILLCELL_X1 PHY_2647 ();
 FILLCELL_X1 PHY_2648 ();
 FILLCELL_X1 PHY_2649 ();
 FILLCELL_X1 PHY_265 ();
 FILLCELL_X1 PHY_2650 ();
 FILLCELL_X1 PHY_2651 ();
 FILLCELL_X1 PHY_2652 ();
 FILLCELL_X1 PHY_2653 ();
 FILLCELL_X1 PHY_2654 ();
 FILLCELL_X1 PHY_2655 ();
 FILLCELL_X1 PHY_2656 ();
 FILLCELL_X1 PHY_2657 ();
 FILLCELL_X1 PHY_2658 ();
 FILLCELL_X1 PHY_2659 ();
 FILLCELL_X1 PHY_266 ();
 FILLCELL_X1 PHY_2660 ();
 FILLCELL_X1 PHY_2661 ();
 FILLCELL_X1 PHY_2662 ();
 FILLCELL_X1 PHY_2663 ();
 FILLCELL_X1 PHY_2664 ();
 FILLCELL_X1 PHY_2665 ();
 FILLCELL_X1 PHY_2666 ();
 FILLCELL_X1 PHY_2667 ();
 FILLCELL_X1 PHY_2668 ();
 FILLCELL_X1 PHY_2669 ();
 FILLCELL_X1 PHY_267 ();
 FILLCELL_X1 PHY_2670 ();
 FILLCELL_X1 PHY_2671 ();
 FILLCELL_X1 PHY_2672 ();
 FILLCELL_X1 PHY_2673 ();
 FILLCELL_X1 PHY_2674 ();
 FILLCELL_X1 PHY_2675 ();
 FILLCELL_X1 PHY_2676 ();
 FILLCELL_X1 PHY_2677 ();
 FILLCELL_X1 PHY_2678 ();
 FILLCELL_X1 PHY_2679 ();
 FILLCELL_X1 PHY_268 ();
 FILLCELL_X1 PHY_2680 ();
 FILLCELL_X1 PHY_2681 ();
 FILLCELL_X1 PHY_2682 ();
 FILLCELL_X1 PHY_2683 ();
 FILLCELL_X1 PHY_2684 ();
 FILLCELL_X1 PHY_2685 ();
 FILLCELL_X1 PHY_2686 ();
 FILLCELL_X1 PHY_2687 ();
 FILLCELL_X1 PHY_2688 ();
 FILLCELL_X1 PHY_2689 ();
 FILLCELL_X1 PHY_269 ();
 FILLCELL_X1 PHY_2690 ();
 FILLCELL_X1 PHY_2691 ();
 FILLCELL_X1 PHY_2692 ();
 FILLCELL_X1 PHY_2693 ();
 FILLCELL_X1 PHY_2694 ();
 FILLCELL_X1 PHY_2695 ();
 FILLCELL_X1 PHY_2696 ();
 FILLCELL_X1 PHY_2697 ();
 FILLCELL_X1 PHY_2698 ();
 FILLCELL_X1 PHY_2699 ();
 FILLCELL_X1 PHY_27 ();
 FILLCELL_X1 PHY_270 ();
 FILLCELL_X1 PHY_2700 ();
 FILLCELL_X1 PHY_2701 ();
 FILLCELL_X1 PHY_2702 ();
 FILLCELL_X1 PHY_2703 ();
 FILLCELL_X1 PHY_2704 ();
 FILLCELL_X1 PHY_2705 ();
 FILLCELL_X1 PHY_2706 ();
 FILLCELL_X1 PHY_2707 ();
 FILLCELL_X1 PHY_2708 ();
 FILLCELL_X1 PHY_2709 ();
 FILLCELL_X1 PHY_271 ();
 FILLCELL_X1 PHY_2710 ();
 FILLCELL_X1 PHY_2711 ();
 FILLCELL_X1 PHY_2712 ();
 FILLCELL_X1 PHY_2713 ();
 FILLCELL_X1 PHY_2714 ();
 FILLCELL_X1 PHY_2715 ();
 FILLCELL_X1 PHY_2716 ();
 FILLCELL_X1 PHY_2717 ();
 FILLCELL_X1 PHY_2718 ();
 FILLCELL_X1 PHY_2719 ();
 FILLCELL_X1 PHY_272 ();
 FILLCELL_X1 PHY_2720 ();
 FILLCELL_X1 PHY_2721 ();
 FILLCELL_X1 PHY_2722 ();
 FILLCELL_X1 PHY_2723 ();
 FILLCELL_X1 PHY_2724 ();
 FILLCELL_X1 PHY_2725 ();
 FILLCELL_X1 PHY_2726 ();
 FILLCELL_X1 PHY_2727 ();
 FILLCELL_X1 PHY_2728 ();
 FILLCELL_X1 PHY_2729 ();
 FILLCELL_X1 PHY_273 ();
 FILLCELL_X1 PHY_2730 ();
 FILLCELL_X1 PHY_2731 ();
 FILLCELL_X1 PHY_2732 ();
 FILLCELL_X1 PHY_2733 ();
 FILLCELL_X1 PHY_2734 ();
 FILLCELL_X1 PHY_2735 ();
 FILLCELL_X1 PHY_2736 ();
 FILLCELL_X1 PHY_2737 ();
 FILLCELL_X1 PHY_2738 ();
 FILLCELL_X1 PHY_2739 ();
 FILLCELL_X1 PHY_274 ();
 FILLCELL_X1 PHY_2740 ();
 FILLCELL_X1 PHY_2741 ();
 FILLCELL_X1 PHY_2742 ();
 FILLCELL_X1 PHY_2743 ();
 FILLCELL_X1 PHY_2744 ();
 FILLCELL_X1 PHY_2745 ();
 FILLCELL_X1 PHY_2746 ();
 FILLCELL_X1 PHY_2747 ();
 FILLCELL_X1 PHY_2748 ();
 FILLCELL_X1 PHY_2749 ();
 FILLCELL_X1 PHY_275 ();
 FILLCELL_X1 PHY_2750 ();
 FILLCELL_X1 PHY_2751 ();
 FILLCELL_X1 PHY_2752 ();
 FILLCELL_X1 PHY_2753 ();
 FILLCELL_X1 PHY_2754 ();
 FILLCELL_X1 PHY_2755 ();
 FILLCELL_X1 PHY_2756 ();
 FILLCELL_X1 PHY_2757 ();
 FILLCELL_X1 PHY_2758 ();
 FILLCELL_X1 PHY_2759 ();
 FILLCELL_X1 PHY_276 ();
 FILLCELL_X1 PHY_2760 ();
 FILLCELL_X1 PHY_2761 ();
 FILLCELL_X1 PHY_2762 ();
 FILLCELL_X1 PHY_2763 ();
 FILLCELL_X1 PHY_2764 ();
 FILLCELL_X1 PHY_2765 ();
 FILLCELL_X1 PHY_2766 ();
 FILLCELL_X1 PHY_2767 ();
 FILLCELL_X1 PHY_2768 ();
 FILLCELL_X1 PHY_2769 ();
 FILLCELL_X1 PHY_277 ();
 FILLCELL_X1 PHY_2770 ();
 FILLCELL_X1 PHY_2771 ();
 FILLCELL_X1 PHY_2772 ();
 FILLCELL_X1 PHY_2773 ();
 FILLCELL_X1 PHY_2774 ();
 FILLCELL_X1 PHY_2775 ();
 FILLCELL_X1 PHY_2776 ();
 FILLCELL_X1 PHY_2777 ();
 FILLCELL_X1 PHY_2778 ();
 FILLCELL_X1 PHY_2779 ();
 FILLCELL_X1 PHY_278 ();
 FILLCELL_X1 PHY_2780 ();
 FILLCELL_X1 PHY_2781 ();
 FILLCELL_X1 PHY_2782 ();
 FILLCELL_X1 PHY_2783 ();
 FILLCELL_X1 PHY_2784 ();
 FILLCELL_X1 PHY_2785 ();
 FILLCELL_X1 PHY_2786 ();
 FILLCELL_X1 PHY_2787 ();
 FILLCELL_X1 PHY_2788 ();
 FILLCELL_X1 PHY_2789 ();
 FILLCELL_X1 PHY_279 ();
 FILLCELL_X1 PHY_2790 ();
 FILLCELL_X1 PHY_2791 ();
 FILLCELL_X1 PHY_2792 ();
 FILLCELL_X1 PHY_2793 ();
 FILLCELL_X1 PHY_2794 ();
 FILLCELL_X1 PHY_2795 ();
 FILLCELL_X1 PHY_2796 ();
 FILLCELL_X1 PHY_2797 ();
 FILLCELL_X1 PHY_2798 ();
 FILLCELL_X1 PHY_2799 ();
 FILLCELL_X1 PHY_28 ();
 FILLCELL_X1 PHY_280 ();
 FILLCELL_X1 PHY_2800 ();
 FILLCELL_X1 PHY_2801 ();
 FILLCELL_X1 PHY_2802 ();
 FILLCELL_X1 PHY_2803 ();
 FILLCELL_X1 PHY_2804 ();
 FILLCELL_X1 PHY_2805 ();
 FILLCELL_X1 PHY_2806 ();
 FILLCELL_X1 PHY_2807 ();
 FILLCELL_X1 PHY_2808 ();
 FILLCELL_X1 PHY_2809 ();
 FILLCELL_X1 PHY_281 ();
 FILLCELL_X1 PHY_2810 ();
 FILLCELL_X1 PHY_2811 ();
 FILLCELL_X1 PHY_2812 ();
 FILLCELL_X1 PHY_2813 ();
 FILLCELL_X1 PHY_2814 ();
 FILLCELL_X1 PHY_2815 ();
 FILLCELL_X1 PHY_2816 ();
 FILLCELL_X1 PHY_2817 ();
 FILLCELL_X1 PHY_2818 ();
 FILLCELL_X1 PHY_2819 ();
 FILLCELL_X1 PHY_282 ();
 FILLCELL_X1 PHY_2820 ();
 FILLCELL_X1 PHY_2821 ();
 FILLCELL_X1 PHY_2822 ();
 FILLCELL_X1 PHY_2823 ();
 FILLCELL_X1 PHY_2824 ();
 FILLCELL_X1 PHY_2825 ();
 FILLCELL_X1 PHY_2826 ();
 FILLCELL_X1 PHY_2827 ();
 FILLCELL_X1 PHY_2828 ();
 FILLCELL_X1 PHY_2829 ();
 FILLCELL_X1 PHY_283 ();
 FILLCELL_X1 PHY_2830 ();
 FILLCELL_X1 PHY_2831 ();
 FILLCELL_X1 PHY_2832 ();
 FILLCELL_X1 PHY_2833 ();
 FILLCELL_X1 PHY_2834 ();
 FILLCELL_X1 PHY_2835 ();
 FILLCELL_X1 PHY_2836 ();
 FILLCELL_X1 PHY_2837 ();
 FILLCELL_X1 PHY_2838 ();
 FILLCELL_X1 PHY_2839 ();
 FILLCELL_X1 PHY_284 ();
 FILLCELL_X1 PHY_2840 ();
 FILLCELL_X1 PHY_2841 ();
 FILLCELL_X1 PHY_2842 ();
 FILLCELL_X1 PHY_2843 ();
 FILLCELL_X1 PHY_2844 ();
 FILLCELL_X1 PHY_2845 ();
 FILLCELL_X1 PHY_2846 ();
 FILLCELL_X1 PHY_2847 ();
 FILLCELL_X1 PHY_2848 ();
 FILLCELL_X1 PHY_2849 ();
 FILLCELL_X1 PHY_285 ();
 FILLCELL_X1 PHY_2850 ();
 FILLCELL_X1 PHY_2851 ();
 FILLCELL_X1 PHY_2852 ();
 FILLCELL_X1 PHY_2853 ();
 FILLCELL_X1 PHY_2854 ();
 FILLCELL_X1 PHY_2855 ();
 FILLCELL_X1 PHY_2856 ();
 FILLCELL_X1 PHY_2857 ();
 FILLCELL_X1 PHY_2858 ();
 FILLCELL_X1 PHY_2859 ();
 FILLCELL_X1 PHY_286 ();
 FILLCELL_X1 PHY_2860 ();
 FILLCELL_X1 PHY_2861 ();
 FILLCELL_X1 PHY_2862 ();
 FILLCELL_X1 PHY_2863 ();
 FILLCELL_X1 PHY_2864 ();
 FILLCELL_X1 PHY_2865 ();
 FILLCELL_X1 PHY_2866 ();
 FILLCELL_X1 PHY_2867 ();
 FILLCELL_X1 PHY_2868 ();
 FILLCELL_X1 PHY_2869 ();
 FILLCELL_X1 PHY_287 ();
 FILLCELL_X1 PHY_2870 ();
 FILLCELL_X1 PHY_2871 ();
 FILLCELL_X1 PHY_2872 ();
 FILLCELL_X1 PHY_2873 ();
 FILLCELL_X1 PHY_2874 ();
 FILLCELL_X1 PHY_2875 ();
 FILLCELL_X1 PHY_2876 ();
 FILLCELL_X1 PHY_2877 ();
 FILLCELL_X1 PHY_2878 ();
 FILLCELL_X1 PHY_2879 ();
 FILLCELL_X1 PHY_288 ();
 FILLCELL_X1 PHY_2880 ();
 FILLCELL_X1 PHY_2881 ();
 FILLCELL_X1 PHY_2882 ();
 FILLCELL_X1 PHY_2883 ();
 FILLCELL_X1 PHY_2884 ();
 FILLCELL_X1 PHY_2885 ();
 FILLCELL_X1 PHY_2886 ();
 FILLCELL_X1 PHY_2887 ();
 FILLCELL_X1 PHY_2888 ();
 FILLCELL_X1 PHY_2889 ();
 FILLCELL_X1 PHY_289 ();
 FILLCELL_X1 PHY_2890 ();
 FILLCELL_X1 PHY_2891 ();
 FILLCELL_X1 PHY_2892 ();
 FILLCELL_X1 PHY_2893 ();
 FILLCELL_X1 PHY_2894 ();
 FILLCELL_X1 PHY_2895 ();
 FILLCELL_X1 PHY_2896 ();
 FILLCELL_X1 PHY_2897 ();
 FILLCELL_X1 PHY_2898 ();
 FILLCELL_X1 PHY_2899 ();
 FILLCELL_X1 PHY_29 ();
 FILLCELL_X1 PHY_290 ();
 FILLCELL_X1 PHY_2900 ();
 FILLCELL_X1 PHY_2901 ();
 FILLCELL_X1 PHY_2902 ();
 FILLCELL_X1 PHY_2903 ();
 FILLCELL_X1 PHY_2904 ();
 FILLCELL_X1 PHY_2905 ();
 FILLCELL_X1 PHY_2906 ();
 FILLCELL_X1 PHY_2907 ();
 FILLCELL_X1 PHY_2908 ();
 FILLCELL_X1 PHY_2909 ();
 FILLCELL_X1 PHY_291 ();
 FILLCELL_X1 PHY_2910 ();
 FILLCELL_X1 PHY_2911 ();
 FILLCELL_X1 PHY_2912 ();
 FILLCELL_X1 PHY_2913 ();
 FILLCELL_X1 PHY_2914 ();
 FILLCELL_X1 PHY_2915 ();
 FILLCELL_X1 PHY_2916 ();
 FILLCELL_X1 PHY_2917 ();
 FILLCELL_X1 PHY_2918 ();
 FILLCELL_X1 PHY_2919 ();
 FILLCELL_X1 PHY_292 ();
 FILLCELL_X1 PHY_2920 ();
 FILLCELL_X1 PHY_2921 ();
 FILLCELL_X1 PHY_2922 ();
 FILLCELL_X1 PHY_2923 ();
 FILLCELL_X1 PHY_2924 ();
 FILLCELL_X1 PHY_2925 ();
 FILLCELL_X1 PHY_2926 ();
 FILLCELL_X1 PHY_2927 ();
 FILLCELL_X1 PHY_2928 ();
 FILLCELL_X1 PHY_2929 ();
 FILLCELL_X1 PHY_293 ();
 FILLCELL_X1 PHY_2930 ();
 FILLCELL_X1 PHY_2931 ();
 FILLCELL_X1 PHY_2932 ();
 FILLCELL_X1 PHY_2933 ();
 FILLCELL_X1 PHY_2934 ();
 FILLCELL_X1 PHY_2935 ();
 FILLCELL_X1 PHY_2936 ();
 FILLCELL_X1 PHY_2937 ();
 FILLCELL_X1 PHY_2938 ();
 FILLCELL_X1 PHY_2939 ();
 FILLCELL_X1 PHY_294 ();
 FILLCELL_X1 PHY_2940 ();
 FILLCELL_X1 PHY_2941 ();
 FILLCELL_X1 PHY_2942 ();
 FILLCELL_X1 PHY_2943 ();
 FILLCELL_X1 PHY_2944 ();
 FILLCELL_X1 PHY_2945 ();
 FILLCELL_X1 PHY_2946 ();
 FILLCELL_X1 PHY_2947 ();
 FILLCELL_X1 PHY_2948 ();
 FILLCELL_X1 PHY_2949 ();
 FILLCELL_X1 PHY_295 ();
 FILLCELL_X1 PHY_2950 ();
 FILLCELL_X1 PHY_2951 ();
 FILLCELL_X1 PHY_2952 ();
 FILLCELL_X1 PHY_2953 ();
 FILLCELL_X1 PHY_2954 ();
 FILLCELL_X1 PHY_2955 ();
 FILLCELL_X1 PHY_2956 ();
 FILLCELL_X1 PHY_2957 ();
 FILLCELL_X1 PHY_2958 ();
 FILLCELL_X1 PHY_2959 ();
 FILLCELL_X1 PHY_296 ();
 FILLCELL_X1 PHY_2960 ();
 FILLCELL_X1 PHY_2961 ();
 FILLCELL_X1 PHY_2962 ();
 FILLCELL_X1 PHY_2963 ();
 FILLCELL_X1 PHY_2964 ();
 FILLCELL_X1 PHY_2965 ();
 FILLCELL_X1 PHY_2966 ();
 FILLCELL_X1 PHY_2967 ();
 FILLCELL_X1 PHY_2968 ();
 FILLCELL_X1 PHY_2969 ();
 FILLCELL_X1 PHY_297 ();
 FILLCELL_X1 PHY_2970 ();
 FILLCELL_X1 PHY_2971 ();
 FILLCELL_X1 PHY_2972 ();
 FILLCELL_X1 PHY_2973 ();
 FILLCELL_X1 PHY_2974 ();
 FILLCELL_X1 PHY_2975 ();
 FILLCELL_X1 PHY_2976 ();
 FILLCELL_X1 PHY_2977 ();
 FILLCELL_X1 PHY_2978 ();
 FILLCELL_X1 PHY_2979 ();
 FILLCELL_X1 PHY_298 ();
 FILLCELL_X1 PHY_2980 ();
 FILLCELL_X1 PHY_2981 ();
 FILLCELL_X1 PHY_2982 ();
 FILLCELL_X1 PHY_2983 ();
 FILLCELL_X1 PHY_2984 ();
 FILLCELL_X1 PHY_2985 ();
 FILLCELL_X1 PHY_2986 ();
 FILLCELL_X1 PHY_2987 ();
 FILLCELL_X1 PHY_2988 ();
 FILLCELL_X1 PHY_2989 ();
 FILLCELL_X1 PHY_299 ();
 FILLCELL_X1 PHY_2990 ();
 FILLCELL_X1 PHY_2991 ();
 FILLCELL_X1 PHY_2992 ();
 FILLCELL_X1 PHY_2993 ();
 FILLCELL_X1 PHY_2994 ();
 FILLCELL_X1 PHY_2995 ();
 FILLCELL_X1 PHY_2996 ();
 FILLCELL_X1 PHY_2997 ();
 FILLCELL_X1 PHY_2998 ();
 FILLCELL_X1 PHY_2999 ();
 FILLCELL_X1 PHY_3 ();
 FILLCELL_X1 PHY_30 ();
 FILLCELL_X1 PHY_300 ();
 FILLCELL_X1 PHY_3000 ();
 FILLCELL_X1 PHY_3001 ();
 FILLCELL_X1 PHY_3002 ();
 FILLCELL_X1 PHY_3003 ();
 FILLCELL_X1 PHY_3004 ();
 FILLCELL_X1 PHY_3005 ();
 FILLCELL_X1 PHY_3006 ();
 FILLCELL_X1 PHY_3007 ();
 FILLCELL_X1 PHY_3008 ();
 FILLCELL_X1 PHY_3009 ();
 FILLCELL_X1 PHY_301 ();
 FILLCELL_X1 PHY_3010 ();
 FILLCELL_X1 PHY_3011 ();
 FILLCELL_X1 PHY_3012 ();
 FILLCELL_X1 PHY_3013 ();
 FILLCELL_X1 PHY_3014 ();
 FILLCELL_X1 PHY_3015 ();
 FILLCELL_X1 PHY_3016 ();
 FILLCELL_X1 PHY_3017 ();
 FILLCELL_X1 PHY_3018 ();
 FILLCELL_X1 PHY_3019 ();
 FILLCELL_X1 PHY_302 ();
 FILLCELL_X1 PHY_3020 ();
 FILLCELL_X1 PHY_3021 ();
 FILLCELL_X1 PHY_3022 ();
 FILLCELL_X1 PHY_3023 ();
 FILLCELL_X1 PHY_3024 ();
 FILLCELL_X1 PHY_3025 ();
 FILLCELL_X1 PHY_3026 ();
 FILLCELL_X1 PHY_3027 ();
 FILLCELL_X1 PHY_3028 ();
 FILLCELL_X1 PHY_3029 ();
 FILLCELL_X1 PHY_303 ();
 FILLCELL_X1 PHY_3030 ();
 FILLCELL_X1 PHY_3031 ();
 FILLCELL_X1 PHY_3032 ();
 FILLCELL_X1 PHY_3033 ();
 FILLCELL_X1 PHY_3034 ();
 FILLCELL_X1 PHY_3035 ();
 FILLCELL_X1 PHY_3036 ();
 FILLCELL_X1 PHY_3037 ();
 FILLCELL_X1 PHY_3038 ();
 FILLCELL_X1 PHY_3039 ();
 FILLCELL_X1 PHY_304 ();
 FILLCELL_X1 PHY_3040 ();
 FILLCELL_X1 PHY_3041 ();
 FILLCELL_X1 PHY_3042 ();
 FILLCELL_X1 PHY_3043 ();
 FILLCELL_X1 PHY_3044 ();
 FILLCELL_X1 PHY_3045 ();
 FILLCELL_X1 PHY_3046 ();
 FILLCELL_X1 PHY_3047 ();
 FILLCELL_X1 PHY_3048 ();
 FILLCELL_X1 PHY_3049 ();
 FILLCELL_X1 PHY_305 ();
 FILLCELL_X1 PHY_3050 ();
 FILLCELL_X1 PHY_3051 ();
 FILLCELL_X1 PHY_3052 ();
 FILLCELL_X1 PHY_3053 ();
 FILLCELL_X1 PHY_3054 ();
 FILLCELL_X1 PHY_3055 ();
 FILLCELL_X1 PHY_3056 ();
 FILLCELL_X1 PHY_3057 ();
 FILLCELL_X1 PHY_3058 ();
 FILLCELL_X1 PHY_3059 ();
 FILLCELL_X1 PHY_306 ();
 FILLCELL_X1 PHY_3060 ();
 FILLCELL_X1 PHY_3061 ();
 FILLCELL_X1 PHY_3062 ();
 FILLCELL_X1 PHY_3063 ();
 FILLCELL_X1 PHY_3064 ();
 FILLCELL_X1 PHY_3065 ();
 FILLCELL_X1 PHY_3066 ();
 FILLCELL_X1 PHY_3067 ();
 FILLCELL_X1 PHY_3068 ();
 FILLCELL_X1 PHY_3069 ();
 FILLCELL_X1 PHY_307 ();
 FILLCELL_X1 PHY_3070 ();
 FILLCELL_X1 PHY_3071 ();
 FILLCELL_X1 PHY_3072 ();
 FILLCELL_X1 PHY_3073 ();
 FILLCELL_X1 PHY_3074 ();
 FILLCELL_X1 PHY_3075 ();
 FILLCELL_X1 PHY_3076 ();
 FILLCELL_X1 PHY_3077 ();
 FILLCELL_X1 PHY_3078 ();
 FILLCELL_X1 PHY_3079 ();
 FILLCELL_X1 PHY_308 ();
 FILLCELL_X1 PHY_3080 ();
 FILLCELL_X1 PHY_3081 ();
 FILLCELL_X1 PHY_3082 ();
 FILLCELL_X1 PHY_3083 ();
 FILLCELL_X1 PHY_3084 ();
 FILLCELL_X1 PHY_3085 ();
 FILLCELL_X1 PHY_3086 ();
 FILLCELL_X1 PHY_3087 ();
 FILLCELL_X1 PHY_3088 ();
 FILLCELL_X1 PHY_3089 ();
 FILLCELL_X1 PHY_309 ();
 FILLCELL_X1 PHY_3090 ();
 FILLCELL_X1 PHY_3091 ();
 FILLCELL_X1 PHY_3092 ();
 FILLCELL_X1 PHY_3093 ();
 FILLCELL_X1 PHY_3094 ();
 FILLCELL_X1 PHY_3095 ();
 FILLCELL_X1 PHY_3096 ();
 FILLCELL_X1 PHY_3097 ();
 FILLCELL_X1 PHY_3098 ();
 FILLCELL_X1 PHY_3099 ();
 FILLCELL_X1 PHY_31 ();
 FILLCELL_X1 PHY_310 ();
 FILLCELL_X1 PHY_3100 ();
 FILLCELL_X1 PHY_3101 ();
 FILLCELL_X1 PHY_3102 ();
 FILLCELL_X1 PHY_3103 ();
 FILLCELL_X1 PHY_3104 ();
 FILLCELL_X1 PHY_3105 ();
 FILLCELL_X1 PHY_3106 ();
 FILLCELL_X1 PHY_3107 ();
 FILLCELL_X1 PHY_3108 ();
 FILLCELL_X1 PHY_3109 ();
 FILLCELL_X1 PHY_311 ();
 FILLCELL_X1 PHY_3110 ();
 FILLCELL_X1 PHY_3111 ();
 FILLCELL_X1 PHY_3112 ();
 FILLCELL_X1 PHY_3113 ();
 FILLCELL_X1 PHY_3114 ();
 FILLCELL_X1 PHY_3115 ();
 FILLCELL_X1 PHY_3116 ();
 FILLCELL_X1 PHY_3117 ();
 FILLCELL_X1 PHY_3118 ();
 FILLCELL_X1 PHY_3119 ();
 FILLCELL_X1 PHY_312 ();
 FILLCELL_X1 PHY_3120 ();
 FILLCELL_X1 PHY_3121 ();
 FILLCELL_X1 PHY_3122 ();
 FILLCELL_X1 PHY_3123 ();
 FILLCELL_X1 PHY_3124 ();
 FILLCELL_X1 PHY_3125 ();
 FILLCELL_X1 PHY_3126 ();
 FILLCELL_X1 PHY_3127 ();
 FILLCELL_X1 PHY_3128 ();
 FILLCELL_X1 PHY_3129 ();
 FILLCELL_X1 PHY_313 ();
 FILLCELL_X1 PHY_3130 ();
 FILLCELL_X1 PHY_3131 ();
 FILLCELL_X1 PHY_3132 ();
 FILLCELL_X1 PHY_3133 ();
 FILLCELL_X1 PHY_3134 ();
 FILLCELL_X1 PHY_3135 ();
 FILLCELL_X1 PHY_3136 ();
 FILLCELL_X1 PHY_3137 ();
 FILLCELL_X1 PHY_3138 ();
 FILLCELL_X1 PHY_3139 ();
 FILLCELL_X1 PHY_314 ();
 FILLCELL_X1 PHY_3140 ();
 FILLCELL_X1 PHY_3141 ();
 FILLCELL_X1 PHY_3142 ();
 FILLCELL_X1 PHY_3143 ();
 FILLCELL_X1 PHY_3144 ();
 FILLCELL_X1 PHY_3145 ();
 FILLCELL_X1 PHY_3146 ();
 FILLCELL_X1 PHY_3147 ();
 FILLCELL_X1 PHY_3148 ();
 FILLCELL_X1 PHY_3149 ();
 FILLCELL_X1 PHY_315 ();
 FILLCELL_X1 PHY_3150 ();
 FILLCELL_X1 PHY_3151 ();
 FILLCELL_X1 PHY_3152 ();
 FILLCELL_X1 PHY_3153 ();
 FILLCELL_X1 PHY_3154 ();
 FILLCELL_X1 PHY_3155 ();
 FILLCELL_X1 PHY_3156 ();
 FILLCELL_X1 PHY_3157 ();
 FILLCELL_X1 PHY_3158 ();
 FILLCELL_X1 PHY_3159 ();
 FILLCELL_X1 PHY_316 ();
 FILLCELL_X1 PHY_3160 ();
 FILLCELL_X1 PHY_3161 ();
 FILLCELL_X1 PHY_3162 ();
 FILLCELL_X1 PHY_3163 ();
 FILLCELL_X1 PHY_3164 ();
 FILLCELL_X1 PHY_3165 ();
 FILLCELL_X1 PHY_3166 ();
 FILLCELL_X1 PHY_3167 ();
 FILLCELL_X1 PHY_3168 ();
 FILLCELL_X1 PHY_3169 ();
 FILLCELL_X1 PHY_317 ();
 FILLCELL_X1 PHY_3170 ();
 FILLCELL_X1 PHY_3171 ();
 FILLCELL_X1 PHY_3172 ();
 FILLCELL_X1 PHY_3173 ();
 FILLCELL_X1 PHY_3174 ();
 FILLCELL_X1 PHY_3175 ();
 FILLCELL_X1 PHY_3176 ();
 FILLCELL_X1 PHY_3177 ();
 FILLCELL_X1 PHY_3178 ();
 FILLCELL_X1 PHY_3179 ();
 FILLCELL_X1 PHY_318 ();
 FILLCELL_X1 PHY_3180 ();
 FILLCELL_X1 PHY_3181 ();
 FILLCELL_X1 PHY_3182 ();
 FILLCELL_X1 PHY_3183 ();
 FILLCELL_X1 PHY_3184 ();
 FILLCELL_X1 PHY_3185 ();
 FILLCELL_X1 PHY_3186 ();
 FILLCELL_X1 PHY_3187 ();
 FILLCELL_X1 PHY_3188 ();
 FILLCELL_X1 PHY_3189 ();
 FILLCELL_X1 PHY_319 ();
 FILLCELL_X1 PHY_3190 ();
 FILLCELL_X1 PHY_3191 ();
 FILLCELL_X1 PHY_3192 ();
 FILLCELL_X1 PHY_3193 ();
 FILLCELL_X1 PHY_3194 ();
 FILLCELL_X1 PHY_3195 ();
 FILLCELL_X1 PHY_3196 ();
 FILLCELL_X1 PHY_3197 ();
 FILLCELL_X1 PHY_3198 ();
 FILLCELL_X1 PHY_3199 ();
 FILLCELL_X1 PHY_32 ();
 FILLCELL_X1 PHY_320 ();
 FILLCELL_X1 PHY_3200 ();
 FILLCELL_X1 PHY_3201 ();
 FILLCELL_X1 PHY_3202 ();
 FILLCELL_X1 PHY_3203 ();
 FILLCELL_X1 PHY_3204 ();
 FILLCELL_X1 PHY_3205 ();
 FILLCELL_X1 PHY_3206 ();
 FILLCELL_X1 PHY_3207 ();
 FILLCELL_X1 PHY_3208 ();
 FILLCELL_X1 PHY_3209 ();
 FILLCELL_X1 PHY_321 ();
 FILLCELL_X1 PHY_3210 ();
 FILLCELL_X1 PHY_3211 ();
 FILLCELL_X1 PHY_3212 ();
 FILLCELL_X1 PHY_3213 ();
 FILLCELL_X1 PHY_3214 ();
 FILLCELL_X1 PHY_3215 ();
 FILLCELL_X1 PHY_3216 ();
 FILLCELL_X1 PHY_3217 ();
 FILLCELL_X1 PHY_3218 ();
 FILLCELL_X1 PHY_3219 ();
 FILLCELL_X1 PHY_322 ();
 FILLCELL_X1 PHY_3220 ();
 FILLCELL_X1 PHY_3221 ();
 FILLCELL_X1 PHY_3222 ();
 FILLCELL_X1 PHY_3223 ();
 FILLCELL_X1 PHY_3224 ();
 FILLCELL_X1 PHY_3225 ();
 FILLCELL_X1 PHY_3226 ();
 FILLCELL_X1 PHY_3227 ();
 FILLCELL_X1 PHY_3228 ();
 FILLCELL_X1 PHY_3229 ();
 FILLCELL_X1 PHY_323 ();
 FILLCELL_X1 PHY_3230 ();
 FILLCELL_X1 PHY_3231 ();
 FILLCELL_X1 PHY_3232 ();
 FILLCELL_X1 PHY_3233 ();
 FILLCELL_X1 PHY_3234 ();
 FILLCELL_X1 PHY_3235 ();
 FILLCELL_X1 PHY_3236 ();
 FILLCELL_X1 PHY_3237 ();
 FILLCELL_X1 PHY_3238 ();
 FILLCELL_X1 PHY_3239 ();
 FILLCELL_X1 PHY_324 ();
 FILLCELL_X1 PHY_3240 ();
 FILLCELL_X1 PHY_3241 ();
 FILLCELL_X1 PHY_3242 ();
 FILLCELL_X1 PHY_3243 ();
 FILLCELL_X1 PHY_3244 ();
 FILLCELL_X1 PHY_3245 ();
 FILLCELL_X1 PHY_3246 ();
 FILLCELL_X1 PHY_3247 ();
 FILLCELL_X1 PHY_3248 ();
 FILLCELL_X1 PHY_3249 ();
 FILLCELL_X1 PHY_325 ();
 FILLCELL_X1 PHY_3250 ();
 FILLCELL_X1 PHY_3251 ();
 FILLCELL_X1 PHY_3252 ();
 FILLCELL_X1 PHY_3253 ();
 FILLCELL_X1 PHY_3254 ();
 FILLCELL_X1 PHY_3255 ();
 FILLCELL_X1 PHY_3256 ();
 FILLCELL_X1 PHY_3257 ();
 FILLCELL_X1 PHY_3258 ();
 FILLCELL_X1 PHY_3259 ();
 FILLCELL_X1 PHY_326 ();
 FILLCELL_X1 PHY_3260 ();
 FILLCELL_X1 PHY_3261 ();
 FILLCELL_X1 PHY_3262 ();
 FILLCELL_X1 PHY_3263 ();
 FILLCELL_X1 PHY_3264 ();
 FILLCELL_X1 PHY_3265 ();
 FILLCELL_X1 PHY_3266 ();
 FILLCELL_X1 PHY_3267 ();
 FILLCELL_X1 PHY_3268 ();
 FILLCELL_X1 PHY_3269 ();
 FILLCELL_X1 PHY_327 ();
 FILLCELL_X1 PHY_3270 ();
 FILLCELL_X1 PHY_3271 ();
 FILLCELL_X1 PHY_3272 ();
 FILLCELL_X1 PHY_3273 ();
 FILLCELL_X1 PHY_3274 ();
 FILLCELL_X1 PHY_3275 ();
 FILLCELL_X1 PHY_3276 ();
 FILLCELL_X1 PHY_3277 ();
 FILLCELL_X1 PHY_3278 ();
 FILLCELL_X1 PHY_3279 ();
 FILLCELL_X1 PHY_328 ();
 FILLCELL_X1 PHY_3280 ();
 FILLCELL_X1 PHY_3281 ();
 FILLCELL_X1 PHY_3282 ();
 FILLCELL_X1 PHY_3283 ();
 FILLCELL_X1 PHY_3284 ();
 FILLCELL_X1 PHY_3285 ();
 FILLCELL_X1 PHY_3286 ();
 FILLCELL_X1 PHY_3287 ();
 FILLCELL_X1 PHY_3288 ();
 FILLCELL_X1 PHY_3289 ();
 FILLCELL_X1 PHY_329 ();
 FILLCELL_X1 PHY_3290 ();
 FILLCELL_X1 PHY_3291 ();
 FILLCELL_X1 PHY_3292 ();
 FILLCELL_X1 PHY_3293 ();
 FILLCELL_X1 PHY_3294 ();
 FILLCELL_X1 PHY_3295 ();
 FILLCELL_X1 PHY_3296 ();
 FILLCELL_X1 PHY_3297 ();
 FILLCELL_X1 PHY_3298 ();
 FILLCELL_X1 PHY_3299 ();
 FILLCELL_X1 PHY_33 ();
 FILLCELL_X1 PHY_330 ();
 FILLCELL_X1 PHY_3300 ();
 FILLCELL_X1 PHY_3301 ();
 FILLCELL_X1 PHY_3302 ();
 FILLCELL_X1 PHY_3303 ();
 FILLCELL_X1 PHY_3304 ();
 FILLCELL_X1 PHY_3305 ();
 FILLCELL_X1 PHY_3306 ();
 FILLCELL_X1 PHY_3307 ();
 FILLCELL_X1 PHY_3308 ();
 FILLCELL_X1 PHY_3309 ();
 FILLCELL_X1 PHY_331 ();
 FILLCELL_X1 PHY_3310 ();
 FILLCELL_X1 PHY_3311 ();
 FILLCELL_X1 PHY_3312 ();
 FILLCELL_X1 PHY_3313 ();
 FILLCELL_X1 PHY_3314 ();
 FILLCELL_X1 PHY_3315 ();
 FILLCELL_X1 PHY_3316 ();
 FILLCELL_X1 PHY_3317 ();
 FILLCELL_X1 PHY_3318 ();
 FILLCELL_X1 PHY_3319 ();
 FILLCELL_X1 PHY_332 ();
 FILLCELL_X1 PHY_3320 ();
 FILLCELL_X1 PHY_3321 ();
 FILLCELL_X1 PHY_3322 ();
 FILLCELL_X1 PHY_3323 ();
 FILLCELL_X1 PHY_3324 ();
 FILLCELL_X1 PHY_3325 ();
 FILLCELL_X1 PHY_3326 ();
 FILLCELL_X1 PHY_3327 ();
 FILLCELL_X1 PHY_3328 ();
 FILLCELL_X1 PHY_3329 ();
 FILLCELL_X1 PHY_333 ();
 FILLCELL_X1 PHY_3330 ();
 FILLCELL_X1 PHY_3331 ();
 FILLCELL_X1 PHY_3332 ();
 FILLCELL_X1 PHY_3333 ();
 FILLCELL_X1 PHY_3334 ();
 FILLCELL_X1 PHY_3335 ();
 FILLCELL_X1 PHY_3336 ();
 FILLCELL_X1 PHY_3337 ();
 FILLCELL_X1 PHY_3338 ();
 FILLCELL_X1 PHY_3339 ();
 FILLCELL_X1 PHY_334 ();
 FILLCELL_X1 PHY_3340 ();
 FILLCELL_X1 PHY_3341 ();
 FILLCELL_X1 PHY_3342 ();
 FILLCELL_X1 PHY_3343 ();
 FILLCELL_X1 PHY_3344 ();
 FILLCELL_X1 PHY_3345 ();
 FILLCELL_X1 PHY_3346 ();
 FILLCELL_X1 PHY_3347 ();
 FILLCELL_X1 PHY_3348 ();
 FILLCELL_X1 PHY_3349 ();
 FILLCELL_X1 PHY_335 ();
 FILLCELL_X1 PHY_3350 ();
 FILLCELL_X1 PHY_3351 ();
 FILLCELL_X1 PHY_3352 ();
 FILLCELL_X1 PHY_3353 ();
 FILLCELL_X1 PHY_3354 ();
 FILLCELL_X1 PHY_3355 ();
 FILLCELL_X1 PHY_3356 ();
 FILLCELL_X1 PHY_3357 ();
 FILLCELL_X1 PHY_3358 ();
 FILLCELL_X1 PHY_3359 ();
 FILLCELL_X1 PHY_336 ();
 FILLCELL_X1 PHY_3360 ();
 FILLCELL_X1 PHY_3361 ();
 FILLCELL_X1 PHY_3362 ();
 FILLCELL_X1 PHY_3363 ();
 FILLCELL_X1 PHY_3364 ();
 FILLCELL_X1 PHY_3365 ();
 FILLCELL_X1 PHY_3366 ();
 FILLCELL_X1 PHY_3367 ();
 FILLCELL_X1 PHY_3368 ();
 FILLCELL_X1 PHY_3369 ();
 FILLCELL_X1 PHY_337 ();
 FILLCELL_X1 PHY_3370 ();
 FILLCELL_X1 PHY_3371 ();
 FILLCELL_X1 PHY_3372 ();
 FILLCELL_X1 PHY_3373 ();
 FILLCELL_X1 PHY_3374 ();
 FILLCELL_X1 PHY_3375 ();
 FILLCELL_X1 PHY_3376 ();
 FILLCELL_X1 PHY_3377 ();
 FILLCELL_X1 PHY_3378 ();
 FILLCELL_X1 PHY_3379 ();
 FILLCELL_X1 PHY_338 ();
 FILLCELL_X1 PHY_3380 ();
 FILLCELL_X1 PHY_3381 ();
 FILLCELL_X1 PHY_3382 ();
 FILLCELL_X1 PHY_3383 ();
 FILLCELL_X1 PHY_3384 ();
 FILLCELL_X1 PHY_3385 ();
 FILLCELL_X1 PHY_3386 ();
 FILLCELL_X1 PHY_3387 ();
 FILLCELL_X1 PHY_3388 ();
 FILLCELL_X1 PHY_3389 ();
 FILLCELL_X1 PHY_339 ();
 FILLCELL_X1 PHY_3390 ();
 FILLCELL_X1 PHY_3391 ();
 FILLCELL_X1 PHY_3392 ();
 FILLCELL_X1 PHY_3393 ();
 FILLCELL_X1 PHY_3394 ();
 FILLCELL_X1 PHY_3395 ();
 FILLCELL_X1 PHY_3396 ();
 FILLCELL_X1 PHY_3397 ();
 FILLCELL_X1 PHY_3398 ();
 FILLCELL_X1 PHY_3399 ();
 FILLCELL_X1 PHY_34 ();
 FILLCELL_X1 PHY_340 ();
 FILLCELL_X1 PHY_3400 ();
 FILLCELL_X1 PHY_3401 ();
 FILLCELL_X1 PHY_3402 ();
 FILLCELL_X1 PHY_3403 ();
 FILLCELL_X1 PHY_3404 ();
 FILLCELL_X1 PHY_3405 ();
 FILLCELL_X1 PHY_3406 ();
 FILLCELL_X1 PHY_3407 ();
 FILLCELL_X1 PHY_3408 ();
 FILLCELL_X1 PHY_3409 ();
 FILLCELL_X1 PHY_341 ();
 FILLCELL_X1 PHY_3410 ();
 FILLCELL_X1 PHY_3411 ();
 FILLCELL_X1 PHY_3412 ();
 FILLCELL_X1 PHY_3413 ();
 FILLCELL_X1 PHY_3414 ();
 FILLCELL_X1 PHY_3415 ();
 FILLCELL_X1 PHY_3416 ();
 FILLCELL_X1 PHY_3417 ();
 FILLCELL_X1 PHY_3418 ();
 FILLCELL_X1 PHY_3419 ();
 FILLCELL_X1 PHY_342 ();
 FILLCELL_X1 PHY_3420 ();
 FILLCELL_X1 PHY_3421 ();
 FILLCELL_X1 PHY_3422 ();
 FILLCELL_X1 PHY_3423 ();
 FILLCELL_X1 PHY_3424 ();
 FILLCELL_X1 PHY_3425 ();
 FILLCELL_X1 PHY_3426 ();
 FILLCELL_X1 PHY_3427 ();
 FILLCELL_X1 PHY_3428 ();
 FILLCELL_X1 PHY_3429 ();
 FILLCELL_X1 PHY_343 ();
 FILLCELL_X1 PHY_3430 ();
 FILLCELL_X1 PHY_3431 ();
 FILLCELL_X1 PHY_3432 ();
 FILLCELL_X1 PHY_3433 ();
 FILLCELL_X1 PHY_3434 ();
 FILLCELL_X1 PHY_3435 ();
 FILLCELL_X1 PHY_3436 ();
 FILLCELL_X1 PHY_3437 ();
 FILLCELL_X1 PHY_3438 ();
 FILLCELL_X1 PHY_3439 ();
 FILLCELL_X1 PHY_344 ();
 FILLCELL_X1 PHY_3440 ();
 FILLCELL_X1 PHY_3441 ();
 FILLCELL_X1 PHY_3442 ();
 FILLCELL_X1 PHY_3443 ();
 FILLCELL_X1 PHY_3444 ();
 FILLCELL_X1 PHY_3445 ();
 FILLCELL_X1 PHY_3446 ();
 FILLCELL_X1 PHY_3447 ();
 FILLCELL_X1 PHY_3448 ();
 FILLCELL_X1 PHY_3449 ();
 FILLCELL_X1 PHY_345 ();
 FILLCELL_X1 PHY_3450 ();
 FILLCELL_X1 PHY_3451 ();
 FILLCELL_X1 PHY_3452 ();
 FILLCELL_X1 PHY_3453 ();
 FILLCELL_X1 PHY_3454 ();
 FILLCELL_X1 PHY_3455 ();
 FILLCELL_X1 PHY_3456 ();
 FILLCELL_X1 PHY_3457 ();
 FILLCELL_X1 PHY_3458 ();
 FILLCELL_X1 PHY_3459 ();
 FILLCELL_X1 PHY_346 ();
 FILLCELL_X1 PHY_3460 ();
 FILLCELL_X1 PHY_3461 ();
 FILLCELL_X1 PHY_3462 ();
 FILLCELL_X1 PHY_3463 ();
 FILLCELL_X1 PHY_3464 ();
 FILLCELL_X1 PHY_3465 ();
 FILLCELL_X1 PHY_3466 ();
 FILLCELL_X1 PHY_3467 ();
 FILLCELL_X1 PHY_3468 ();
 FILLCELL_X1 PHY_3469 ();
 FILLCELL_X1 PHY_347 ();
 FILLCELL_X1 PHY_3470 ();
 FILLCELL_X1 PHY_3471 ();
 FILLCELL_X1 PHY_3472 ();
 FILLCELL_X1 PHY_3473 ();
 FILLCELL_X1 PHY_3474 ();
 FILLCELL_X1 PHY_3475 ();
 FILLCELL_X1 PHY_3476 ();
 FILLCELL_X1 PHY_3477 ();
 FILLCELL_X1 PHY_3478 ();
 FILLCELL_X1 PHY_3479 ();
 FILLCELL_X1 PHY_348 ();
 FILLCELL_X1 PHY_3480 ();
 FILLCELL_X1 PHY_3481 ();
 FILLCELL_X1 PHY_3482 ();
 FILLCELL_X1 PHY_3483 ();
 FILLCELL_X1 PHY_3484 ();
 FILLCELL_X1 PHY_3485 ();
 FILLCELL_X1 PHY_3486 ();
 FILLCELL_X1 PHY_3487 ();
 FILLCELL_X1 PHY_3488 ();
 FILLCELL_X1 PHY_3489 ();
 FILLCELL_X1 PHY_349 ();
 FILLCELL_X1 PHY_3490 ();
 FILLCELL_X1 PHY_3491 ();
 FILLCELL_X1 PHY_3492 ();
 FILLCELL_X1 PHY_3493 ();
 FILLCELL_X1 PHY_3494 ();
 FILLCELL_X1 PHY_3495 ();
 FILLCELL_X1 PHY_3496 ();
 FILLCELL_X1 PHY_3497 ();
 FILLCELL_X1 PHY_3498 ();
 FILLCELL_X1 PHY_3499 ();
 FILLCELL_X1 PHY_35 ();
 FILLCELL_X1 PHY_350 ();
 FILLCELL_X1 PHY_3500 ();
 FILLCELL_X1 PHY_3501 ();
 FILLCELL_X1 PHY_3502 ();
 FILLCELL_X1 PHY_3503 ();
 FILLCELL_X1 PHY_3504 ();
 FILLCELL_X1 PHY_3505 ();
 FILLCELL_X1 PHY_3506 ();
 FILLCELL_X1 PHY_3507 ();
 FILLCELL_X1 PHY_3508 ();
 FILLCELL_X1 PHY_3509 ();
 FILLCELL_X1 PHY_351 ();
 FILLCELL_X1 PHY_3510 ();
 FILLCELL_X1 PHY_3511 ();
 FILLCELL_X1 PHY_3512 ();
 FILLCELL_X1 PHY_3513 ();
 FILLCELL_X1 PHY_3514 ();
 FILLCELL_X1 PHY_3515 ();
 FILLCELL_X1 PHY_3516 ();
 FILLCELL_X1 PHY_3517 ();
 FILLCELL_X1 PHY_3518 ();
 FILLCELL_X1 PHY_3519 ();
 FILLCELL_X1 PHY_352 ();
 FILLCELL_X1 PHY_3520 ();
 FILLCELL_X1 PHY_3521 ();
 FILLCELL_X1 PHY_3522 ();
 FILLCELL_X1 PHY_3523 ();
 FILLCELL_X1 PHY_3524 ();
 FILLCELL_X1 PHY_3525 ();
 FILLCELL_X1 PHY_3526 ();
 FILLCELL_X1 PHY_3527 ();
 FILLCELL_X1 PHY_3528 ();
 FILLCELL_X1 PHY_3529 ();
 FILLCELL_X1 PHY_353 ();
 FILLCELL_X1 PHY_3530 ();
 FILLCELL_X1 PHY_3531 ();
 FILLCELL_X1 PHY_3532 ();
 FILLCELL_X1 PHY_3533 ();
 FILLCELL_X1 PHY_3534 ();
 FILLCELL_X1 PHY_3535 ();
 FILLCELL_X1 PHY_3536 ();
 FILLCELL_X1 PHY_3537 ();
 FILLCELL_X1 PHY_3538 ();
 FILLCELL_X1 PHY_3539 ();
 FILLCELL_X1 PHY_354 ();
 FILLCELL_X1 PHY_3540 ();
 FILLCELL_X1 PHY_3541 ();
 FILLCELL_X1 PHY_3542 ();
 FILLCELL_X1 PHY_3543 ();
 FILLCELL_X1 PHY_3544 ();
 FILLCELL_X1 PHY_3545 ();
 FILLCELL_X1 PHY_3546 ();
 FILLCELL_X1 PHY_3547 ();
 FILLCELL_X1 PHY_3548 ();
 FILLCELL_X1 PHY_3549 ();
 FILLCELL_X1 PHY_355 ();
 FILLCELL_X1 PHY_3550 ();
 FILLCELL_X1 PHY_3551 ();
 FILLCELL_X1 PHY_3552 ();
 FILLCELL_X1 PHY_3553 ();
 FILLCELL_X1 PHY_3554 ();
 FILLCELL_X1 PHY_3555 ();
 FILLCELL_X1 PHY_3556 ();
 FILLCELL_X1 PHY_3557 ();
 FILLCELL_X1 PHY_3558 ();
 FILLCELL_X1 PHY_3559 ();
 FILLCELL_X1 PHY_356 ();
 FILLCELL_X1 PHY_3560 ();
 FILLCELL_X1 PHY_3561 ();
 FILLCELL_X1 PHY_3562 ();
 FILLCELL_X1 PHY_3563 ();
 FILLCELL_X1 PHY_3564 ();
 FILLCELL_X1 PHY_3565 ();
 FILLCELL_X1 PHY_3566 ();
 FILLCELL_X1 PHY_3567 ();
 FILLCELL_X1 PHY_3568 ();
 FILLCELL_X1 PHY_3569 ();
 FILLCELL_X1 PHY_357 ();
 FILLCELL_X1 PHY_3570 ();
 FILLCELL_X1 PHY_3571 ();
 FILLCELL_X1 PHY_3572 ();
 FILLCELL_X1 PHY_3573 ();
 FILLCELL_X1 PHY_3574 ();
 FILLCELL_X1 PHY_3575 ();
 FILLCELL_X1 PHY_3576 ();
 FILLCELL_X1 PHY_3577 ();
 FILLCELL_X1 PHY_3578 ();
 FILLCELL_X1 PHY_3579 ();
 FILLCELL_X1 PHY_358 ();
 FILLCELL_X1 PHY_3580 ();
 FILLCELL_X1 PHY_3581 ();
 FILLCELL_X1 PHY_3582 ();
 FILLCELL_X1 PHY_3583 ();
 FILLCELL_X1 PHY_3584 ();
 FILLCELL_X1 PHY_3585 ();
 FILLCELL_X1 PHY_3586 ();
 FILLCELL_X1 PHY_3587 ();
 FILLCELL_X1 PHY_3588 ();
 FILLCELL_X1 PHY_3589 ();
 FILLCELL_X1 PHY_359 ();
 FILLCELL_X1 PHY_3590 ();
 FILLCELL_X1 PHY_3591 ();
 FILLCELL_X1 PHY_3592 ();
 FILLCELL_X1 PHY_3593 ();
 FILLCELL_X1 PHY_3594 ();
 FILLCELL_X1 PHY_3595 ();
 FILLCELL_X1 PHY_3596 ();
 FILLCELL_X1 PHY_3597 ();
 FILLCELL_X1 PHY_3598 ();
 FILLCELL_X1 PHY_3599 ();
 FILLCELL_X1 PHY_36 ();
 FILLCELL_X1 PHY_360 ();
 FILLCELL_X1 PHY_3600 ();
 FILLCELL_X1 PHY_3601 ();
 FILLCELL_X1 PHY_3602 ();
 FILLCELL_X1 PHY_3603 ();
 FILLCELL_X1 PHY_3604 ();
 FILLCELL_X1 PHY_3605 ();
 FILLCELL_X1 PHY_3606 ();
 FILLCELL_X1 PHY_3607 ();
 FILLCELL_X1 PHY_3608 ();
 FILLCELL_X1 PHY_3609 ();
 FILLCELL_X1 PHY_361 ();
 FILLCELL_X1 PHY_3610 ();
 FILLCELL_X1 PHY_3611 ();
 FILLCELL_X1 PHY_3612 ();
 FILLCELL_X1 PHY_3613 ();
 FILLCELL_X1 PHY_3614 ();
 FILLCELL_X1 PHY_3615 ();
 FILLCELL_X1 PHY_3616 ();
 FILLCELL_X1 PHY_3617 ();
 FILLCELL_X1 PHY_3618 ();
 FILLCELL_X1 PHY_3619 ();
 FILLCELL_X1 PHY_362 ();
 FILLCELL_X1 PHY_3620 ();
 FILLCELL_X1 PHY_3621 ();
 FILLCELL_X1 PHY_3622 ();
 FILLCELL_X1 PHY_3623 ();
 FILLCELL_X1 PHY_3624 ();
 FILLCELL_X1 PHY_3625 ();
 FILLCELL_X1 PHY_3626 ();
 FILLCELL_X1 PHY_3627 ();
 FILLCELL_X1 PHY_3628 ();
 FILLCELL_X1 PHY_3629 ();
 FILLCELL_X1 PHY_363 ();
 FILLCELL_X1 PHY_3630 ();
 FILLCELL_X1 PHY_3631 ();
 FILLCELL_X1 PHY_3632 ();
 FILLCELL_X1 PHY_3633 ();
 FILLCELL_X1 PHY_3634 ();
 FILLCELL_X1 PHY_3635 ();
 FILLCELL_X1 PHY_3636 ();
 FILLCELL_X1 PHY_3637 ();
 FILLCELL_X1 PHY_3638 ();
 FILLCELL_X1 PHY_3639 ();
 FILLCELL_X1 PHY_364 ();
 FILLCELL_X1 PHY_3640 ();
 FILLCELL_X1 PHY_3641 ();
 FILLCELL_X1 PHY_3642 ();
 FILLCELL_X1 PHY_3643 ();
 FILLCELL_X1 PHY_3644 ();
 FILLCELL_X1 PHY_3645 ();
 FILLCELL_X1 PHY_3646 ();
 FILLCELL_X1 PHY_3647 ();
 FILLCELL_X1 PHY_3648 ();
 FILLCELL_X1 PHY_3649 ();
 FILLCELL_X1 PHY_365 ();
 FILLCELL_X1 PHY_3650 ();
 FILLCELL_X1 PHY_3651 ();
 FILLCELL_X1 PHY_3652 ();
 FILLCELL_X1 PHY_3653 ();
 FILLCELL_X1 PHY_3654 ();
 FILLCELL_X1 PHY_3655 ();
 FILLCELL_X1 PHY_3656 ();
 FILLCELL_X1 PHY_3657 ();
 FILLCELL_X1 PHY_3658 ();
 FILLCELL_X1 PHY_3659 ();
 FILLCELL_X1 PHY_366 ();
 FILLCELL_X1 PHY_3660 ();
 FILLCELL_X1 PHY_3661 ();
 FILLCELL_X1 PHY_3662 ();
 FILLCELL_X1 PHY_3663 ();
 FILLCELL_X1 PHY_3664 ();
 FILLCELL_X1 PHY_3665 ();
 FILLCELL_X1 PHY_3666 ();
 FILLCELL_X1 PHY_3667 ();
 FILLCELL_X1 PHY_3668 ();
 FILLCELL_X1 PHY_3669 ();
 FILLCELL_X1 PHY_367 ();
 FILLCELL_X1 PHY_3670 ();
 FILLCELL_X1 PHY_3671 ();
 FILLCELL_X1 PHY_3672 ();
 FILLCELL_X1 PHY_3673 ();
 FILLCELL_X1 PHY_3674 ();
 FILLCELL_X1 PHY_3675 ();
 FILLCELL_X1 PHY_3676 ();
 FILLCELL_X1 PHY_3677 ();
 FILLCELL_X1 PHY_3678 ();
 FILLCELL_X1 PHY_3679 ();
 FILLCELL_X1 PHY_368 ();
 FILLCELL_X1 PHY_3680 ();
 FILLCELL_X1 PHY_3681 ();
 FILLCELL_X1 PHY_3682 ();
 FILLCELL_X1 PHY_3683 ();
 FILLCELL_X1 PHY_3684 ();
 FILLCELL_X1 PHY_3685 ();
 FILLCELL_X1 PHY_3686 ();
 FILLCELL_X1 PHY_3687 ();
 FILLCELL_X1 PHY_3688 ();
 FILLCELL_X1 PHY_3689 ();
 FILLCELL_X1 PHY_369 ();
 FILLCELL_X1 PHY_3690 ();
 FILLCELL_X1 PHY_3691 ();
 FILLCELL_X1 PHY_3692 ();
 FILLCELL_X1 PHY_3693 ();
 FILLCELL_X1 PHY_3694 ();
 FILLCELL_X1 PHY_3695 ();
 FILLCELL_X1 PHY_3696 ();
 FILLCELL_X1 PHY_3697 ();
 FILLCELL_X1 PHY_3698 ();
 FILLCELL_X1 PHY_3699 ();
 FILLCELL_X1 PHY_37 ();
 FILLCELL_X1 PHY_370 ();
 FILLCELL_X1 PHY_3700 ();
 FILLCELL_X1 PHY_3701 ();
 FILLCELL_X1 PHY_3702 ();
 FILLCELL_X1 PHY_3703 ();
 FILLCELL_X1 PHY_3704 ();
 FILLCELL_X1 PHY_3705 ();
 FILLCELL_X1 PHY_3706 ();
 FILLCELL_X1 PHY_3707 ();
 FILLCELL_X1 PHY_3708 ();
 FILLCELL_X1 PHY_3709 ();
 FILLCELL_X1 PHY_371 ();
 FILLCELL_X1 PHY_3710 ();
 FILLCELL_X1 PHY_3711 ();
 FILLCELL_X1 PHY_3712 ();
 FILLCELL_X1 PHY_3713 ();
 FILLCELL_X1 PHY_3714 ();
 FILLCELL_X1 PHY_3715 ();
 FILLCELL_X1 PHY_3716 ();
 FILLCELL_X1 PHY_3717 ();
 FILLCELL_X1 PHY_3718 ();
 FILLCELL_X1 PHY_3719 ();
 FILLCELL_X1 PHY_372 ();
 FILLCELL_X1 PHY_3720 ();
 FILLCELL_X1 PHY_3721 ();
 FILLCELL_X1 PHY_3722 ();
 FILLCELL_X1 PHY_3723 ();
 FILLCELL_X1 PHY_3724 ();
 FILLCELL_X1 PHY_3725 ();
 FILLCELL_X1 PHY_3726 ();
 FILLCELL_X1 PHY_3727 ();
 FILLCELL_X1 PHY_3728 ();
 FILLCELL_X1 PHY_3729 ();
 FILLCELL_X1 PHY_373 ();
 FILLCELL_X1 PHY_3730 ();
 FILLCELL_X1 PHY_3731 ();
 FILLCELL_X1 PHY_3732 ();
 FILLCELL_X1 PHY_3733 ();
 FILLCELL_X1 PHY_3734 ();
 FILLCELL_X1 PHY_3735 ();
 FILLCELL_X1 PHY_3736 ();
 FILLCELL_X1 PHY_3737 ();
 FILLCELL_X1 PHY_3738 ();
 FILLCELL_X1 PHY_3739 ();
 FILLCELL_X1 PHY_374 ();
 FILLCELL_X1 PHY_3740 ();
 FILLCELL_X1 PHY_3741 ();
 FILLCELL_X1 PHY_3742 ();
 FILLCELL_X1 PHY_3743 ();
 FILLCELL_X1 PHY_3744 ();
 FILLCELL_X1 PHY_3745 ();
 FILLCELL_X1 PHY_3746 ();
 FILLCELL_X1 PHY_3747 ();
 FILLCELL_X1 PHY_3748 ();
 FILLCELL_X1 PHY_3749 ();
 FILLCELL_X1 PHY_375 ();
 FILLCELL_X1 PHY_3750 ();
 FILLCELL_X1 PHY_3751 ();
 FILLCELL_X1 PHY_3752 ();
 FILLCELL_X1 PHY_3753 ();
 FILLCELL_X1 PHY_3754 ();
 FILLCELL_X1 PHY_3755 ();
 FILLCELL_X1 PHY_3756 ();
 FILLCELL_X1 PHY_3757 ();
 FILLCELL_X1 PHY_3758 ();
 FILLCELL_X1 PHY_3759 ();
 FILLCELL_X1 PHY_376 ();
 FILLCELL_X1 PHY_3760 ();
 FILLCELL_X1 PHY_3761 ();
 FILLCELL_X1 PHY_3762 ();
 FILLCELL_X1 PHY_3763 ();
 FILLCELL_X1 PHY_3764 ();
 FILLCELL_X1 PHY_3765 ();
 FILLCELL_X1 PHY_3766 ();
 FILLCELL_X1 PHY_3767 ();
 FILLCELL_X1 PHY_3768 ();
 FILLCELL_X1 PHY_3769 ();
 FILLCELL_X1 PHY_377 ();
 FILLCELL_X1 PHY_3770 ();
 FILLCELL_X1 PHY_3771 ();
 FILLCELL_X1 PHY_3772 ();
 FILLCELL_X1 PHY_3773 ();
 FILLCELL_X1 PHY_3774 ();
 FILLCELL_X1 PHY_3775 ();
 FILLCELL_X1 PHY_3776 ();
 FILLCELL_X1 PHY_3777 ();
 FILLCELL_X1 PHY_3778 ();
 FILLCELL_X1 PHY_3779 ();
 FILLCELL_X1 PHY_378 ();
 FILLCELL_X1 PHY_3780 ();
 FILLCELL_X1 PHY_3781 ();
 FILLCELL_X1 PHY_3782 ();
 FILLCELL_X1 PHY_3783 ();
 FILLCELL_X1 PHY_3784 ();
 FILLCELL_X1 PHY_3785 ();
 FILLCELL_X1 PHY_3786 ();
 FILLCELL_X1 PHY_3787 ();
 FILLCELL_X1 PHY_3788 ();
 FILLCELL_X1 PHY_3789 ();
 FILLCELL_X1 PHY_379 ();
 FILLCELL_X1 PHY_3790 ();
 FILLCELL_X1 PHY_3791 ();
 FILLCELL_X1 PHY_3792 ();
 FILLCELL_X1 PHY_3793 ();
 FILLCELL_X1 PHY_3794 ();
 FILLCELL_X1 PHY_3795 ();
 FILLCELL_X1 PHY_3796 ();
 FILLCELL_X1 PHY_3797 ();
 FILLCELL_X1 PHY_3798 ();
 FILLCELL_X1 PHY_3799 ();
 FILLCELL_X1 PHY_38 ();
 FILLCELL_X1 PHY_380 ();
 FILLCELL_X1 PHY_3800 ();
 FILLCELL_X1 PHY_3801 ();
 FILLCELL_X1 PHY_3802 ();
 FILLCELL_X1 PHY_3803 ();
 FILLCELL_X1 PHY_3804 ();
 FILLCELL_X1 PHY_3805 ();
 FILLCELL_X1 PHY_3806 ();
 FILLCELL_X1 PHY_3807 ();
 FILLCELL_X1 PHY_3808 ();
 FILLCELL_X1 PHY_3809 ();
 FILLCELL_X1 PHY_381 ();
 FILLCELL_X1 PHY_3810 ();
 FILLCELL_X1 PHY_3811 ();
 FILLCELL_X1 PHY_3812 ();
 FILLCELL_X1 PHY_3813 ();
 FILLCELL_X1 PHY_3814 ();
 FILLCELL_X1 PHY_3815 ();
 FILLCELL_X1 PHY_3816 ();
 FILLCELL_X1 PHY_3817 ();
 FILLCELL_X1 PHY_3818 ();
 FILLCELL_X1 PHY_3819 ();
 FILLCELL_X1 PHY_382 ();
 FILLCELL_X1 PHY_3820 ();
 FILLCELL_X1 PHY_3821 ();
 FILLCELL_X1 PHY_3822 ();
 FILLCELL_X1 PHY_3823 ();
 FILLCELL_X1 PHY_3824 ();
 FILLCELL_X1 PHY_3825 ();
 FILLCELL_X1 PHY_3826 ();
 FILLCELL_X1 PHY_3827 ();
 FILLCELL_X1 PHY_3828 ();
 FILLCELL_X1 PHY_3829 ();
 FILLCELL_X1 PHY_383 ();
 FILLCELL_X1 PHY_3830 ();
 FILLCELL_X1 PHY_3831 ();
 FILLCELL_X1 PHY_3832 ();
 FILLCELL_X1 PHY_3833 ();
 FILLCELL_X1 PHY_3834 ();
 FILLCELL_X1 PHY_3835 ();
 FILLCELL_X1 PHY_3836 ();
 FILLCELL_X1 PHY_3837 ();
 FILLCELL_X1 PHY_3838 ();
 FILLCELL_X1 PHY_3839 ();
 FILLCELL_X1 PHY_384 ();
 FILLCELL_X1 PHY_3840 ();
 FILLCELL_X1 PHY_3841 ();
 FILLCELL_X1 PHY_3842 ();
 FILLCELL_X1 PHY_3843 ();
 FILLCELL_X1 PHY_3844 ();
 FILLCELL_X1 PHY_3845 ();
 FILLCELL_X1 PHY_3846 ();
 FILLCELL_X1 PHY_3847 ();
 FILLCELL_X1 PHY_3848 ();
 FILLCELL_X1 PHY_3849 ();
 FILLCELL_X1 PHY_385 ();
 FILLCELL_X1 PHY_3850 ();
 FILLCELL_X1 PHY_3851 ();
 FILLCELL_X1 PHY_3852 ();
 FILLCELL_X1 PHY_3853 ();
 FILLCELL_X1 PHY_3854 ();
 FILLCELL_X1 PHY_3855 ();
 FILLCELL_X1 PHY_3856 ();
 FILLCELL_X1 PHY_3857 ();
 FILLCELL_X1 PHY_3858 ();
 FILLCELL_X1 PHY_3859 ();
 FILLCELL_X1 PHY_386 ();
 FILLCELL_X1 PHY_3860 ();
 FILLCELL_X1 PHY_3861 ();
 FILLCELL_X1 PHY_3862 ();
 FILLCELL_X1 PHY_3863 ();
 FILLCELL_X1 PHY_3864 ();
 FILLCELL_X1 PHY_3865 ();
 FILLCELL_X1 PHY_3866 ();
 FILLCELL_X1 PHY_3867 ();
 FILLCELL_X1 PHY_3868 ();
 FILLCELL_X1 PHY_3869 ();
 FILLCELL_X1 PHY_387 ();
 FILLCELL_X1 PHY_3870 ();
 FILLCELL_X1 PHY_3871 ();
 FILLCELL_X1 PHY_3872 ();
 FILLCELL_X1 PHY_3873 ();
 FILLCELL_X1 PHY_3874 ();
 FILLCELL_X1 PHY_3875 ();
 FILLCELL_X1 PHY_3876 ();
 FILLCELL_X1 PHY_3877 ();
 FILLCELL_X1 PHY_3878 ();
 FILLCELL_X1 PHY_3879 ();
 FILLCELL_X1 PHY_388 ();
 FILLCELL_X1 PHY_3880 ();
 FILLCELL_X1 PHY_3881 ();
 FILLCELL_X1 PHY_3882 ();
 FILLCELL_X1 PHY_3883 ();
 FILLCELL_X1 PHY_3884 ();
 FILLCELL_X1 PHY_3885 ();
 FILLCELL_X1 PHY_3886 ();
 FILLCELL_X1 PHY_3887 ();
 FILLCELL_X1 PHY_3888 ();
 FILLCELL_X1 PHY_3889 ();
 FILLCELL_X1 PHY_389 ();
 FILLCELL_X1 PHY_3890 ();
 FILLCELL_X1 PHY_3891 ();
 FILLCELL_X1 PHY_3892 ();
 FILLCELL_X1 PHY_3893 ();
 FILLCELL_X1 PHY_3894 ();
 FILLCELL_X1 PHY_3895 ();
 FILLCELL_X1 PHY_3896 ();
 FILLCELL_X1 PHY_3897 ();
 FILLCELL_X1 PHY_3898 ();
 FILLCELL_X1 PHY_3899 ();
 FILLCELL_X1 PHY_39 ();
 FILLCELL_X1 PHY_390 ();
 FILLCELL_X1 PHY_3900 ();
 FILLCELL_X1 PHY_3901 ();
 FILLCELL_X1 PHY_3902 ();
 FILLCELL_X1 PHY_3903 ();
 FILLCELL_X1 PHY_3904 ();
 FILLCELL_X1 PHY_3905 ();
 FILLCELL_X1 PHY_3906 ();
 FILLCELL_X1 PHY_3907 ();
 FILLCELL_X1 PHY_3908 ();
 FILLCELL_X1 PHY_3909 ();
 FILLCELL_X1 PHY_391 ();
 FILLCELL_X1 PHY_3910 ();
 FILLCELL_X1 PHY_3911 ();
 FILLCELL_X1 PHY_3912 ();
 FILLCELL_X1 PHY_3913 ();
 FILLCELL_X1 PHY_3914 ();
 FILLCELL_X1 PHY_3915 ();
 FILLCELL_X1 PHY_3916 ();
 FILLCELL_X1 PHY_3917 ();
 FILLCELL_X1 PHY_3918 ();
 FILLCELL_X1 PHY_3919 ();
 FILLCELL_X1 PHY_392 ();
 FILLCELL_X1 PHY_3920 ();
 FILLCELL_X1 PHY_3921 ();
 FILLCELL_X1 PHY_3922 ();
 FILLCELL_X1 PHY_3923 ();
 FILLCELL_X1 PHY_3924 ();
 FILLCELL_X1 PHY_3925 ();
 FILLCELL_X1 PHY_3926 ();
 FILLCELL_X1 PHY_3927 ();
 FILLCELL_X1 PHY_3928 ();
 FILLCELL_X1 PHY_3929 ();
 FILLCELL_X1 PHY_393 ();
 FILLCELL_X1 PHY_3930 ();
 FILLCELL_X1 PHY_3931 ();
 FILLCELL_X1 PHY_3932 ();
 FILLCELL_X1 PHY_3933 ();
 FILLCELL_X1 PHY_3934 ();
 FILLCELL_X1 PHY_3935 ();
 FILLCELL_X1 PHY_3936 ();
 FILLCELL_X1 PHY_3937 ();
 FILLCELL_X1 PHY_3938 ();
 FILLCELL_X1 PHY_3939 ();
 FILLCELL_X1 PHY_394 ();
 FILLCELL_X1 PHY_3940 ();
 FILLCELL_X1 PHY_3941 ();
 FILLCELL_X1 PHY_3942 ();
 FILLCELL_X1 PHY_3943 ();
 FILLCELL_X1 PHY_3944 ();
 FILLCELL_X1 PHY_3945 ();
 FILLCELL_X1 PHY_3946 ();
 FILLCELL_X1 PHY_3947 ();
 FILLCELL_X1 PHY_3948 ();
 FILLCELL_X1 PHY_3949 ();
 FILLCELL_X1 PHY_395 ();
 FILLCELL_X1 PHY_3950 ();
 FILLCELL_X1 PHY_3951 ();
 FILLCELL_X1 PHY_3952 ();
 FILLCELL_X1 PHY_3953 ();
 FILLCELL_X1 PHY_3954 ();
 FILLCELL_X1 PHY_3955 ();
 FILLCELL_X1 PHY_3956 ();
 FILLCELL_X1 PHY_3957 ();
 FILLCELL_X1 PHY_3958 ();
 FILLCELL_X1 PHY_3959 ();
 FILLCELL_X1 PHY_396 ();
 FILLCELL_X1 PHY_3960 ();
 FILLCELL_X1 PHY_3961 ();
 FILLCELL_X1 PHY_3962 ();
 FILLCELL_X1 PHY_3963 ();
 FILLCELL_X1 PHY_3964 ();
 FILLCELL_X1 PHY_3965 ();
 FILLCELL_X1 PHY_3966 ();
 FILLCELL_X1 PHY_3967 ();
 FILLCELL_X1 PHY_3968 ();
 FILLCELL_X1 PHY_3969 ();
 FILLCELL_X1 PHY_397 ();
 FILLCELL_X1 PHY_3970 ();
 FILLCELL_X1 PHY_3971 ();
 FILLCELL_X1 PHY_3972 ();
 FILLCELL_X1 PHY_3973 ();
 FILLCELL_X1 PHY_3974 ();
 FILLCELL_X1 PHY_3975 ();
 FILLCELL_X1 PHY_3976 ();
 FILLCELL_X1 PHY_3977 ();
 FILLCELL_X1 PHY_3978 ();
 FILLCELL_X1 PHY_3979 ();
 FILLCELL_X1 PHY_398 ();
 FILLCELL_X1 PHY_3980 ();
 FILLCELL_X1 PHY_3981 ();
 FILLCELL_X1 PHY_3982 ();
 FILLCELL_X1 PHY_3983 ();
 FILLCELL_X1 PHY_3984 ();
 FILLCELL_X1 PHY_3985 ();
 FILLCELL_X1 PHY_3986 ();
 FILLCELL_X1 PHY_3987 ();
 FILLCELL_X1 PHY_3988 ();
 FILLCELL_X1 PHY_3989 ();
 FILLCELL_X1 PHY_399 ();
 FILLCELL_X1 PHY_3990 ();
 FILLCELL_X1 PHY_3991 ();
 FILLCELL_X1 PHY_3992 ();
 FILLCELL_X1 PHY_3993 ();
 FILLCELL_X1 PHY_3994 ();
 FILLCELL_X1 PHY_3995 ();
 FILLCELL_X1 PHY_3996 ();
 FILLCELL_X1 PHY_3997 ();
 FILLCELL_X1 PHY_3998 ();
 FILLCELL_X1 PHY_3999 ();
 FILLCELL_X1 PHY_4 ();
 FILLCELL_X1 PHY_40 ();
 FILLCELL_X1 PHY_400 ();
 FILLCELL_X1 PHY_4000 ();
 FILLCELL_X1 PHY_4001 ();
 FILLCELL_X1 PHY_4002 ();
 FILLCELL_X1 PHY_4003 ();
 FILLCELL_X1 PHY_4004 ();
 FILLCELL_X1 PHY_4005 ();
 FILLCELL_X1 PHY_4006 ();
 FILLCELL_X1 PHY_4007 ();
 FILLCELL_X1 PHY_4008 ();
 FILLCELL_X1 PHY_4009 ();
 FILLCELL_X1 PHY_401 ();
 FILLCELL_X1 PHY_4010 ();
 FILLCELL_X1 PHY_4011 ();
 FILLCELL_X1 PHY_4012 ();
 FILLCELL_X1 PHY_4013 ();
 FILLCELL_X1 PHY_4014 ();
 FILLCELL_X1 PHY_4015 ();
 FILLCELL_X1 PHY_4016 ();
 FILLCELL_X1 PHY_4017 ();
 FILLCELL_X1 PHY_4018 ();
 FILLCELL_X1 PHY_4019 ();
 FILLCELL_X1 PHY_402 ();
 FILLCELL_X1 PHY_4020 ();
 FILLCELL_X1 PHY_4021 ();
 FILLCELL_X1 PHY_4022 ();
 FILLCELL_X1 PHY_4023 ();
 FILLCELL_X1 PHY_4024 ();
 FILLCELL_X1 PHY_4025 ();
 FILLCELL_X1 PHY_4026 ();
 FILLCELL_X1 PHY_4027 ();
 FILLCELL_X1 PHY_4028 ();
 FILLCELL_X1 PHY_4029 ();
 FILLCELL_X1 PHY_403 ();
 FILLCELL_X1 PHY_4030 ();
 FILLCELL_X1 PHY_4031 ();
 FILLCELL_X1 PHY_4032 ();
 FILLCELL_X1 PHY_4033 ();
 FILLCELL_X1 PHY_4034 ();
 FILLCELL_X1 PHY_4035 ();
 FILLCELL_X1 PHY_4036 ();
 FILLCELL_X1 PHY_4037 ();
 FILLCELL_X1 PHY_4038 ();
 FILLCELL_X1 PHY_4039 ();
 FILLCELL_X1 PHY_404 ();
 FILLCELL_X1 PHY_4040 ();
 FILLCELL_X1 PHY_4041 ();
 FILLCELL_X1 PHY_4042 ();
 FILLCELL_X1 PHY_4043 ();
 FILLCELL_X1 PHY_4044 ();
 FILLCELL_X1 PHY_4045 ();
 FILLCELL_X1 PHY_4046 ();
 FILLCELL_X1 PHY_4047 ();
 FILLCELL_X1 PHY_4048 ();
 FILLCELL_X1 PHY_4049 ();
 FILLCELL_X1 PHY_405 ();
 FILLCELL_X1 PHY_4050 ();
 FILLCELL_X1 PHY_4051 ();
 FILLCELL_X1 PHY_4052 ();
 FILLCELL_X1 PHY_4053 ();
 FILLCELL_X1 PHY_4054 ();
 FILLCELL_X1 PHY_4055 ();
 FILLCELL_X1 PHY_4056 ();
 FILLCELL_X1 PHY_4057 ();
 FILLCELL_X1 PHY_4058 ();
 FILLCELL_X1 PHY_4059 ();
 FILLCELL_X1 PHY_406 ();
 FILLCELL_X1 PHY_4060 ();
 FILLCELL_X1 PHY_4061 ();
 FILLCELL_X1 PHY_4062 ();
 FILLCELL_X1 PHY_4063 ();
 FILLCELL_X1 PHY_4064 ();
 FILLCELL_X1 PHY_4065 ();
 FILLCELL_X1 PHY_4066 ();
 FILLCELL_X1 PHY_4067 ();
 FILLCELL_X1 PHY_4068 ();
 FILLCELL_X1 PHY_4069 ();
 FILLCELL_X1 PHY_407 ();
 FILLCELL_X1 PHY_4070 ();
 FILLCELL_X1 PHY_4071 ();
 FILLCELL_X1 PHY_4072 ();
 FILLCELL_X1 PHY_4073 ();
 FILLCELL_X1 PHY_4074 ();
 FILLCELL_X1 PHY_4075 ();
 FILLCELL_X1 PHY_4076 ();
 FILLCELL_X1 PHY_4077 ();
 FILLCELL_X1 PHY_4078 ();
 FILLCELL_X1 PHY_4079 ();
 FILLCELL_X1 PHY_408 ();
 FILLCELL_X1 PHY_4080 ();
 FILLCELL_X1 PHY_4081 ();
 FILLCELL_X1 PHY_4082 ();
 FILLCELL_X1 PHY_4083 ();
 FILLCELL_X1 PHY_4084 ();
 FILLCELL_X1 PHY_4085 ();
 FILLCELL_X1 PHY_4086 ();
 FILLCELL_X1 PHY_4087 ();
 FILLCELL_X1 PHY_4088 ();
 FILLCELL_X1 PHY_4089 ();
 FILLCELL_X1 PHY_409 ();
 FILLCELL_X1 PHY_4090 ();
 FILLCELL_X1 PHY_4091 ();
 FILLCELL_X1 PHY_4092 ();
 FILLCELL_X1 PHY_4093 ();
 FILLCELL_X1 PHY_4094 ();
 FILLCELL_X1 PHY_4095 ();
 FILLCELL_X1 PHY_4096 ();
 FILLCELL_X1 PHY_4097 ();
 FILLCELL_X1 PHY_4098 ();
 FILLCELL_X1 PHY_4099 ();
 FILLCELL_X1 PHY_41 ();
 FILLCELL_X1 PHY_410 ();
 FILLCELL_X1 PHY_4100 ();
 FILLCELL_X1 PHY_4101 ();
 FILLCELL_X1 PHY_4102 ();
 FILLCELL_X1 PHY_4103 ();
 FILLCELL_X1 PHY_4104 ();
 FILLCELL_X1 PHY_4105 ();
 FILLCELL_X1 PHY_4106 ();
 FILLCELL_X1 PHY_4107 ();
 FILLCELL_X1 PHY_4108 ();
 FILLCELL_X1 PHY_4109 ();
 FILLCELL_X1 PHY_411 ();
 FILLCELL_X1 PHY_4110 ();
 FILLCELL_X1 PHY_4111 ();
 FILLCELL_X1 PHY_4112 ();
 FILLCELL_X1 PHY_4113 ();
 FILLCELL_X1 PHY_4114 ();
 FILLCELL_X1 PHY_4115 ();
 FILLCELL_X1 PHY_4116 ();
 FILLCELL_X1 PHY_4117 ();
 FILLCELL_X1 PHY_4118 ();
 FILLCELL_X1 PHY_4119 ();
 FILLCELL_X1 PHY_412 ();
 FILLCELL_X1 PHY_4120 ();
 FILLCELL_X1 PHY_4121 ();
 FILLCELL_X1 PHY_4122 ();
 FILLCELL_X1 PHY_4123 ();
 FILLCELL_X1 PHY_4124 ();
 FILLCELL_X1 PHY_4125 ();
 FILLCELL_X1 PHY_4126 ();
 FILLCELL_X1 PHY_4127 ();
 FILLCELL_X1 PHY_4128 ();
 FILLCELL_X1 PHY_4129 ();
 FILLCELL_X1 PHY_413 ();
 FILLCELL_X1 PHY_4130 ();
 FILLCELL_X1 PHY_4131 ();
 FILLCELL_X1 PHY_4132 ();
 FILLCELL_X1 PHY_4133 ();
 FILLCELL_X1 PHY_4134 ();
 FILLCELL_X1 PHY_4135 ();
 FILLCELL_X1 PHY_4136 ();
 FILLCELL_X1 PHY_4137 ();
 FILLCELL_X1 PHY_4138 ();
 FILLCELL_X1 PHY_4139 ();
 FILLCELL_X1 PHY_414 ();
 FILLCELL_X1 PHY_4140 ();
 FILLCELL_X1 PHY_4141 ();
 FILLCELL_X1 PHY_4142 ();
 FILLCELL_X1 PHY_4143 ();
 FILLCELL_X1 PHY_4144 ();
 FILLCELL_X1 PHY_4145 ();
 FILLCELL_X1 PHY_4146 ();
 FILLCELL_X1 PHY_4147 ();
 FILLCELL_X1 PHY_4148 ();
 FILLCELL_X1 PHY_4149 ();
 FILLCELL_X1 PHY_415 ();
 FILLCELL_X1 PHY_4150 ();
 FILLCELL_X1 PHY_4151 ();
 FILLCELL_X1 PHY_4152 ();
 FILLCELL_X1 PHY_4153 ();
 FILLCELL_X1 PHY_4154 ();
 FILLCELL_X1 PHY_4155 ();
 FILLCELL_X1 PHY_4156 ();
 FILLCELL_X1 PHY_4157 ();
 FILLCELL_X1 PHY_4158 ();
 FILLCELL_X1 PHY_4159 ();
 FILLCELL_X1 PHY_416 ();
 FILLCELL_X1 PHY_4160 ();
 FILLCELL_X1 PHY_4161 ();
 FILLCELL_X1 PHY_4162 ();
 FILLCELL_X1 PHY_4163 ();
 FILLCELL_X1 PHY_4164 ();
 FILLCELL_X1 PHY_4165 ();
 FILLCELL_X1 PHY_4166 ();
 FILLCELL_X1 PHY_4167 ();
 FILLCELL_X1 PHY_4168 ();
 FILLCELL_X1 PHY_4169 ();
 FILLCELL_X1 PHY_417 ();
 FILLCELL_X1 PHY_4170 ();
 FILLCELL_X1 PHY_4171 ();
 FILLCELL_X1 PHY_4172 ();
 FILLCELL_X1 PHY_4173 ();
 FILLCELL_X1 PHY_4174 ();
 FILLCELL_X1 PHY_4175 ();
 FILLCELL_X1 PHY_4176 ();
 FILLCELL_X1 PHY_4177 ();
 FILLCELL_X1 PHY_4178 ();
 FILLCELL_X1 PHY_4179 ();
 FILLCELL_X1 PHY_418 ();
 FILLCELL_X1 PHY_4180 ();
 FILLCELL_X1 PHY_4181 ();
 FILLCELL_X1 PHY_4182 ();
 FILLCELL_X1 PHY_4183 ();
 FILLCELL_X1 PHY_4184 ();
 FILLCELL_X1 PHY_4185 ();
 FILLCELL_X1 PHY_4186 ();
 FILLCELL_X1 PHY_4187 ();
 FILLCELL_X1 PHY_4188 ();
 FILLCELL_X1 PHY_4189 ();
 FILLCELL_X1 PHY_419 ();
 FILLCELL_X1 PHY_4190 ();
 FILLCELL_X1 PHY_4191 ();
 FILLCELL_X1 PHY_4192 ();
 FILLCELL_X1 PHY_4193 ();
 FILLCELL_X1 PHY_4194 ();
 FILLCELL_X1 PHY_4195 ();
 FILLCELL_X1 PHY_4196 ();
 FILLCELL_X1 PHY_4197 ();
 FILLCELL_X1 PHY_4198 ();
 FILLCELL_X1 PHY_4199 ();
 FILLCELL_X1 PHY_42 ();
 FILLCELL_X1 PHY_420 ();
 FILLCELL_X1 PHY_4200 ();
 FILLCELL_X1 PHY_4201 ();
 FILLCELL_X1 PHY_4202 ();
 FILLCELL_X1 PHY_4203 ();
 FILLCELL_X1 PHY_4204 ();
 FILLCELL_X1 PHY_4205 ();
 FILLCELL_X1 PHY_4206 ();
 FILLCELL_X1 PHY_4207 ();
 FILLCELL_X1 PHY_4208 ();
 FILLCELL_X1 PHY_4209 ();
 FILLCELL_X1 PHY_421 ();
 FILLCELL_X1 PHY_4210 ();
 FILLCELL_X1 PHY_4211 ();
 FILLCELL_X1 PHY_4212 ();
 FILLCELL_X1 PHY_4213 ();
 FILLCELL_X1 PHY_4214 ();
 FILLCELL_X1 PHY_4215 ();
 FILLCELL_X1 PHY_4216 ();
 FILLCELL_X1 PHY_4217 ();
 FILLCELL_X1 PHY_4218 ();
 FILLCELL_X1 PHY_4219 ();
 FILLCELL_X1 PHY_422 ();
 FILLCELL_X1 PHY_4220 ();
 FILLCELL_X1 PHY_4221 ();
 FILLCELL_X1 PHY_4222 ();
 FILLCELL_X1 PHY_4223 ();
 FILLCELL_X1 PHY_4224 ();
 FILLCELL_X1 PHY_4225 ();
 FILLCELL_X1 PHY_4226 ();
 FILLCELL_X1 PHY_4227 ();
 FILLCELL_X1 PHY_4228 ();
 FILLCELL_X1 PHY_4229 ();
 FILLCELL_X1 PHY_423 ();
 FILLCELL_X1 PHY_4230 ();
 FILLCELL_X1 PHY_4231 ();
 FILLCELL_X1 PHY_4232 ();
 FILLCELL_X1 PHY_4233 ();
 FILLCELL_X1 PHY_4234 ();
 FILLCELL_X1 PHY_4235 ();
 FILLCELL_X1 PHY_4236 ();
 FILLCELL_X1 PHY_4237 ();
 FILLCELL_X1 PHY_4238 ();
 FILLCELL_X1 PHY_4239 ();
 FILLCELL_X1 PHY_424 ();
 FILLCELL_X1 PHY_4240 ();
 FILLCELL_X1 PHY_4241 ();
 FILLCELL_X1 PHY_4242 ();
 FILLCELL_X1 PHY_4243 ();
 FILLCELL_X1 PHY_4244 ();
 FILLCELL_X1 PHY_4245 ();
 FILLCELL_X1 PHY_4246 ();
 FILLCELL_X1 PHY_4247 ();
 FILLCELL_X1 PHY_4248 ();
 FILLCELL_X1 PHY_4249 ();
 FILLCELL_X1 PHY_425 ();
 FILLCELL_X1 PHY_4250 ();
 FILLCELL_X1 PHY_4251 ();
 FILLCELL_X1 PHY_4252 ();
 FILLCELL_X1 PHY_4253 ();
 FILLCELL_X1 PHY_4254 ();
 FILLCELL_X1 PHY_4255 ();
 FILLCELL_X1 PHY_4256 ();
 FILLCELL_X1 PHY_4257 ();
 FILLCELL_X1 PHY_4258 ();
 FILLCELL_X1 PHY_4259 ();
 FILLCELL_X1 PHY_426 ();
 FILLCELL_X1 PHY_4260 ();
 FILLCELL_X1 PHY_4261 ();
 FILLCELL_X1 PHY_4262 ();
 FILLCELL_X1 PHY_4263 ();
 FILLCELL_X1 PHY_4264 ();
 FILLCELL_X1 PHY_4265 ();
 FILLCELL_X1 PHY_4266 ();
 FILLCELL_X1 PHY_4267 ();
 FILLCELL_X1 PHY_4268 ();
 FILLCELL_X1 PHY_4269 ();
 FILLCELL_X1 PHY_427 ();
 FILLCELL_X1 PHY_4270 ();
 FILLCELL_X1 PHY_4271 ();
 FILLCELL_X1 PHY_4272 ();
 FILLCELL_X1 PHY_4273 ();
 FILLCELL_X1 PHY_4274 ();
 FILLCELL_X1 PHY_4275 ();
 FILLCELL_X1 PHY_4276 ();
 FILLCELL_X1 PHY_4277 ();
 FILLCELL_X1 PHY_4278 ();
 FILLCELL_X1 PHY_4279 ();
 FILLCELL_X1 PHY_428 ();
 FILLCELL_X1 PHY_4280 ();
 FILLCELL_X1 PHY_4281 ();
 FILLCELL_X1 PHY_4282 ();
 FILLCELL_X1 PHY_4283 ();
 FILLCELL_X1 PHY_4284 ();
 FILLCELL_X1 PHY_4285 ();
 FILLCELL_X1 PHY_4286 ();
 FILLCELL_X1 PHY_4287 ();
 FILLCELL_X1 PHY_4288 ();
 FILLCELL_X1 PHY_4289 ();
 FILLCELL_X1 PHY_429 ();
 FILLCELL_X1 PHY_4290 ();
 FILLCELL_X1 PHY_4291 ();
 FILLCELL_X1 PHY_4292 ();
 FILLCELL_X1 PHY_4293 ();
 FILLCELL_X1 PHY_4294 ();
 FILLCELL_X1 PHY_4295 ();
 FILLCELL_X1 PHY_4296 ();
 FILLCELL_X1 PHY_4297 ();
 FILLCELL_X1 PHY_4298 ();
 FILLCELL_X1 PHY_4299 ();
 FILLCELL_X1 PHY_43 ();
 FILLCELL_X1 PHY_430 ();
 FILLCELL_X1 PHY_4300 ();
 FILLCELL_X1 PHY_4301 ();
 FILLCELL_X1 PHY_4302 ();
 FILLCELL_X1 PHY_4303 ();
 FILLCELL_X1 PHY_4304 ();
 FILLCELL_X1 PHY_4305 ();
 FILLCELL_X1 PHY_4306 ();
 FILLCELL_X1 PHY_4307 ();
 FILLCELL_X1 PHY_4308 ();
 FILLCELL_X1 PHY_4309 ();
 FILLCELL_X1 PHY_431 ();
 FILLCELL_X1 PHY_4310 ();
 FILLCELL_X1 PHY_4311 ();
 FILLCELL_X1 PHY_4312 ();
 FILLCELL_X1 PHY_4313 ();
 FILLCELL_X1 PHY_4314 ();
 FILLCELL_X1 PHY_4315 ();
 FILLCELL_X1 PHY_4316 ();
 FILLCELL_X1 PHY_4317 ();
 FILLCELL_X1 PHY_4318 ();
 FILLCELL_X1 PHY_4319 ();
 FILLCELL_X1 PHY_432 ();
 FILLCELL_X1 PHY_4320 ();
 FILLCELL_X1 PHY_4321 ();
 FILLCELL_X1 PHY_4322 ();
 FILLCELL_X1 PHY_4323 ();
 FILLCELL_X1 PHY_4324 ();
 FILLCELL_X1 PHY_4325 ();
 FILLCELL_X1 PHY_4326 ();
 FILLCELL_X1 PHY_4327 ();
 FILLCELL_X1 PHY_4328 ();
 FILLCELL_X1 PHY_4329 ();
 FILLCELL_X1 PHY_433 ();
 FILLCELL_X1 PHY_4330 ();
 FILLCELL_X1 PHY_4331 ();
 FILLCELL_X1 PHY_4332 ();
 FILLCELL_X1 PHY_4333 ();
 FILLCELL_X1 PHY_4334 ();
 FILLCELL_X1 PHY_4335 ();
 FILLCELL_X1 PHY_4336 ();
 FILLCELL_X1 PHY_4337 ();
 FILLCELL_X1 PHY_4338 ();
 FILLCELL_X1 PHY_4339 ();
 FILLCELL_X1 PHY_434 ();
 FILLCELL_X1 PHY_4340 ();
 FILLCELL_X1 PHY_4341 ();
 FILLCELL_X1 PHY_4342 ();
 FILLCELL_X1 PHY_4343 ();
 FILLCELL_X1 PHY_4344 ();
 FILLCELL_X1 PHY_4345 ();
 FILLCELL_X1 PHY_4346 ();
 FILLCELL_X1 PHY_4347 ();
 FILLCELL_X1 PHY_4348 ();
 FILLCELL_X1 PHY_4349 ();
 FILLCELL_X1 PHY_435 ();
 FILLCELL_X1 PHY_4350 ();
 FILLCELL_X1 PHY_4351 ();
 FILLCELL_X1 PHY_4352 ();
 FILLCELL_X1 PHY_4353 ();
 FILLCELL_X1 PHY_4354 ();
 FILLCELL_X1 PHY_4355 ();
 FILLCELL_X1 PHY_4356 ();
 FILLCELL_X1 PHY_4357 ();
 FILLCELL_X1 PHY_4358 ();
 FILLCELL_X1 PHY_4359 ();
 FILLCELL_X1 PHY_436 ();
 FILLCELL_X1 PHY_4360 ();
 FILLCELL_X1 PHY_4361 ();
 FILLCELL_X1 PHY_4362 ();
 FILLCELL_X1 PHY_4363 ();
 FILLCELL_X1 PHY_4364 ();
 FILLCELL_X1 PHY_4365 ();
 FILLCELL_X1 PHY_4366 ();
 FILLCELL_X1 PHY_4367 ();
 FILLCELL_X1 PHY_4368 ();
 FILLCELL_X1 PHY_4369 ();
 FILLCELL_X1 PHY_437 ();
 FILLCELL_X1 PHY_4370 ();
 FILLCELL_X1 PHY_4371 ();
 FILLCELL_X1 PHY_4372 ();
 FILLCELL_X1 PHY_4373 ();
 FILLCELL_X1 PHY_4374 ();
 FILLCELL_X1 PHY_4375 ();
 FILLCELL_X1 PHY_4376 ();
 FILLCELL_X1 PHY_4377 ();
 FILLCELL_X1 PHY_4378 ();
 FILLCELL_X1 PHY_4379 ();
 FILLCELL_X1 PHY_438 ();
 FILLCELL_X1 PHY_4380 ();
 FILLCELL_X1 PHY_4381 ();
 FILLCELL_X1 PHY_4382 ();
 FILLCELL_X1 PHY_4383 ();
 FILLCELL_X1 PHY_4384 ();
 FILLCELL_X1 PHY_4385 ();
 FILLCELL_X1 PHY_4386 ();
 FILLCELL_X1 PHY_4387 ();
 FILLCELL_X1 PHY_4388 ();
 FILLCELL_X1 PHY_4389 ();
 FILLCELL_X1 PHY_439 ();
 FILLCELL_X1 PHY_4390 ();
 FILLCELL_X1 PHY_4391 ();
 FILLCELL_X1 PHY_4392 ();
 FILLCELL_X1 PHY_4393 ();
 FILLCELL_X1 PHY_4394 ();
 FILLCELL_X1 PHY_4395 ();
 FILLCELL_X1 PHY_4396 ();
 FILLCELL_X1 PHY_4397 ();
 FILLCELL_X1 PHY_4398 ();
 FILLCELL_X1 PHY_4399 ();
 FILLCELL_X1 PHY_44 ();
 FILLCELL_X1 PHY_440 ();
 FILLCELL_X1 PHY_4400 ();
 FILLCELL_X1 PHY_4401 ();
 FILLCELL_X1 PHY_4402 ();
 FILLCELL_X1 PHY_4403 ();
 FILLCELL_X1 PHY_4404 ();
 FILLCELL_X1 PHY_4405 ();
 FILLCELL_X1 PHY_4406 ();
 FILLCELL_X1 PHY_4407 ();
 FILLCELL_X1 PHY_4408 ();
 FILLCELL_X1 PHY_4409 ();
 FILLCELL_X1 PHY_441 ();
 FILLCELL_X1 PHY_4410 ();
 FILLCELL_X1 PHY_4411 ();
 FILLCELL_X1 PHY_4412 ();
 FILLCELL_X1 PHY_4413 ();
 FILLCELL_X1 PHY_4414 ();
 FILLCELL_X1 PHY_4415 ();
 FILLCELL_X1 PHY_4416 ();
 FILLCELL_X1 PHY_4417 ();
 FILLCELL_X1 PHY_4418 ();
 FILLCELL_X1 PHY_4419 ();
 FILLCELL_X1 PHY_442 ();
 FILLCELL_X1 PHY_4420 ();
 FILLCELL_X1 PHY_4421 ();
 FILLCELL_X1 PHY_4422 ();
 FILLCELL_X1 PHY_4423 ();
 FILLCELL_X1 PHY_4424 ();
 FILLCELL_X1 PHY_4425 ();
 FILLCELL_X1 PHY_4426 ();
 FILLCELL_X1 PHY_4427 ();
 FILLCELL_X1 PHY_4428 ();
 FILLCELL_X1 PHY_4429 ();
 FILLCELL_X1 PHY_443 ();
 FILLCELL_X1 PHY_4430 ();
 FILLCELL_X1 PHY_4431 ();
 FILLCELL_X1 PHY_4432 ();
 FILLCELL_X1 PHY_4433 ();
 FILLCELL_X1 PHY_4434 ();
 FILLCELL_X1 PHY_4435 ();
 FILLCELL_X1 PHY_4436 ();
 FILLCELL_X1 PHY_4437 ();
 FILLCELL_X1 PHY_4438 ();
 FILLCELL_X1 PHY_4439 ();
 FILLCELL_X1 PHY_444 ();
 FILLCELL_X1 PHY_4440 ();
 FILLCELL_X1 PHY_4441 ();
 FILLCELL_X1 PHY_4442 ();
 FILLCELL_X1 PHY_4443 ();
 FILLCELL_X1 PHY_4444 ();
 FILLCELL_X1 PHY_4445 ();
 FILLCELL_X1 PHY_4446 ();
 FILLCELL_X1 PHY_4447 ();
 FILLCELL_X1 PHY_4448 ();
 FILLCELL_X1 PHY_4449 ();
 FILLCELL_X1 PHY_445 ();
 FILLCELL_X1 PHY_4450 ();
 FILLCELL_X1 PHY_4451 ();
 FILLCELL_X1 PHY_4452 ();
 FILLCELL_X1 PHY_4453 ();
 FILLCELL_X1 PHY_4454 ();
 FILLCELL_X1 PHY_4455 ();
 FILLCELL_X1 PHY_4456 ();
 FILLCELL_X1 PHY_4457 ();
 FILLCELL_X1 PHY_4458 ();
 FILLCELL_X1 PHY_4459 ();
 FILLCELL_X1 PHY_446 ();
 FILLCELL_X1 PHY_4460 ();
 FILLCELL_X1 PHY_4461 ();
 FILLCELL_X1 PHY_4462 ();
 FILLCELL_X1 PHY_4463 ();
 FILLCELL_X1 PHY_4464 ();
 FILLCELL_X1 PHY_4465 ();
 FILLCELL_X1 PHY_4466 ();
 FILLCELL_X1 PHY_4467 ();
 FILLCELL_X1 PHY_4468 ();
 FILLCELL_X1 PHY_4469 ();
 FILLCELL_X1 PHY_447 ();
 FILLCELL_X1 PHY_4470 ();
 FILLCELL_X1 PHY_4471 ();
 FILLCELL_X1 PHY_4472 ();
 FILLCELL_X1 PHY_4473 ();
 FILLCELL_X1 PHY_4474 ();
 FILLCELL_X1 PHY_4475 ();
 FILLCELL_X1 PHY_4476 ();
 FILLCELL_X1 PHY_4477 ();
 FILLCELL_X1 PHY_4478 ();
 FILLCELL_X1 PHY_4479 ();
 FILLCELL_X1 PHY_448 ();
 FILLCELL_X1 PHY_4480 ();
 FILLCELL_X1 PHY_4481 ();
 FILLCELL_X1 PHY_4482 ();
 FILLCELL_X1 PHY_4483 ();
 FILLCELL_X1 PHY_4484 ();
 FILLCELL_X1 PHY_4485 ();
 FILLCELL_X1 PHY_4486 ();
 FILLCELL_X1 PHY_4487 ();
 FILLCELL_X1 PHY_4488 ();
 FILLCELL_X1 PHY_4489 ();
 FILLCELL_X1 PHY_449 ();
 FILLCELL_X1 PHY_4490 ();
 FILLCELL_X1 PHY_4491 ();
 FILLCELL_X1 PHY_4492 ();
 FILLCELL_X1 PHY_4493 ();
 FILLCELL_X1 PHY_4494 ();
 FILLCELL_X1 PHY_4495 ();
 FILLCELL_X1 PHY_4496 ();
 FILLCELL_X1 PHY_4497 ();
 FILLCELL_X1 PHY_4498 ();
 FILLCELL_X1 PHY_4499 ();
 FILLCELL_X1 PHY_45 ();
 FILLCELL_X1 PHY_450 ();
 FILLCELL_X1 PHY_4500 ();
 FILLCELL_X1 PHY_4501 ();
 FILLCELL_X1 PHY_4502 ();
 FILLCELL_X1 PHY_4503 ();
 FILLCELL_X1 PHY_4504 ();
 FILLCELL_X1 PHY_4505 ();
 FILLCELL_X1 PHY_4506 ();
 FILLCELL_X1 PHY_4507 ();
 FILLCELL_X1 PHY_4508 ();
 FILLCELL_X1 PHY_4509 ();
 FILLCELL_X1 PHY_451 ();
 FILLCELL_X1 PHY_4510 ();
 FILLCELL_X1 PHY_4511 ();
 FILLCELL_X1 PHY_4512 ();
 FILLCELL_X1 PHY_4513 ();
 FILLCELL_X1 PHY_4514 ();
 FILLCELL_X1 PHY_4515 ();
 FILLCELL_X1 PHY_4516 ();
 FILLCELL_X1 PHY_4517 ();
 FILLCELL_X1 PHY_4518 ();
 FILLCELL_X1 PHY_4519 ();
 FILLCELL_X1 PHY_452 ();
 FILLCELL_X1 PHY_4520 ();
 FILLCELL_X1 PHY_4521 ();
 FILLCELL_X1 PHY_4522 ();
 FILLCELL_X1 PHY_4523 ();
 FILLCELL_X1 PHY_4524 ();
 FILLCELL_X1 PHY_4525 ();
 FILLCELL_X1 PHY_4526 ();
 FILLCELL_X1 PHY_4527 ();
 FILLCELL_X1 PHY_4528 ();
 FILLCELL_X1 PHY_4529 ();
 FILLCELL_X1 PHY_453 ();
 FILLCELL_X1 PHY_4530 ();
 FILLCELL_X1 PHY_4531 ();
 FILLCELL_X1 PHY_4532 ();
 FILLCELL_X1 PHY_4533 ();
 FILLCELL_X1 PHY_4534 ();
 FILLCELL_X1 PHY_4535 ();
 FILLCELL_X1 PHY_4536 ();
 FILLCELL_X1 PHY_4537 ();
 FILLCELL_X1 PHY_4538 ();
 FILLCELL_X1 PHY_4539 ();
 FILLCELL_X1 PHY_454 ();
 FILLCELL_X1 PHY_4540 ();
 FILLCELL_X1 PHY_4541 ();
 FILLCELL_X1 PHY_4542 ();
 FILLCELL_X1 PHY_4543 ();
 FILLCELL_X1 PHY_4544 ();
 FILLCELL_X1 PHY_4545 ();
 FILLCELL_X1 PHY_4546 ();
 FILLCELL_X1 PHY_4547 ();
 FILLCELL_X1 PHY_4548 ();
 FILLCELL_X1 PHY_4549 ();
 FILLCELL_X1 PHY_455 ();
 FILLCELL_X1 PHY_4550 ();
 FILLCELL_X1 PHY_4551 ();
 FILLCELL_X1 PHY_4552 ();
 FILLCELL_X1 PHY_4553 ();
 FILLCELL_X1 PHY_4554 ();
 FILLCELL_X1 PHY_4555 ();
 FILLCELL_X1 PHY_4556 ();
 FILLCELL_X1 PHY_4557 ();
 FILLCELL_X1 PHY_4558 ();
 FILLCELL_X1 PHY_4559 ();
 FILLCELL_X1 PHY_456 ();
 FILLCELL_X1 PHY_4560 ();
 FILLCELL_X1 PHY_4561 ();
 FILLCELL_X1 PHY_4562 ();
 FILLCELL_X1 PHY_4563 ();
 FILLCELL_X1 PHY_4564 ();
 FILLCELL_X1 PHY_4565 ();
 FILLCELL_X1 PHY_4566 ();
 FILLCELL_X1 PHY_4567 ();
 FILLCELL_X1 PHY_4568 ();
 FILLCELL_X1 PHY_4569 ();
 FILLCELL_X1 PHY_457 ();
 FILLCELL_X1 PHY_4570 ();
 FILLCELL_X1 PHY_4571 ();
 FILLCELL_X1 PHY_4572 ();
 FILLCELL_X1 PHY_4573 ();
 FILLCELL_X1 PHY_4574 ();
 FILLCELL_X1 PHY_4575 ();
 FILLCELL_X1 PHY_4576 ();
 FILLCELL_X1 PHY_4577 ();
 FILLCELL_X1 PHY_4578 ();
 FILLCELL_X1 PHY_4579 ();
 FILLCELL_X1 PHY_458 ();
 FILLCELL_X1 PHY_4580 ();
 FILLCELL_X1 PHY_4581 ();
 FILLCELL_X1 PHY_4582 ();
 FILLCELL_X1 PHY_4583 ();
 FILLCELL_X1 PHY_4584 ();
 FILLCELL_X1 PHY_4585 ();
 FILLCELL_X1 PHY_4586 ();
 FILLCELL_X1 PHY_4587 ();
 FILLCELL_X1 PHY_4588 ();
 FILLCELL_X1 PHY_4589 ();
 FILLCELL_X1 PHY_459 ();
 FILLCELL_X1 PHY_4590 ();
 FILLCELL_X1 PHY_4591 ();
 FILLCELL_X1 PHY_4592 ();
 FILLCELL_X1 PHY_4593 ();
 FILLCELL_X1 PHY_4594 ();
 FILLCELL_X1 PHY_4595 ();
 FILLCELL_X1 PHY_4596 ();
 FILLCELL_X1 PHY_4597 ();
 FILLCELL_X1 PHY_4598 ();
 FILLCELL_X1 PHY_4599 ();
 FILLCELL_X1 PHY_46 ();
 FILLCELL_X1 PHY_460 ();
 FILLCELL_X1 PHY_4600 ();
 FILLCELL_X1 PHY_4601 ();
 FILLCELL_X1 PHY_4602 ();
 FILLCELL_X1 PHY_4603 ();
 FILLCELL_X1 PHY_4604 ();
 FILLCELL_X1 PHY_4605 ();
 FILLCELL_X1 PHY_4606 ();
 FILLCELL_X1 PHY_4607 ();
 FILLCELL_X1 PHY_4608 ();
 FILLCELL_X1 PHY_4609 ();
 FILLCELL_X1 PHY_461 ();
 FILLCELL_X1 PHY_4610 ();
 FILLCELL_X1 PHY_4611 ();
 FILLCELL_X1 PHY_4612 ();
 FILLCELL_X1 PHY_4613 ();
 FILLCELL_X1 PHY_4614 ();
 FILLCELL_X1 PHY_4615 ();
 FILLCELL_X1 PHY_4616 ();
 FILLCELL_X1 PHY_4617 ();
 FILLCELL_X1 PHY_4618 ();
 FILLCELL_X1 PHY_4619 ();
 FILLCELL_X1 PHY_462 ();
 FILLCELL_X1 PHY_4620 ();
 FILLCELL_X1 PHY_4621 ();
 FILLCELL_X1 PHY_4622 ();
 FILLCELL_X1 PHY_4623 ();
 FILLCELL_X1 PHY_4624 ();
 FILLCELL_X1 PHY_4625 ();
 FILLCELL_X1 PHY_4626 ();
 FILLCELL_X1 PHY_4627 ();
 FILLCELL_X1 PHY_4628 ();
 FILLCELL_X1 PHY_4629 ();
 FILLCELL_X1 PHY_463 ();
 FILLCELL_X1 PHY_4630 ();
 FILLCELL_X1 PHY_4631 ();
 FILLCELL_X1 PHY_4632 ();
 FILLCELL_X1 PHY_4633 ();
 FILLCELL_X1 PHY_4634 ();
 FILLCELL_X1 PHY_4635 ();
 FILLCELL_X1 PHY_4636 ();
 FILLCELL_X1 PHY_4637 ();
 FILLCELL_X1 PHY_4638 ();
 FILLCELL_X1 PHY_4639 ();
 FILLCELL_X1 PHY_464 ();
 FILLCELL_X1 PHY_4640 ();
 FILLCELL_X1 PHY_4641 ();
 FILLCELL_X1 PHY_4642 ();
 FILLCELL_X1 PHY_4643 ();
 FILLCELL_X1 PHY_4644 ();
 FILLCELL_X1 PHY_4645 ();
 FILLCELL_X1 PHY_4646 ();
 FILLCELL_X1 PHY_4647 ();
 FILLCELL_X1 PHY_4648 ();
 FILLCELL_X1 PHY_4649 ();
 FILLCELL_X1 PHY_465 ();
 FILLCELL_X1 PHY_4650 ();
 FILLCELL_X1 PHY_4651 ();
 FILLCELL_X1 PHY_4652 ();
 FILLCELL_X1 PHY_4653 ();
 FILLCELL_X1 PHY_4654 ();
 FILLCELL_X1 PHY_4655 ();
 FILLCELL_X1 PHY_4656 ();
 FILLCELL_X1 PHY_4657 ();
 FILLCELL_X1 PHY_4658 ();
 FILLCELL_X1 PHY_4659 ();
 FILLCELL_X1 PHY_466 ();
 FILLCELL_X1 PHY_4660 ();
 FILLCELL_X1 PHY_4661 ();
 FILLCELL_X1 PHY_4662 ();
 FILLCELL_X1 PHY_4663 ();
 FILLCELL_X1 PHY_4664 ();
 FILLCELL_X1 PHY_4665 ();
 FILLCELL_X1 PHY_4666 ();
 FILLCELL_X1 PHY_4667 ();
 FILLCELL_X1 PHY_4668 ();
 FILLCELL_X1 PHY_4669 ();
 FILLCELL_X1 PHY_467 ();
 FILLCELL_X1 PHY_4670 ();
 FILLCELL_X1 PHY_4671 ();
 FILLCELL_X1 PHY_4672 ();
 FILLCELL_X1 PHY_4673 ();
 FILLCELL_X1 PHY_4674 ();
 FILLCELL_X1 PHY_4675 ();
 FILLCELL_X1 PHY_4676 ();
 FILLCELL_X1 PHY_4677 ();
 FILLCELL_X1 PHY_4678 ();
 FILLCELL_X1 PHY_4679 ();
 FILLCELL_X1 PHY_468 ();
 FILLCELL_X1 PHY_4680 ();
 FILLCELL_X1 PHY_4681 ();
 FILLCELL_X1 PHY_4682 ();
 FILLCELL_X1 PHY_4683 ();
 FILLCELL_X1 PHY_4684 ();
 FILLCELL_X1 PHY_4685 ();
 FILLCELL_X1 PHY_4686 ();
 FILLCELL_X1 PHY_4687 ();
 FILLCELL_X1 PHY_4688 ();
 FILLCELL_X1 PHY_4689 ();
 FILLCELL_X1 PHY_469 ();
 FILLCELL_X1 PHY_4690 ();
 FILLCELL_X1 PHY_4691 ();
 FILLCELL_X1 PHY_4692 ();
 FILLCELL_X1 PHY_4693 ();
 FILLCELL_X1 PHY_4694 ();
 FILLCELL_X1 PHY_4695 ();
 FILLCELL_X1 PHY_4696 ();
 FILLCELL_X1 PHY_4697 ();
 FILLCELL_X1 PHY_4698 ();
 FILLCELL_X1 PHY_4699 ();
 FILLCELL_X1 PHY_47 ();
 FILLCELL_X1 PHY_470 ();
 FILLCELL_X1 PHY_4700 ();
 FILLCELL_X1 PHY_4701 ();
 FILLCELL_X1 PHY_4702 ();
 FILLCELL_X1 PHY_4703 ();
 FILLCELL_X1 PHY_4704 ();
 FILLCELL_X1 PHY_4705 ();
 FILLCELL_X1 PHY_4706 ();
 FILLCELL_X1 PHY_4707 ();
 FILLCELL_X1 PHY_4708 ();
 FILLCELL_X1 PHY_4709 ();
 FILLCELL_X1 PHY_471 ();
 FILLCELL_X1 PHY_4710 ();
 FILLCELL_X1 PHY_4711 ();
 FILLCELL_X1 PHY_4712 ();
 FILLCELL_X1 PHY_4713 ();
 FILLCELL_X1 PHY_4714 ();
 FILLCELL_X1 PHY_4715 ();
 FILLCELL_X1 PHY_4716 ();
 FILLCELL_X1 PHY_4717 ();
 FILLCELL_X1 PHY_4718 ();
 FILLCELL_X1 PHY_4719 ();
 FILLCELL_X1 PHY_472 ();
 FILLCELL_X1 PHY_4720 ();
 FILLCELL_X1 PHY_4721 ();
 FILLCELL_X1 PHY_4722 ();
 FILLCELL_X1 PHY_4723 ();
 FILLCELL_X1 PHY_4724 ();
 FILLCELL_X1 PHY_4725 ();
 FILLCELL_X1 PHY_4726 ();
 FILLCELL_X1 PHY_4727 ();
 FILLCELL_X1 PHY_4728 ();
 FILLCELL_X1 PHY_4729 ();
 FILLCELL_X1 PHY_473 ();
 FILLCELL_X1 PHY_4730 ();
 FILLCELL_X1 PHY_4731 ();
 FILLCELL_X1 PHY_4732 ();
 FILLCELL_X1 PHY_4733 ();
 FILLCELL_X1 PHY_4734 ();
 FILLCELL_X1 PHY_4735 ();
 FILLCELL_X1 PHY_4736 ();
 FILLCELL_X1 PHY_4737 ();
 FILLCELL_X1 PHY_4738 ();
 FILLCELL_X1 PHY_4739 ();
 FILLCELL_X1 PHY_474 ();
 FILLCELL_X1 PHY_4740 ();
 FILLCELL_X1 PHY_4741 ();
 FILLCELL_X1 PHY_4742 ();
 FILLCELL_X1 PHY_4743 ();
 FILLCELL_X1 PHY_4744 ();
 FILLCELL_X1 PHY_4745 ();
 FILLCELL_X1 PHY_4746 ();
 FILLCELL_X1 PHY_4747 ();
 FILLCELL_X1 PHY_4748 ();
 FILLCELL_X1 PHY_4749 ();
 FILLCELL_X1 PHY_475 ();
 FILLCELL_X1 PHY_4750 ();
 FILLCELL_X1 PHY_4751 ();
 FILLCELL_X1 PHY_4752 ();
 FILLCELL_X1 PHY_4753 ();
 FILLCELL_X1 PHY_4754 ();
 FILLCELL_X1 PHY_4755 ();
 FILLCELL_X1 PHY_4756 ();
 FILLCELL_X1 PHY_4757 ();
 FILLCELL_X1 PHY_4758 ();
 FILLCELL_X1 PHY_4759 ();
 FILLCELL_X1 PHY_476 ();
 FILLCELL_X1 PHY_4760 ();
 FILLCELL_X1 PHY_4761 ();
 FILLCELL_X1 PHY_4762 ();
 FILLCELL_X1 PHY_4763 ();
 FILLCELL_X1 PHY_4764 ();
 FILLCELL_X1 PHY_4765 ();
 FILLCELL_X1 PHY_4766 ();
 FILLCELL_X1 PHY_4767 ();
 FILLCELL_X1 PHY_4768 ();
 FILLCELL_X1 PHY_4769 ();
 FILLCELL_X1 PHY_477 ();
 FILLCELL_X1 PHY_4770 ();
 FILLCELL_X1 PHY_4771 ();
 FILLCELL_X1 PHY_4772 ();
 FILLCELL_X1 PHY_4773 ();
 FILLCELL_X1 PHY_4774 ();
 FILLCELL_X1 PHY_4775 ();
 FILLCELL_X1 PHY_4776 ();
 FILLCELL_X1 PHY_4777 ();
 FILLCELL_X1 PHY_4778 ();
 FILLCELL_X1 PHY_4779 ();
 FILLCELL_X1 PHY_478 ();
 FILLCELL_X1 PHY_4780 ();
 FILLCELL_X1 PHY_4781 ();
 FILLCELL_X1 PHY_4782 ();
 FILLCELL_X1 PHY_4783 ();
 FILLCELL_X1 PHY_4784 ();
 FILLCELL_X1 PHY_4785 ();
 FILLCELL_X1 PHY_4786 ();
 FILLCELL_X1 PHY_4787 ();
 FILLCELL_X1 PHY_4788 ();
 FILLCELL_X1 PHY_4789 ();
 FILLCELL_X1 PHY_479 ();
 FILLCELL_X1 PHY_4790 ();
 FILLCELL_X1 PHY_4791 ();
 FILLCELL_X1 PHY_4792 ();
 FILLCELL_X1 PHY_4793 ();
 FILLCELL_X1 PHY_4794 ();
 FILLCELL_X1 PHY_4795 ();
 FILLCELL_X1 PHY_4796 ();
 FILLCELL_X1 PHY_4797 ();
 FILLCELL_X1 PHY_4798 ();
 FILLCELL_X1 PHY_4799 ();
 FILLCELL_X1 PHY_48 ();
 FILLCELL_X1 PHY_480 ();
 FILLCELL_X1 PHY_4800 ();
 FILLCELL_X1 PHY_4801 ();
 FILLCELL_X1 PHY_4802 ();
 FILLCELL_X1 PHY_4803 ();
 FILLCELL_X1 PHY_4804 ();
 FILLCELL_X1 PHY_4805 ();
 FILLCELL_X1 PHY_4806 ();
 FILLCELL_X1 PHY_4807 ();
 FILLCELL_X1 PHY_4808 ();
 FILLCELL_X1 PHY_4809 ();
 FILLCELL_X1 PHY_481 ();
 FILLCELL_X1 PHY_4810 ();
 FILLCELL_X1 PHY_4811 ();
 FILLCELL_X1 PHY_4812 ();
 FILLCELL_X1 PHY_4813 ();
 FILLCELL_X1 PHY_4814 ();
 FILLCELL_X1 PHY_4815 ();
 FILLCELL_X1 PHY_4816 ();
 FILLCELL_X1 PHY_4817 ();
 FILLCELL_X1 PHY_4818 ();
 FILLCELL_X1 PHY_4819 ();
 FILLCELL_X1 PHY_482 ();
 FILLCELL_X1 PHY_4820 ();
 FILLCELL_X1 PHY_4821 ();
 FILLCELL_X1 PHY_4822 ();
 FILLCELL_X1 PHY_4823 ();
 FILLCELL_X1 PHY_4824 ();
 FILLCELL_X1 PHY_4825 ();
 FILLCELL_X1 PHY_4826 ();
 FILLCELL_X1 PHY_4827 ();
 FILLCELL_X1 PHY_4828 ();
 FILLCELL_X1 PHY_4829 ();
 FILLCELL_X1 PHY_483 ();
 FILLCELL_X1 PHY_4830 ();
 FILLCELL_X1 PHY_4831 ();
 FILLCELL_X1 PHY_4832 ();
 FILLCELL_X1 PHY_4833 ();
 FILLCELL_X1 PHY_4834 ();
 FILLCELL_X1 PHY_4835 ();
 FILLCELL_X1 PHY_4836 ();
 FILLCELL_X1 PHY_4837 ();
 FILLCELL_X1 PHY_4838 ();
 FILLCELL_X1 PHY_4839 ();
 FILLCELL_X1 PHY_484 ();
 FILLCELL_X1 PHY_4840 ();
 FILLCELL_X1 PHY_4841 ();
 FILLCELL_X1 PHY_4842 ();
 FILLCELL_X1 PHY_4843 ();
 FILLCELL_X1 PHY_4844 ();
 FILLCELL_X1 PHY_4845 ();
 FILLCELL_X1 PHY_4846 ();
 FILLCELL_X1 PHY_4847 ();
 FILLCELL_X1 PHY_4848 ();
 FILLCELL_X1 PHY_4849 ();
 FILLCELL_X1 PHY_485 ();
 FILLCELL_X1 PHY_4850 ();
 FILLCELL_X1 PHY_4851 ();
 FILLCELL_X1 PHY_4852 ();
 FILLCELL_X1 PHY_4853 ();
 FILLCELL_X1 PHY_4854 ();
 FILLCELL_X1 PHY_4855 ();
 FILLCELL_X1 PHY_4856 ();
 FILLCELL_X1 PHY_4857 ();
 FILLCELL_X1 PHY_4858 ();
 FILLCELL_X1 PHY_4859 ();
 FILLCELL_X1 PHY_486 ();
 FILLCELL_X1 PHY_4860 ();
 FILLCELL_X1 PHY_4861 ();
 FILLCELL_X1 PHY_4862 ();
 FILLCELL_X1 PHY_4863 ();
 FILLCELL_X1 PHY_4864 ();
 FILLCELL_X1 PHY_4865 ();
 FILLCELL_X1 PHY_4866 ();
 FILLCELL_X1 PHY_4867 ();
 FILLCELL_X1 PHY_4868 ();
 FILLCELL_X1 PHY_4869 ();
 FILLCELL_X1 PHY_487 ();
 FILLCELL_X1 PHY_4870 ();
 FILLCELL_X1 PHY_4871 ();
 FILLCELL_X1 PHY_4872 ();
 FILLCELL_X1 PHY_4873 ();
 FILLCELL_X1 PHY_4874 ();
 FILLCELL_X1 PHY_4875 ();
 FILLCELL_X1 PHY_4876 ();
 FILLCELL_X1 PHY_4877 ();
 FILLCELL_X1 PHY_4878 ();
 FILLCELL_X1 PHY_4879 ();
 FILLCELL_X1 PHY_488 ();
 FILLCELL_X1 PHY_4880 ();
 FILLCELL_X1 PHY_4881 ();
 FILLCELL_X1 PHY_4882 ();
 FILLCELL_X1 PHY_4883 ();
 FILLCELL_X1 PHY_4884 ();
 FILLCELL_X1 PHY_4885 ();
 FILLCELL_X1 PHY_4886 ();
 FILLCELL_X1 PHY_4887 ();
 FILLCELL_X1 PHY_4888 ();
 FILLCELL_X1 PHY_4889 ();
 FILLCELL_X1 PHY_489 ();
 FILLCELL_X1 PHY_4890 ();
 FILLCELL_X1 PHY_4891 ();
 FILLCELL_X1 PHY_4892 ();
 FILLCELL_X1 PHY_4893 ();
 FILLCELL_X1 PHY_4894 ();
 FILLCELL_X1 PHY_4895 ();
 FILLCELL_X1 PHY_4896 ();
 FILLCELL_X1 PHY_4897 ();
 FILLCELL_X1 PHY_4898 ();
 FILLCELL_X1 PHY_4899 ();
 FILLCELL_X1 PHY_49 ();
 FILLCELL_X1 PHY_490 ();
 FILLCELL_X1 PHY_4900 ();
 FILLCELL_X1 PHY_4901 ();
 FILLCELL_X1 PHY_4902 ();
 FILLCELL_X1 PHY_4903 ();
 FILLCELL_X1 PHY_4904 ();
 FILLCELL_X1 PHY_4905 ();
 FILLCELL_X1 PHY_4906 ();
 FILLCELL_X1 PHY_4907 ();
 FILLCELL_X1 PHY_4908 ();
 FILLCELL_X1 PHY_4909 ();
 FILLCELL_X1 PHY_491 ();
 FILLCELL_X1 PHY_4910 ();
 FILLCELL_X1 PHY_4911 ();
 FILLCELL_X1 PHY_4912 ();
 FILLCELL_X1 PHY_4913 ();
 FILLCELL_X1 PHY_4914 ();
 FILLCELL_X1 PHY_4915 ();
 FILLCELL_X1 PHY_4916 ();
 FILLCELL_X1 PHY_4917 ();
 FILLCELL_X1 PHY_4918 ();
 FILLCELL_X1 PHY_4919 ();
 FILLCELL_X1 PHY_492 ();
 FILLCELL_X1 PHY_4920 ();
 FILLCELL_X1 PHY_4921 ();
 FILLCELL_X1 PHY_4922 ();
 FILLCELL_X1 PHY_4923 ();
 FILLCELL_X1 PHY_4924 ();
 FILLCELL_X1 PHY_4925 ();
 FILLCELL_X1 PHY_4926 ();
 FILLCELL_X1 PHY_4927 ();
 FILLCELL_X1 PHY_4928 ();
 FILLCELL_X1 PHY_4929 ();
 FILLCELL_X1 PHY_493 ();
 FILLCELL_X1 PHY_4930 ();
 FILLCELL_X1 PHY_4931 ();
 FILLCELL_X1 PHY_4932 ();
 FILLCELL_X1 PHY_4933 ();
 FILLCELL_X1 PHY_4934 ();
 FILLCELL_X1 PHY_4935 ();
 FILLCELL_X1 PHY_4936 ();
 FILLCELL_X1 PHY_4937 ();
 FILLCELL_X1 PHY_4938 ();
 FILLCELL_X1 PHY_4939 ();
 FILLCELL_X1 PHY_494 ();
 FILLCELL_X1 PHY_4940 ();
 FILLCELL_X1 PHY_4941 ();
 FILLCELL_X1 PHY_4942 ();
 FILLCELL_X1 PHY_4943 ();
 FILLCELL_X1 PHY_4944 ();
 FILLCELL_X1 PHY_4945 ();
 FILLCELL_X1 PHY_4946 ();
 FILLCELL_X1 PHY_4947 ();
 FILLCELL_X1 PHY_4948 ();
 FILLCELL_X1 PHY_4949 ();
 FILLCELL_X1 PHY_495 ();
 FILLCELL_X1 PHY_4950 ();
 FILLCELL_X1 PHY_4951 ();
 FILLCELL_X1 PHY_4952 ();
 FILLCELL_X1 PHY_4953 ();
 FILLCELL_X1 PHY_4954 ();
 FILLCELL_X1 PHY_4955 ();
 FILLCELL_X1 PHY_4956 ();
 FILLCELL_X1 PHY_4957 ();
 FILLCELL_X1 PHY_4958 ();
 FILLCELL_X1 PHY_4959 ();
 FILLCELL_X1 PHY_496 ();
 FILLCELL_X1 PHY_4960 ();
 FILLCELL_X1 PHY_4961 ();
 FILLCELL_X1 PHY_4962 ();
 FILLCELL_X1 PHY_4963 ();
 FILLCELL_X1 PHY_4964 ();
 FILLCELL_X1 PHY_4965 ();
 FILLCELL_X1 PHY_4966 ();
 FILLCELL_X1 PHY_4967 ();
 FILLCELL_X1 PHY_4968 ();
 FILLCELL_X1 PHY_4969 ();
 FILLCELL_X1 PHY_497 ();
 FILLCELL_X1 PHY_4970 ();
 FILLCELL_X1 PHY_4971 ();
 FILLCELL_X1 PHY_4972 ();
 FILLCELL_X1 PHY_4973 ();
 FILLCELL_X1 PHY_4974 ();
 FILLCELL_X1 PHY_4975 ();
 FILLCELL_X1 PHY_4976 ();
 FILLCELL_X1 PHY_4977 ();
 FILLCELL_X1 PHY_4978 ();
 FILLCELL_X1 PHY_4979 ();
 FILLCELL_X1 PHY_498 ();
 FILLCELL_X1 PHY_4980 ();
 FILLCELL_X1 PHY_4981 ();
 FILLCELL_X1 PHY_4982 ();
 FILLCELL_X1 PHY_4983 ();
 FILLCELL_X1 PHY_4984 ();
 FILLCELL_X1 PHY_4985 ();
 FILLCELL_X1 PHY_4986 ();
 FILLCELL_X1 PHY_4987 ();
 FILLCELL_X1 PHY_4988 ();
 FILLCELL_X1 PHY_4989 ();
 FILLCELL_X1 PHY_499 ();
 FILLCELL_X1 PHY_4990 ();
 FILLCELL_X1 PHY_4991 ();
 FILLCELL_X1 PHY_4992 ();
 FILLCELL_X1 PHY_4993 ();
 FILLCELL_X1 PHY_4994 ();
 FILLCELL_X1 PHY_4995 ();
 FILLCELL_X1 PHY_4996 ();
 FILLCELL_X1 PHY_4997 ();
 FILLCELL_X1 PHY_4998 ();
 FILLCELL_X1 PHY_4999 ();
 FILLCELL_X1 PHY_5 ();
 FILLCELL_X1 PHY_50 ();
 FILLCELL_X1 PHY_500 ();
 FILLCELL_X1 PHY_5000 ();
 FILLCELL_X1 PHY_5001 ();
 FILLCELL_X1 PHY_5002 ();
 FILLCELL_X1 PHY_5003 ();
 FILLCELL_X1 PHY_5004 ();
 FILLCELL_X1 PHY_5005 ();
 FILLCELL_X1 PHY_5006 ();
 FILLCELL_X1 PHY_5007 ();
 FILLCELL_X1 PHY_5008 ();
 FILLCELL_X1 PHY_5009 ();
 FILLCELL_X1 PHY_501 ();
 FILLCELL_X1 PHY_5010 ();
 FILLCELL_X1 PHY_5011 ();
 FILLCELL_X1 PHY_5012 ();
 FILLCELL_X1 PHY_5013 ();
 FILLCELL_X1 PHY_5014 ();
 FILLCELL_X1 PHY_5015 ();
 FILLCELL_X1 PHY_5016 ();
 FILLCELL_X1 PHY_5017 ();
 FILLCELL_X1 PHY_5018 ();
 FILLCELL_X1 PHY_5019 ();
 FILLCELL_X1 PHY_502 ();
 FILLCELL_X1 PHY_5020 ();
 FILLCELL_X1 PHY_5021 ();
 FILLCELL_X1 PHY_5022 ();
 FILLCELL_X1 PHY_5023 ();
 FILLCELL_X1 PHY_5024 ();
 FILLCELL_X1 PHY_5025 ();
 FILLCELL_X1 PHY_5026 ();
 FILLCELL_X1 PHY_5027 ();
 FILLCELL_X1 PHY_5028 ();
 FILLCELL_X1 PHY_5029 ();
 FILLCELL_X1 PHY_503 ();
 FILLCELL_X1 PHY_5030 ();
 FILLCELL_X1 PHY_5031 ();
 FILLCELL_X1 PHY_5032 ();
 FILLCELL_X1 PHY_5033 ();
 FILLCELL_X1 PHY_5034 ();
 FILLCELL_X1 PHY_5035 ();
 FILLCELL_X1 PHY_5036 ();
 FILLCELL_X1 PHY_5037 ();
 FILLCELL_X1 PHY_5038 ();
 FILLCELL_X1 PHY_5039 ();
 FILLCELL_X1 PHY_504 ();
 FILLCELL_X1 PHY_5040 ();
 FILLCELL_X1 PHY_5041 ();
 FILLCELL_X1 PHY_5042 ();
 FILLCELL_X1 PHY_5043 ();
 FILLCELL_X1 PHY_5044 ();
 FILLCELL_X1 PHY_5045 ();
 FILLCELL_X1 PHY_5046 ();
 FILLCELL_X1 PHY_5047 ();
 FILLCELL_X1 PHY_5048 ();
 FILLCELL_X1 PHY_5049 ();
 FILLCELL_X1 PHY_505 ();
 FILLCELL_X1 PHY_5050 ();
 FILLCELL_X1 PHY_5051 ();
 FILLCELL_X1 PHY_5052 ();
 FILLCELL_X1 PHY_5053 ();
 FILLCELL_X1 PHY_5054 ();
 FILLCELL_X1 PHY_5055 ();
 FILLCELL_X1 PHY_5056 ();
 FILLCELL_X1 PHY_5057 ();
 FILLCELL_X1 PHY_5058 ();
 FILLCELL_X1 PHY_5059 ();
 FILLCELL_X1 PHY_506 ();
 FILLCELL_X1 PHY_5060 ();
 FILLCELL_X1 PHY_5061 ();
 FILLCELL_X1 PHY_5062 ();
 FILLCELL_X1 PHY_5063 ();
 FILLCELL_X1 PHY_5064 ();
 FILLCELL_X1 PHY_5065 ();
 FILLCELL_X1 PHY_5066 ();
 FILLCELL_X1 PHY_5067 ();
 FILLCELL_X1 PHY_5068 ();
 FILLCELL_X1 PHY_5069 ();
 FILLCELL_X1 PHY_507 ();
 FILLCELL_X1 PHY_5070 ();
 FILLCELL_X1 PHY_5071 ();
 FILLCELL_X1 PHY_5072 ();
 FILLCELL_X1 PHY_5073 ();
 FILLCELL_X1 PHY_5074 ();
 FILLCELL_X1 PHY_5075 ();
 FILLCELL_X1 PHY_5076 ();
 FILLCELL_X1 PHY_5077 ();
 FILLCELL_X1 PHY_5078 ();
 FILLCELL_X1 PHY_5079 ();
 FILLCELL_X1 PHY_508 ();
 FILLCELL_X1 PHY_5080 ();
 FILLCELL_X1 PHY_5081 ();
 FILLCELL_X1 PHY_5082 ();
 FILLCELL_X1 PHY_5083 ();
 FILLCELL_X1 PHY_5084 ();
 FILLCELL_X1 PHY_5085 ();
 FILLCELL_X1 PHY_5086 ();
 FILLCELL_X1 PHY_5087 ();
 FILLCELL_X1 PHY_5088 ();
 FILLCELL_X1 PHY_5089 ();
 FILLCELL_X1 PHY_509 ();
 FILLCELL_X1 PHY_5090 ();
 FILLCELL_X1 PHY_5091 ();
 FILLCELL_X1 PHY_5092 ();
 FILLCELL_X1 PHY_5093 ();
 FILLCELL_X1 PHY_5094 ();
 FILLCELL_X1 PHY_5095 ();
 FILLCELL_X1 PHY_5096 ();
 FILLCELL_X1 PHY_5097 ();
 FILLCELL_X1 PHY_5098 ();
 FILLCELL_X1 PHY_5099 ();
 FILLCELL_X1 PHY_51 ();
 FILLCELL_X1 PHY_510 ();
 FILLCELL_X1 PHY_5100 ();
 FILLCELL_X1 PHY_5101 ();
 FILLCELL_X1 PHY_5102 ();
 FILLCELL_X1 PHY_5103 ();
 FILLCELL_X1 PHY_5104 ();
 FILLCELL_X1 PHY_5105 ();
 FILLCELL_X1 PHY_5106 ();
 FILLCELL_X1 PHY_5107 ();
 FILLCELL_X1 PHY_5108 ();
 FILLCELL_X1 PHY_5109 ();
 FILLCELL_X1 PHY_511 ();
 FILLCELL_X1 PHY_5110 ();
 FILLCELL_X1 PHY_5111 ();
 FILLCELL_X1 PHY_5112 ();
 FILLCELL_X1 PHY_5113 ();
 FILLCELL_X1 PHY_5114 ();
 FILLCELL_X1 PHY_5115 ();
 FILLCELL_X1 PHY_5116 ();
 FILLCELL_X1 PHY_5117 ();
 FILLCELL_X1 PHY_5118 ();
 FILLCELL_X1 PHY_5119 ();
 FILLCELL_X1 PHY_512 ();
 FILLCELL_X1 PHY_5120 ();
 FILLCELL_X1 PHY_5121 ();
 FILLCELL_X1 PHY_5122 ();
 FILLCELL_X1 PHY_5123 ();
 FILLCELL_X1 PHY_5124 ();
 FILLCELL_X1 PHY_5125 ();
 FILLCELL_X1 PHY_5126 ();
 FILLCELL_X1 PHY_5127 ();
 FILLCELL_X1 PHY_5128 ();
 FILLCELL_X1 PHY_5129 ();
 FILLCELL_X1 PHY_513 ();
 FILLCELL_X1 PHY_5130 ();
 FILLCELL_X1 PHY_5131 ();
 FILLCELL_X1 PHY_5132 ();
 FILLCELL_X1 PHY_5133 ();
 FILLCELL_X1 PHY_5134 ();
 FILLCELL_X1 PHY_5135 ();
 FILLCELL_X1 PHY_5136 ();
 FILLCELL_X1 PHY_5137 ();
 FILLCELL_X1 PHY_5138 ();
 FILLCELL_X1 PHY_5139 ();
 FILLCELL_X1 PHY_514 ();
 FILLCELL_X1 PHY_5140 ();
 FILLCELL_X1 PHY_5141 ();
 FILLCELL_X1 PHY_5142 ();
 FILLCELL_X1 PHY_5143 ();
 FILLCELL_X1 PHY_5144 ();
 FILLCELL_X1 PHY_5145 ();
 FILLCELL_X1 PHY_5146 ();
 FILLCELL_X1 PHY_5147 ();
 FILLCELL_X1 PHY_5148 ();
 FILLCELL_X1 PHY_5149 ();
 FILLCELL_X1 PHY_515 ();
 FILLCELL_X1 PHY_5150 ();
 FILLCELL_X1 PHY_5151 ();
 FILLCELL_X1 PHY_5152 ();
 FILLCELL_X1 PHY_5153 ();
 FILLCELL_X1 PHY_5154 ();
 FILLCELL_X1 PHY_5155 ();
 FILLCELL_X1 PHY_5156 ();
 FILLCELL_X1 PHY_5157 ();
 FILLCELL_X1 PHY_5158 ();
 FILLCELL_X1 PHY_5159 ();
 FILLCELL_X1 PHY_516 ();
 FILLCELL_X1 PHY_5160 ();
 FILLCELL_X1 PHY_5161 ();
 FILLCELL_X1 PHY_5162 ();
 FILLCELL_X1 PHY_5163 ();
 FILLCELL_X1 PHY_5164 ();
 FILLCELL_X1 PHY_5165 ();
 FILLCELL_X1 PHY_5166 ();
 FILLCELL_X1 PHY_5167 ();
 FILLCELL_X1 PHY_5168 ();
 FILLCELL_X1 PHY_5169 ();
 FILLCELL_X1 PHY_517 ();
 FILLCELL_X1 PHY_5170 ();
 FILLCELL_X1 PHY_5171 ();
 FILLCELL_X1 PHY_5172 ();
 FILLCELL_X1 PHY_5173 ();
 FILLCELL_X1 PHY_5174 ();
 FILLCELL_X1 PHY_5175 ();
 FILLCELL_X1 PHY_5176 ();
 FILLCELL_X1 PHY_5177 ();
 FILLCELL_X1 PHY_5178 ();
 FILLCELL_X1 PHY_5179 ();
 FILLCELL_X1 PHY_518 ();
 FILLCELL_X1 PHY_5180 ();
 FILLCELL_X1 PHY_5181 ();
 FILLCELL_X1 PHY_5182 ();
 FILLCELL_X1 PHY_5183 ();
 FILLCELL_X1 PHY_5184 ();
 FILLCELL_X1 PHY_5185 ();
 FILLCELL_X1 PHY_5186 ();
 FILLCELL_X1 PHY_5187 ();
 FILLCELL_X1 PHY_5188 ();
 FILLCELL_X1 PHY_5189 ();
 FILLCELL_X1 PHY_519 ();
 FILLCELL_X1 PHY_5190 ();
 FILLCELL_X1 PHY_5191 ();
 FILLCELL_X1 PHY_5192 ();
 FILLCELL_X1 PHY_5193 ();
 FILLCELL_X1 PHY_5194 ();
 FILLCELL_X1 PHY_5195 ();
 FILLCELL_X1 PHY_5196 ();
 FILLCELL_X1 PHY_5197 ();
 FILLCELL_X1 PHY_5198 ();
 FILLCELL_X1 PHY_5199 ();
 FILLCELL_X1 PHY_52 ();
 FILLCELL_X1 PHY_520 ();
 FILLCELL_X1 PHY_5200 ();
 FILLCELL_X1 PHY_5201 ();
 FILLCELL_X1 PHY_5202 ();
 FILLCELL_X1 PHY_5203 ();
 FILLCELL_X1 PHY_5204 ();
 FILLCELL_X1 PHY_5205 ();
 FILLCELL_X1 PHY_5206 ();
 FILLCELL_X1 PHY_5207 ();
 FILLCELL_X1 PHY_5208 ();
 FILLCELL_X1 PHY_5209 ();
 FILLCELL_X1 PHY_521 ();
 FILLCELL_X1 PHY_5210 ();
 FILLCELL_X1 PHY_5211 ();
 FILLCELL_X1 PHY_5212 ();
 FILLCELL_X1 PHY_5213 ();
 FILLCELL_X1 PHY_5214 ();
 FILLCELL_X1 PHY_5215 ();
 FILLCELL_X1 PHY_5216 ();
 FILLCELL_X1 PHY_5217 ();
 FILLCELL_X1 PHY_5218 ();
 FILLCELL_X1 PHY_5219 ();
 FILLCELL_X1 PHY_522 ();
 FILLCELL_X1 PHY_5220 ();
 FILLCELL_X1 PHY_5221 ();
 FILLCELL_X1 PHY_5222 ();
 FILLCELL_X1 PHY_5223 ();
 FILLCELL_X1 PHY_5224 ();
 FILLCELL_X1 PHY_5225 ();
 FILLCELL_X1 PHY_5226 ();
 FILLCELL_X1 PHY_5227 ();
 FILLCELL_X1 PHY_5228 ();
 FILLCELL_X1 PHY_5229 ();
 FILLCELL_X1 PHY_523 ();
 FILLCELL_X1 PHY_5230 ();
 FILLCELL_X1 PHY_5231 ();
 FILLCELL_X1 PHY_5232 ();
 FILLCELL_X1 PHY_5233 ();
 FILLCELL_X1 PHY_5234 ();
 FILLCELL_X1 PHY_5235 ();
 FILLCELL_X1 PHY_5236 ();
 FILLCELL_X1 PHY_5237 ();
 FILLCELL_X1 PHY_5238 ();
 FILLCELL_X1 PHY_5239 ();
 FILLCELL_X1 PHY_524 ();
 FILLCELL_X1 PHY_5240 ();
 FILLCELL_X1 PHY_5241 ();
 FILLCELL_X1 PHY_5242 ();
 FILLCELL_X1 PHY_5243 ();
 FILLCELL_X1 PHY_5244 ();
 FILLCELL_X1 PHY_5245 ();
 FILLCELL_X1 PHY_5246 ();
 FILLCELL_X1 PHY_5247 ();
 FILLCELL_X1 PHY_5248 ();
 FILLCELL_X1 PHY_5249 ();
 FILLCELL_X1 PHY_525 ();
 FILLCELL_X1 PHY_5250 ();
 FILLCELL_X1 PHY_5251 ();
 FILLCELL_X1 PHY_5252 ();
 FILLCELL_X1 PHY_5253 ();
 FILLCELL_X1 PHY_5254 ();
 FILLCELL_X1 PHY_5255 ();
 FILLCELL_X1 PHY_5256 ();
 FILLCELL_X1 PHY_5257 ();
 FILLCELL_X1 PHY_5258 ();
 FILLCELL_X1 PHY_5259 ();
 FILLCELL_X1 PHY_526 ();
 FILLCELL_X1 PHY_5260 ();
 FILLCELL_X1 PHY_5261 ();
 FILLCELL_X1 PHY_5262 ();
 FILLCELL_X1 PHY_5263 ();
 FILLCELL_X1 PHY_5264 ();
 FILLCELL_X1 PHY_5265 ();
 FILLCELL_X1 PHY_5266 ();
 FILLCELL_X1 PHY_5267 ();
 FILLCELL_X1 PHY_5268 ();
 FILLCELL_X1 PHY_5269 ();
 FILLCELL_X1 PHY_527 ();
 FILLCELL_X1 PHY_5270 ();
 FILLCELL_X1 PHY_5271 ();
 FILLCELL_X1 PHY_5272 ();
 FILLCELL_X1 PHY_5273 ();
 FILLCELL_X1 PHY_5274 ();
 FILLCELL_X1 PHY_5275 ();
 FILLCELL_X1 PHY_5276 ();
 FILLCELL_X1 PHY_5277 ();
 FILLCELL_X1 PHY_5278 ();
 FILLCELL_X1 PHY_5279 ();
 FILLCELL_X1 PHY_528 ();
 FILLCELL_X1 PHY_5280 ();
 FILLCELL_X1 PHY_5281 ();
 FILLCELL_X1 PHY_5282 ();
 FILLCELL_X1 PHY_5283 ();
 FILLCELL_X1 PHY_5284 ();
 FILLCELL_X1 PHY_5285 ();
 FILLCELL_X1 PHY_5286 ();
 FILLCELL_X1 PHY_5287 ();
 FILLCELL_X1 PHY_5288 ();
 FILLCELL_X1 PHY_5289 ();
 FILLCELL_X1 PHY_529 ();
 FILLCELL_X1 PHY_5290 ();
 FILLCELL_X1 PHY_5291 ();
 FILLCELL_X1 PHY_5292 ();
 FILLCELL_X1 PHY_5293 ();
 FILLCELL_X1 PHY_5294 ();
 FILLCELL_X1 PHY_5295 ();
 FILLCELL_X1 PHY_5296 ();
 FILLCELL_X1 PHY_5297 ();
 FILLCELL_X1 PHY_5298 ();
 FILLCELL_X1 PHY_5299 ();
 FILLCELL_X1 PHY_53 ();
 FILLCELL_X1 PHY_530 ();
 FILLCELL_X1 PHY_5300 ();
 FILLCELL_X1 PHY_5301 ();
 FILLCELL_X1 PHY_5302 ();
 FILLCELL_X1 PHY_5303 ();
 FILLCELL_X1 PHY_5304 ();
 FILLCELL_X1 PHY_5305 ();
 FILLCELL_X1 PHY_5306 ();
 FILLCELL_X1 PHY_5307 ();
 FILLCELL_X1 PHY_5308 ();
 FILLCELL_X1 PHY_5309 ();
 FILLCELL_X1 PHY_531 ();
 FILLCELL_X1 PHY_5310 ();
 FILLCELL_X1 PHY_5311 ();
 FILLCELL_X1 PHY_5312 ();
 FILLCELL_X1 PHY_5313 ();
 FILLCELL_X1 PHY_5314 ();
 FILLCELL_X1 PHY_5315 ();
 FILLCELL_X1 PHY_5316 ();
 FILLCELL_X1 PHY_5317 ();
 FILLCELL_X1 PHY_5318 ();
 FILLCELL_X1 PHY_5319 ();
 FILLCELL_X1 PHY_532 ();
 FILLCELL_X1 PHY_5320 ();
 FILLCELL_X1 PHY_5321 ();
 FILLCELL_X1 PHY_5322 ();
 FILLCELL_X1 PHY_5323 ();
 FILLCELL_X1 PHY_5324 ();
 FILLCELL_X1 PHY_5325 ();
 FILLCELL_X1 PHY_5326 ();
 FILLCELL_X1 PHY_5327 ();
 FILLCELL_X1 PHY_5328 ();
 FILLCELL_X1 PHY_5329 ();
 FILLCELL_X1 PHY_533 ();
 FILLCELL_X1 PHY_5330 ();
 FILLCELL_X1 PHY_5331 ();
 FILLCELL_X1 PHY_5332 ();
 FILLCELL_X1 PHY_5333 ();
 FILLCELL_X1 PHY_5334 ();
 FILLCELL_X1 PHY_5335 ();
 FILLCELL_X1 PHY_5336 ();
 FILLCELL_X1 PHY_5337 ();
 FILLCELL_X1 PHY_5338 ();
 FILLCELL_X1 PHY_5339 ();
 FILLCELL_X1 PHY_534 ();
 FILLCELL_X1 PHY_5340 ();
 FILLCELL_X1 PHY_5341 ();
 FILLCELL_X1 PHY_5342 ();
 FILLCELL_X1 PHY_5343 ();
 FILLCELL_X1 PHY_5344 ();
 FILLCELL_X1 PHY_5345 ();
 FILLCELL_X1 PHY_5346 ();
 FILLCELL_X1 PHY_5347 ();
 FILLCELL_X1 PHY_5348 ();
 FILLCELL_X1 PHY_5349 ();
 FILLCELL_X1 PHY_535 ();
 FILLCELL_X1 PHY_5350 ();
 FILLCELL_X1 PHY_5351 ();
 FILLCELL_X1 PHY_5352 ();
 FILLCELL_X1 PHY_5353 ();
 FILLCELL_X1 PHY_5354 ();
 FILLCELL_X1 PHY_5355 ();
 FILLCELL_X1 PHY_5356 ();
 FILLCELL_X1 PHY_5357 ();
 FILLCELL_X1 PHY_5358 ();
 FILLCELL_X1 PHY_5359 ();
 FILLCELL_X1 PHY_536 ();
 FILLCELL_X1 PHY_5360 ();
 FILLCELL_X1 PHY_5361 ();
 FILLCELL_X1 PHY_5362 ();
 FILLCELL_X1 PHY_5363 ();
 FILLCELL_X1 PHY_5364 ();
 FILLCELL_X1 PHY_5365 ();
 FILLCELL_X1 PHY_5366 ();
 FILLCELL_X1 PHY_5367 ();
 FILLCELL_X1 PHY_5368 ();
 FILLCELL_X1 PHY_5369 ();
 FILLCELL_X1 PHY_537 ();
 FILLCELL_X1 PHY_5370 ();
 FILLCELL_X1 PHY_5371 ();
 FILLCELL_X1 PHY_5372 ();
 FILLCELL_X1 PHY_5373 ();
 FILLCELL_X1 PHY_5374 ();
 FILLCELL_X1 PHY_5375 ();
 FILLCELL_X1 PHY_5376 ();
 FILLCELL_X1 PHY_5377 ();
 FILLCELL_X1 PHY_5378 ();
 FILLCELL_X1 PHY_5379 ();
 FILLCELL_X1 PHY_538 ();
 FILLCELL_X1 PHY_5380 ();
 FILLCELL_X1 PHY_5381 ();
 FILLCELL_X1 PHY_5382 ();
 FILLCELL_X1 PHY_5383 ();
 FILLCELL_X1 PHY_5384 ();
 FILLCELL_X1 PHY_5385 ();
 FILLCELL_X1 PHY_5386 ();
 FILLCELL_X1 PHY_5387 ();
 FILLCELL_X1 PHY_5388 ();
 FILLCELL_X1 PHY_5389 ();
 FILLCELL_X1 PHY_539 ();
 FILLCELL_X1 PHY_5390 ();
 FILLCELL_X1 PHY_5391 ();
 FILLCELL_X1 PHY_5392 ();
 FILLCELL_X1 PHY_5393 ();
 FILLCELL_X1 PHY_5394 ();
 FILLCELL_X1 PHY_5395 ();
 FILLCELL_X1 PHY_5396 ();
 FILLCELL_X1 PHY_5397 ();
 FILLCELL_X1 PHY_5398 ();
 FILLCELL_X1 PHY_5399 ();
 FILLCELL_X1 PHY_54 ();
 FILLCELL_X1 PHY_540 ();
 FILLCELL_X1 PHY_5400 ();
 FILLCELL_X1 PHY_5401 ();
 FILLCELL_X1 PHY_5402 ();
 FILLCELL_X1 PHY_5403 ();
 FILLCELL_X1 PHY_5404 ();
 FILLCELL_X1 PHY_5405 ();
 FILLCELL_X1 PHY_5406 ();
 FILLCELL_X1 PHY_5407 ();
 FILLCELL_X1 PHY_5408 ();
 FILLCELL_X1 PHY_5409 ();
 FILLCELL_X1 PHY_541 ();
 FILLCELL_X1 PHY_5410 ();
 FILLCELL_X1 PHY_5411 ();
 FILLCELL_X1 PHY_5412 ();
 FILLCELL_X1 PHY_5413 ();
 FILLCELL_X1 PHY_5414 ();
 FILLCELL_X1 PHY_5415 ();
 FILLCELL_X1 PHY_5416 ();
 FILLCELL_X1 PHY_5417 ();
 FILLCELL_X1 PHY_5418 ();
 FILLCELL_X1 PHY_5419 ();
 FILLCELL_X1 PHY_542 ();
 FILLCELL_X1 PHY_5420 ();
 FILLCELL_X1 PHY_5421 ();
 FILLCELL_X1 PHY_5422 ();
 FILLCELL_X1 PHY_5423 ();
 FILLCELL_X1 PHY_5424 ();
 FILLCELL_X1 PHY_5425 ();
 FILLCELL_X1 PHY_5426 ();
 FILLCELL_X1 PHY_5427 ();
 FILLCELL_X1 PHY_5428 ();
 FILLCELL_X1 PHY_5429 ();
 FILLCELL_X1 PHY_543 ();
 FILLCELL_X1 PHY_5430 ();
 FILLCELL_X1 PHY_5431 ();
 FILLCELL_X1 PHY_5432 ();
 FILLCELL_X1 PHY_5433 ();
 FILLCELL_X1 PHY_5434 ();
 FILLCELL_X1 PHY_5435 ();
 FILLCELL_X1 PHY_5436 ();
 FILLCELL_X1 PHY_5437 ();
 FILLCELL_X1 PHY_5438 ();
 FILLCELL_X1 PHY_5439 ();
 FILLCELL_X1 PHY_544 ();
 FILLCELL_X1 PHY_5440 ();
 FILLCELL_X1 PHY_5441 ();
 FILLCELL_X1 PHY_5442 ();
 FILLCELL_X1 PHY_5443 ();
 FILLCELL_X1 PHY_5444 ();
 FILLCELL_X1 PHY_5445 ();
 FILLCELL_X1 PHY_5446 ();
 FILLCELL_X1 PHY_5447 ();
 FILLCELL_X1 PHY_5448 ();
 FILLCELL_X1 PHY_5449 ();
 FILLCELL_X1 PHY_545 ();
 FILLCELL_X1 PHY_5450 ();
 FILLCELL_X1 PHY_5451 ();
 FILLCELL_X1 PHY_5452 ();
 FILLCELL_X1 PHY_5453 ();
 FILLCELL_X1 PHY_5454 ();
 FILLCELL_X1 PHY_5455 ();
 FILLCELL_X1 PHY_5456 ();
 FILLCELL_X1 PHY_5457 ();
 FILLCELL_X1 PHY_5458 ();
 FILLCELL_X1 PHY_5459 ();
 FILLCELL_X1 PHY_546 ();
 FILLCELL_X1 PHY_5460 ();
 FILLCELL_X1 PHY_5461 ();
 FILLCELL_X1 PHY_5462 ();
 FILLCELL_X1 PHY_5463 ();
 FILLCELL_X1 PHY_5464 ();
 FILLCELL_X1 PHY_5465 ();
 FILLCELL_X1 PHY_5466 ();
 FILLCELL_X1 PHY_5467 ();
 FILLCELL_X1 PHY_5468 ();
 FILLCELL_X1 PHY_5469 ();
 FILLCELL_X1 PHY_547 ();
 FILLCELL_X1 PHY_5470 ();
 FILLCELL_X1 PHY_5471 ();
 FILLCELL_X1 PHY_5472 ();
 FILLCELL_X1 PHY_5473 ();
 FILLCELL_X1 PHY_5474 ();
 FILLCELL_X1 PHY_5475 ();
 FILLCELL_X1 PHY_5476 ();
 FILLCELL_X1 PHY_5477 ();
 FILLCELL_X1 PHY_5478 ();
 FILLCELL_X1 PHY_5479 ();
 FILLCELL_X1 PHY_548 ();
 FILLCELL_X1 PHY_5480 ();
 FILLCELL_X1 PHY_5481 ();
 FILLCELL_X1 PHY_5482 ();
 FILLCELL_X1 PHY_5483 ();
 FILLCELL_X1 PHY_5484 ();
 FILLCELL_X1 PHY_5485 ();
 FILLCELL_X1 PHY_5486 ();
 FILLCELL_X1 PHY_5487 ();
 FILLCELL_X1 PHY_5488 ();
 FILLCELL_X1 PHY_5489 ();
 FILLCELL_X1 PHY_549 ();
 FILLCELL_X1 PHY_5490 ();
 FILLCELL_X1 PHY_5491 ();
 FILLCELL_X1 PHY_5492 ();
 FILLCELL_X1 PHY_5493 ();
 FILLCELL_X1 PHY_5494 ();
 FILLCELL_X1 PHY_5495 ();
 FILLCELL_X1 PHY_5496 ();
 FILLCELL_X1 PHY_5497 ();
 FILLCELL_X1 PHY_5498 ();
 FILLCELL_X1 PHY_5499 ();
 FILLCELL_X1 PHY_55 ();
 FILLCELL_X1 PHY_550 ();
 FILLCELL_X1 PHY_5500 ();
 FILLCELL_X1 PHY_5501 ();
 FILLCELL_X1 PHY_5502 ();
 FILLCELL_X1 PHY_5503 ();
 FILLCELL_X1 PHY_5504 ();
 FILLCELL_X1 PHY_5505 ();
 FILLCELL_X1 PHY_5506 ();
 FILLCELL_X1 PHY_5507 ();
 FILLCELL_X1 PHY_5508 ();
 FILLCELL_X1 PHY_5509 ();
 FILLCELL_X1 PHY_551 ();
 FILLCELL_X1 PHY_5510 ();
 FILLCELL_X1 PHY_5511 ();
 FILLCELL_X1 PHY_5512 ();
 FILLCELL_X1 PHY_5513 ();
 FILLCELL_X1 PHY_5514 ();
 FILLCELL_X1 PHY_5515 ();
 FILLCELL_X1 PHY_5516 ();
 FILLCELL_X1 PHY_5517 ();
 FILLCELL_X1 PHY_5518 ();
 FILLCELL_X1 PHY_5519 ();
 FILLCELL_X1 PHY_552 ();
 FILLCELL_X1 PHY_5520 ();
 FILLCELL_X1 PHY_5521 ();
 FILLCELL_X1 PHY_5522 ();
 FILLCELL_X1 PHY_5523 ();
 FILLCELL_X1 PHY_5524 ();
 FILLCELL_X1 PHY_5525 ();
 FILLCELL_X1 PHY_5526 ();
 FILLCELL_X1 PHY_5527 ();
 FILLCELL_X1 PHY_5528 ();
 FILLCELL_X1 PHY_5529 ();
 FILLCELL_X1 PHY_553 ();
 FILLCELL_X1 PHY_5530 ();
 FILLCELL_X1 PHY_5531 ();
 FILLCELL_X1 PHY_5532 ();
 FILLCELL_X1 PHY_5533 ();
 FILLCELL_X1 PHY_5534 ();
 FILLCELL_X1 PHY_5535 ();
 FILLCELL_X1 PHY_5536 ();
 FILLCELL_X1 PHY_5537 ();
 FILLCELL_X1 PHY_5538 ();
 FILLCELL_X1 PHY_5539 ();
 FILLCELL_X1 PHY_554 ();
 FILLCELL_X1 PHY_5540 ();
 FILLCELL_X1 PHY_5541 ();
 FILLCELL_X1 PHY_5542 ();
 FILLCELL_X1 PHY_5543 ();
 FILLCELL_X1 PHY_5544 ();
 FILLCELL_X1 PHY_5545 ();
 FILLCELL_X1 PHY_5546 ();
 FILLCELL_X1 PHY_5547 ();
 FILLCELL_X1 PHY_5548 ();
 FILLCELL_X1 PHY_5549 ();
 FILLCELL_X1 PHY_555 ();
 FILLCELL_X1 PHY_5550 ();
 FILLCELL_X1 PHY_5551 ();
 FILLCELL_X1 PHY_5552 ();
 FILLCELL_X1 PHY_5553 ();
 FILLCELL_X1 PHY_5554 ();
 FILLCELL_X1 PHY_5555 ();
 FILLCELL_X1 PHY_5556 ();
 FILLCELL_X1 PHY_5557 ();
 FILLCELL_X1 PHY_5558 ();
 FILLCELL_X1 PHY_5559 ();
 FILLCELL_X1 PHY_556 ();
 FILLCELL_X1 PHY_5560 ();
 FILLCELL_X1 PHY_5561 ();
 FILLCELL_X1 PHY_5562 ();
 FILLCELL_X1 PHY_5563 ();
 FILLCELL_X1 PHY_5564 ();
 FILLCELL_X1 PHY_5565 ();
 FILLCELL_X1 PHY_5566 ();
 FILLCELL_X1 PHY_5567 ();
 FILLCELL_X1 PHY_5568 ();
 FILLCELL_X1 PHY_5569 ();
 FILLCELL_X1 PHY_557 ();
 FILLCELL_X1 PHY_5570 ();
 FILLCELL_X1 PHY_5571 ();
 FILLCELL_X1 PHY_5572 ();
 FILLCELL_X1 PHY_5573 ();
 FILLCELL_X1 PHY_5574 ();
 FILLCELL_X1 PHY_5575 ();
 FILLCELL_X1 PHY_5576 ();
 FILLCELL_X1 PHY_5577 ();
 FILLCELL_X1 PHY_5578 ();
 FILLCELL_X1 PHY_5579 ();
 FILLCELL_X1 PHY_558 ();
 FILLCELL_X1 PHY_5580 ();
 FILLCELL_X1 PHY_5581 ();
 FILLCELL_X1 PHY_5582 ();
 FILLCELL_X1 PHY_5583 ();
 FILLCELL_X1 PHY_5584 ();
 FILLCELL_X1 PHY_5585 ();
 FILLCELL_X1 PHY_5586 ();
 FILLCELL_X1 PHY_5587 ();
 FILLCELL_X1 PHY_5588 ();
 FILLCELL_X1 PHY_5589 ();
 FILLCELL_X1 PHY_559 ();
 FILLCELL_X1 PHY_5590 ();
 FILLCELL_X1 PHY_5591 ();
 FILLCELL_X1 PHY_5592 ();
 FILLCELL_X1 PHY_5593 ();
 FILLCELL_X1 PHY_5594 ();
 FILLCELL_X1 PHY_5595 ();
 FILLCELL_X1 PHY_5596 ();
 FILLCELL_X1 PHY_5597 ();
 FILLCELL_X1 PHY_5598 ();
 FILLCELL_X1 PHY_5599 ();
 FILLCELL_X1 PHY_56 ();
 FILLCELL_X1 PHY_560 ();
 FILLCELL_X1 PHY_5600 ();
 FILLCELL_X1 PHY_5601 ();
 FILLCELL_X1 PHY_5602 ();
 FILLCELL_X1 PHY_5603 ();
 FILLCELL_X1 PHY_5604 ();
 FILLCELL_X1 PHY_5605 ();
 FILLCELL_X1 PHY_5606 ();
 FILLCELL_X1 PHY_5607 ();
 FILLCELL_X1 PHY_5608 ();
 FILLCELL_X1 PHY_5609 ();
 FILLCELL_X1 PHY_561 ();
 FILLCELL_X1 PHY_5610 ();
 FILLCELL_X1 PHY_5611 ();
 FILLCELL_X1 PHY_5612 ();
 FILLCELL_X1 PHY_5613 ();
 FILLCELL_X1 PHY_5614 ();
 FILLCELL_X1 PHY_5615 ();
 FILLCELL_X1 PHY_5616 ();
 FILLCELL_X1 PHY_5617 ();
 FILLCELL_X1 PHY_5618 ();
 FILLCELL_X1 PHY_5619 ();
 FILLCELL_X1 PHY_562 ();
 FILLCELL_X1 PHY_5620 ();
 FILLCELL_X1 PHY_5621 ();
 FILLCELL_X1 PHY_5622 ();
 FILLCELL_X1 PHY_5623 ();
 FILLCELL_X1 PHY_5624 ();
 FILLCELL_X1 PHY_5625 ();
 FILLCELL_X1 PHY_5626 ();
 FILLCELL_X1 PHY_5627 ();
 FILLCELL_X1 PHY_5628 ();
 FILLCELL_X1 PHY_5629 ();
 FILLCELL_X1 PHY_563 ();
 FILLCELL_X1 PHY_5630 ();
 FILLCELL_X1 PHY_5631 ();
 FILLCELL_X1 PHY_5632 ();
 FILLCELL_X1 PHY_5633 ();
 FILLCELL_X1 PHY_5634 ();
 FILLCELL_X1 PHY_5635 ();
 FILLCELL_X1 PHY_5636 ();
 FILLCELL_X1 PHY_5637 ();
 FILLCELL_X1 PHY_5638 ();
 FILLCELL_X1 PHY_5639 ();
 FILLCELL_X1 PHY_564 ();
 FILLCELL_X1 PHY_5640 ();
 FILLCELL_X1 PHY_5641 ();
 FILLCELL_X1 PHY_5642 ();
 FILLCELL_X1 PHY_5643 ();
 FILLCELL_X1 PHY_5644 ();
 FILLCELL_X1 PHY_5645 ();
 FILLCELL_X1 PHY_5646 ();
 FILLCELL_X1 PHY_5647 ();
 FILLCELL_X1 PHY_5648 ();
 FILLCELL_X1 PHY_5649 ();
 FILLCELL_X1 PHY_565 ();
 FILLCELL_X1 PHY_5650 ();
 FILLCELL_X1 PHY_5651 ();
 FILLCELL_X1 PHY_5652 ();
 FILLCELL_X1 PHY_5653 ();
 FILLCELL_X1 PHY_5654 ();
 FILLCELL_X1 PHY_5655 ();
 FILLCELL_X1 PHY_5656 ();
 FILLCELL_X1 PHY_5657 ();
 FILLCELL_X1 PHY_5658 ();
 FILLCELL_X1 PHY_5659 ();
 FILLCELL_X1 PHY_566 ();
 FILLCELL_X1 PHY_5660 ();
 FILLCELL_X1 PHY_5661 ();
 FILLCELL_X1 PHY_5662 ();
 FILLCELL_X1 PHY_5663 ();
 FILLCELL_X1 PHY_5664 ();
 FILLCELL_X1 PHY_5665 ();
 FILLCELL_X1 PHY_5666 ();
 FILLCELL_X1 PHY_5667 ();
 FILLCELL_X1 PHY_5668 ();
 FILLCELL_X1 PHY_5669 ();
 FILLCELL_X1 PHY_567 ();
 FILLCELL_X1 PHY_5670 ();
 FILLCELL_X1 PHY_5671 ();
 FILLCELL_X1 PHY_5672 ();
 FILLCELL_X1 PHY_5673 ();
 FILLCELL_X1 PHY_5674 ();
 FILLCELL_X1 PHY_5675 ();
 FILLCELL_X1 PHY_5676 ();
 FILLCELL_X1 PHY_5677 ();
 FILLCELL_X1 PHY_5678 ();
 FILLCELL_X1 PHY_5679 ();
 FILLCELL_X1 PHY_568 ();
 FILLCELL_X1 PHY_5680 ();
 FILLCELL_X1 PHY_5681 ();
 FILLCELL_X1 PHY_5682 ();
 FILLCELL_X1 PHY_5683 ();
 FILLCELL_X1 PHY_5684 ();
 FILLCELL_X1 PHY_5685 ();
 FILLCELL_X1 PHY_5686 ();
 FILLCELL_X1 PHY_5687 ();
 FILLCELL_X1 PHY_5688 ();
 FILLCELL_X1 PHY_5689 ();
 FILLCELL_X1 PHY_569 ();
 FILLCELL_X1 PHY_5690 ();
 FILLCELL_X1 PHY_5691 ();
 FILLCELL_X1 PHY_5692 ();
 FILLCELL_X1 PHY_5693 ();
 FILLCELL_X1 PHY_5694 ();
 FILLCELL_X1 PHY_5695 ();
 FILLCELL_X1 PHY_5696 ();
 FILLCELL_X1 PHY_5697 ();
 FILLCELL_X1 PHY_5698 ();
 FILLCELL_X1 PHY_5699 ();
 FILLCELL_X1 PHY_57 ();
 FILLCELL_X1 PHY_570 ();
 FILLCELL_X1 PHY_5700 ();
 FILLCELL_X1 PHY_5701 ();
 FILLCELL_X1 PHY_5702 ();
 FILLCELL_X1 PHY_5703 ();
 FILLCELL_X1 PHY_5704 ();
 FILLCELL_X1 PHY_5705 ();
 FILLCELL_X1 PHY_5706 ();
 FILLCELL_X1 PHY_5707 ();
 FILLCELL_X1 PHY_5708 ();
 FILLCELL_X1 PHY_5709 ();
 FILLCELL_X1 PHY_571 ();
 FILLCELL_X1 PHY_5710 ();
 FILLCELL_X1 PHY_5711 ();
 FILLCELL_X1 PHY_5712 ();
 FILLCELL_X1 PHY_5713 ();
 FILLCELL_X1 PHY_5714 ();
 FILLCELL_X1 PHY_5715 ();
 FILLCELL_X1 PHY_5716 ();
 FILLCELL_X1 PHY_5717 ();
 FILLCELL_X1 PHY_5718 ();
 FILLCELL_X1 PHY_5719 ();
 FILLCELL_X1 PHY_572 ();
 FILLCELL_X1 PHY_5720 ();
 FILLCELL_X1 PHY_5721 ();
 FILLCELL_X1 PHY_5722 ();
 FILLCELL_X1 PHY_5723 ();
 FILLCELL_X1 PHY_5724 ();
 FILLCELL_X1 PHY_5725 ();
 FILLCELL_X1 PHY_5726 ();
 FILLCELL_X1 PHY_5727 ();
 FILLCELL_X1 PHY_5728 ();
 FILLCELL_X1 PHY_5729 ();
 FILLCELL_X1 PHY_573 ();
 FILLCELL_X1 PHY_5730 ();
 FILLCELL_X1 PHY_5731 ();
 FILLCELL_X1 PHY_5732 ();
 FILLCELL_X1 PHY_5733 ();
 FILLCELL_X1 PHY_5734 ();
 FILLCELL_X1 PHY_5735 ();
 FILLCELL_X1 PHY_5736 ();
 FILLCELL_X1 PHY_5737 ();
 FILLCELL_X1 PHY_5738 ();
 FILLCELL_X1 PHY_5739 ();
 FILLCELL_X1 PHY_574 ();
 FILLCELL_X1 PHY_5740 ();
 FILLCELL_X1 PHY_5741 ();
 FILLCELL_X1 PHY_5742 ();
 FILLCELL_X1 PHY_5743 ();
 FILLCELL_X1 PHY_5744 ();
 FILLCELL_X1 PHY_5745 ();
 FILLCELL_X1 PHY_5746 ();
 FILLCELL_X1 PHY_5747 ();
 FILLCELL_X1 PHY_5748 ();
 FILLCELL_X1 PHY_5749 ();
 FILLCELL_X1 PHY_575 ();
 FILLCELL_X1 PHY_5750 ();
 FILLCELL_X1 PHY_5751 ();
 FILLCELL_X1 PHY_5752 ();
 FILLCELL_X1 PHY_5753 ();
 FILLCELL_X1 PHY_5754 ();
 FILLCELL_X1 PHY_5755 ();
 FILLCELL_X1 PHY_5756 ();
 FILLCELL_X1 PHY_5757 ();
 FILLCELL_X1 PHY_5758 ();
 FILLCELL_X1 PHY_5759 ();
 FILLCELL_X1 PHY_576 ();
 FILLCELL_X1 PHY_5760 ();
 FILLCELL_X1 PHY_5761 ();
 FILLCELL_X1 PHY_5762 ();
 FILLCELL_X1 PHY_5763 ();
 FILLCELL_X1 PHY_5764 ();
 FILLCELL_X1 PHY_5765 ();
 FILLCELL_X1 PHY_5766 ();
 FILLCELL_X1 PHY_5767 ();
 FILLCELL_X1 PHY_5768 ();
 FILLCELL_X1 PHY_5769 ();
 FILLCELL_X1 PHY_577 ();
 FILLCELL_X1 PHY_5770 ();
 FILLCELL_X1 PHY_5771 ();
 FILLCELL_X1 PHY_5772 ();
 FILLCELL_X1 PHY_5773 ();
 FILLCELL_X1 PHY_5774 ();
 FILLCELL_X1 PHY_5775 ();
 FILLCELL_X1 PHY_5776 ();
 FILLCELL_X1 PHY_5777 ();
 FILLCELL_X1 PHY_5778 ();
 FILLCELL_X1 PHY_5779 ();
 FILLCELL_X1 PHY_578 ();
 FILLCELL_X1 PHY_5780 ();
 FILLCELL_X1 PHY_5781 ();
 FILLCELL_X1 PHY_5782 ();
 FILLCELL_X1 PHY_5783 ();
 FILLCELL_X1 PHY_5784 ();
 FILLCELL_X1 PHY_5785 ();
 FILLCELL_X1 PHY_5786 ();
 FILLCELL_X1 PHY_5787 ();
 FILLCELL_X1 PHY_5788 ();
 FILLCELL_X1 PHY_5789 ();
 FILLCELL_X1 PHY_579 ();
 FILLCELL_X1 PHY_5790 ();
 FILLCELL_X1 PHY_5791 ();
 FILLCELL_X1 PHY_5792 ();
 FILLCELL_X1 PHY_5793 ();
 FILLCELL_X1 PHY_5794 ();
 FILLCELL_X1 PHY_5795 ();
 FILLCELL_X1 PHY_5796 ();
 FILLCELL_X1 PHY_5797 ();
 FILLCELL_X1 PHY_5798 ();
 FILLCELL_X1 PHY_5799 ();
 FILLCELL_X1 PHY_58 ();
 FILLCELL_X1 PHY_580 ();
 FILLCELL_X1 PHY_5800 ();
 FILLCELL_X1 PHY_5801 ();
 FILLCELL_X1 PHY_5802 ();
 FILLCELL_X1 PHY_5803 ();
 FILLCELL_X1 PHY_5804 ();
 FILLCELL_X1 PHY_5805 ();
 FILLCELL_X1 PHY_5806 ();
 FILLCELL_X1 PHY_5807 ();
 FILLCELL_X1 PHY_5808 ();
 FILLCELL_X1 PHY_5809 ();
 FILLCELL_X1 PHY_581 ();
 FILLCELL_X1 PHY_5810 ();
 FILLCELL_X1 PHY_5811 ();
 FILLCELL_X1 PHY_5812 ();
 FILLCELL_X1 PHY_5813 ();
 FILLCELL_X1 PHY_5814 ();
 FILLCELL_X1 PHY_5815 ();
 FILLCELL_X1 PHY_5816 ();
 FILLCELL_X1 PHY_5817 ();
 FILLCELL_X1 PHY_5818 ();
 FILLCELL_X1 PHY_5819 ();
 FILLCELL_X1 PHY_582 ();
 FILLCELL_X1 PHY_5820 ();
 FILLCELL_X1 PHY_5821 ();
 FILLCELL_X1 PHY_5822 ();
 FILLCELL_X1 PHY_5823 ();
 FILLCELL_X1 PHY_5824 ();
 FILLCELL_X1 PHY_5825 ();
 FILLCELL_X1 PHY_5826 ();
 FILLCELL_X1 PHY_5827 ();
 FILLCELL_X1 PHY_5828 ();
 FILLCELL_X1 PHY_5829 ();
 FILLCELL_X1 PHY_583 ();
 FILLCELL_X1 PHY_5830 ();
 FILLCELL_X1 PHY_5831 ();
 FILLCELL_X1 PHY_5832 ();
 FILLCELL_X1 PHY_5833 ();
 FILLCELL_X1 PHY_5834 ();
 FILLCELL_X1 PHY_5835 ();
 FILLCELL_X1 PHY_5836 ();
 FILLCELL_X1 PHY_5837 ();
 FILLCELL_X1 PHY_5838 ();
 FILLCELL_X1 PHY_5839 ();
 FILLCELL_X1 PHY_584 ();
 FILLCELL_X1 PHY_5840 ();
 FILLCELL_X1 PHY_5841 ();
 FILLCELL_X1 PHY_5842 ();
 FILLCELL_X1 PHY_5843 ();
 FILLCELL_X1 PHY_5844 ();
 FILLCELL_X1 PHY_5845 ();
 FILLCELL_X1 PHY_5846 ();
 FILLCELL_X1 PHY_5847 ();
 FILLCELL_X1 PHY_5848 ();
 FILLCELL_X1 PHY_5849 ();
 FILLCELL_X1 PHY_585 ();
 FILLCELL_X1 PHY_5850 ();
 FILLCELL_X1 PHY_5851 ();
 FILLCELL_X1 PHY_5852 ();
 FILLCELL_X1 PHY_5853 ();
 FILLCELL_X1 PHY_5854 ();
 FILLCELL_X1 PHY_5855 ();
 FILLCELL_X1 PHY_5856 ();
 FILLCELL_X1 PHY_5857 ();
 FILLCELL_X1 PHY_5858 ();
 FILLCELL_X1 PHY_5859 ();
 FILLCELL_X1 PHY_586 ();
 FILLCELL_X1 PHY_5860 ();
 FILLCELL_X1 PHY_5861 ();
 FILLCELL_X1 PHY_5862 ();
 FILLCELL_X1 PHY_5863 ();
 FILLCELL_X1 PHY_5864 ();
 FILLCELL_X1 PHY_5865 ();
 FILLCELL_X1 PHY_5866 ();
 FILLCELL_X1 PHY_5867 ();
 FILLCELL_X1 PHY_5868 ();
 FILLCELL_X1 PHY_5869 ();
 FILLCELL_X1 PHY_587 ();
 FILLCELL_X1 PHY_5870 ();
 FILLCELL_X1 PHY_5871 ();
 FILLCELL_X1 PHY_5872 ();
 FILLCELL_X1 PHY_5873 ();
 FILLCELL_X1 PHY_5874 ();
 FILLCELL_X1 PHY_5875 ();
 FILLCELL_X1 PHY_5876 ();
 FILLCELL_X1 PHY_5877 ();
 FILLCELL_X1 PHY_5878 ();
 FILLCELL_X1 PHY_5879 ();
 FILLCELL_X1 PHY_588 ();
 FILLCELL_X1 PHY_5880 ();
 FILLCELL_X1 PHY_5881 ();
 FILLCELL_X1 PHY_5882 ();
 FILLCELL_X1 PHY_5883 ();
 FILLCELL_X1 PHY_5884 ();
 FILLCELL_X1 PHY_5885 ();
 FILLCELL_X1 PHY_5886 ();
 FILLCELL_X1 PHY_5887 ();
 FILLCELL_X1 PHY_5888 ();
 FILLCELL_X1 PHY_5889 ();
 FILLCELL_X1 PHY_589 ();
 FILLCELL_X1 PHY_5890 ();
 FILLCELL_X1 PHY_5891 ();
 FILLCELL_X1 PHY_5892 ();
 FILLCELL_X1 PHY_5893 ();
 FILLCELL_X1 PHY_5894 ();
 FILLCELL_X1 PHY_5895 ();
 FILLCELL_X1 PHY_5896 ();
 FILLCELL_X1 PHY_5897 ();
 FILLCELL_X1 PHY_5898 ();
 FILLCELL_X1 PHY_5899 ();
 FILLCELL_X1 PHY_59 ();
 FILLCELL_X1 PHY_590 ();
 FILLCELL_X1 PHY_5900 ();
 FILLCELL_X1 PHY_5901 ();
 FILLCELL_X1 PHY_5902 ();
 FILLCELL_X1 PHY_5903 ();
 FILLCELL_X1 PHY_5904 ();
 FILLCELL_X1 PHY_5905 ();
 FILLCELL_X1 PHY_5906 ();
 FILLCELL_X1 PHY_5907 ();
 FILLCELL_X1 PHY_5908 ();
 FILLCELL_X1 PHY_5909 ();
 FILLCELL_X1 PHY_591 ();
 FILLCELL_X1 PHY_5910 ();
 FILLCELL_X1 PHY_5911 ();
 FILLCELL_X1 PHY_5912 ();
 FILLCELL_X1 PHY_5913 ();
 FILLCELL_X1 PHY_5914 ();
 FILLCELL_X1 PHY_5915 ();
 FILLCELL_X1 PHY_5916 ();
 FILLCELL_X1 PHY_5917 ();
 FILLCELL_X1 PHY_5918 ();
 FILLCELL_X1 PHY_5919 ();
 FILLCELL_X1 PHY_592 ();
 FILLCELL_X1 PHY_5920 ();
 FILLCELL_X1 PHY_5921 ();
 FILLCELL_X1 PHY_5922 ();
 FILLCELL_X1 PHY_5923 ();
 FILLCELL_X1 PHY_5924 ();
 FILLCELL_X1 PHY_5925 ();
 FILLCELL_X1 PHY_5926 ();
 FILLCELL_X1 PHY_5927 ();
 FILLCELL_X1 PHY_5928 ();
 FILLCELL_X1 PHY_5929 ();
 FILLCELL_X1 PHY_593 ();
 FILLCELL_X1 PHY_5930 ();
 FILLCELL_X1 PHY_5931 ();
 FILLCELL_X1 PHY_5932 ();
 FILLCELL_X1 PHY_5933 ();
 FILLCELL_X1 PHY_5934 ();
 FILLCELL_X1 PHY_5935 ();
 FILLCELL_X1 PHY_5936 ();
 FILLCELL_X1 PHY_5937 ();
 FILLCELL_X1 PHY_5938 ();
 FILLCELL_X1 PHY_5939 ();
 FILLCELL_X1 PHY_594 ();
 FILLCELL_X1 PHY_5940 ();
 FILLCELL_X1 PHY_5941 ();
 FILLCELL_X1 PHY_5942 ();
 FILLCELL_X1 PHY_5943 ();
 FILLCELL_X1 PHY_5944 ();
 FILLCELL_X1 PHY_5945 ();
 FILLCELL_X1 PHY_5946 ();
 FILLCELL_X1 PHY_5947 ();
 FILLCELL_X1 PHY_5948 ();
 FILLCELL_X1 PHY_5949 ();
 FILLCELL_X1 PHY_595 ();
 FILLCELL_X1 PHY_5950 ();
 FILLCELL_X1 PHY_5951 ();
 FILLCELL_X1 PHY_5952 ();
 FILLCELL_X1 PHY_5953 ();
 FILLCELL_X1 PHY_5954 ();
 FILLCELL_X1 PHY_5955 ();
 FILLCELL_X1 PHY_5956 ();
 FILLCELL_X1 PHY_5957 ();
 FILLCELL_X1 PHY_5958 ();
 FILLCELL_X1 PHY_5959 ();
 FILLCELL_X1 PHY_596 ();
 FILLCELL_X1 PHY_5960 ();
 FILLCELL_X1 PHY_5961 ();
 FILLCELL_X1 PHY_5962 ();
 FILLCELL_X1 PHY_5963 ();
 FILLCELL_X1 PHY_5964 ();
 FILLCELL_X1 PHY_5965 ();
 FILLCELL_X1 PHY_5966 ();
 FILLCELL_X1 PHY_5967 ();
 FILLCELL_X1 PHY_5968 ();
 FILLCELL_X1 PHY_5969 ();
 FILLCELL_X1 PHY_597 ();
 FILLCELL_X1 PHY_5970 ();
 FILLCELL_X1 PHY_5971 ();
 FILLCELL_X1 PHY_5972 ();
 FILLCELL_X1 PHY_5973 ();
 FILLCELL_X1 PHY_5974 ();
 FILLCELL_X1 PHY_5975 ();
 FILLCELL_X1 PHY_5976 ();
 FILLCELL_X1 PHY_5977 ();
 FILLCELL_X1 PHY_5978 ();
 FILLCELL_X1 PHY_5979 ();
 FILLCELL_X1 PHY_598 ();
 FILLCELL_X1 PHY_5980 ();
 FILLCELL_X1 PHY_5981 ();
 FILLCELL_X1 PHY_5982 ();
 FILLCELL_X1 PHY_5983 ();
 FILLCELL_X1 PHY_5984 ();
 FILLCELL_X1 PHY_5985 ();
 FILLCELL_X1 PHY_5986 ();
 FILLCELL_X1 PHY_5987 ();
 FILLCELL_X1 PHY_5988 ();
 FILLCELL_X1 PHY_5989 ();
 FILLCELL_X1 PHY_599 ();
 FILLCELL_X1 PHY_5990 ();
 FILLCELL_X1 PHY_5991 ();
 FILLCELL_X1 PHY_5992 ();
 FILLCELL_X1 PHY_5993 ();
 FILLCELL_X1 PHY_5994 ();
 FILLCELL_X1 PHY_5995 ();
 FILLCELL_X1 PHY_5996 ();
 FILLCELL_X1 PHY_5997 ();
 FILLCELL_X1 PHY_5998 ();
 FILLCELL_X1 PHY_5999 ();
 FILLCELL_X1 PHY_6 ();
 FILLCELL_X1 PHY_60 ();
 FILLCELL_X1 PHY_600 ();
 FILLCELL_X1 PHY_6000 ();
 FILLCELL_X1 PHY_6001 ();
 FILLCELL_X1 PHY_6002 ();
 FILLCELL_X1 PHY_6003 ();
 FILLCELL_X1 PHY_6004 ();
 FILLCELL_X1 PHY_6005 ();
 FILLCELL_X1 PHY_6006 ();
 FILLCELL_X1 PHY_6007 ();
 FILLCELL_X1 PHY_6008 ();
 FILLCELL_X1 PHY_6009 ();
 FILLCELL_X1 PHY_601 ();
 FILLCELL_X1 PHY_6010 ();
 FILLCELL_X1 PHY_6011 ();
 FILLCELL_X1 PHY_6012 ();
 FILLCELL_X1 PHY_6013 ();
 FILLCELL_X1 PHY_6014 ();
 FILLCELL_X1 PHY_6015 ();
 FILLCELL_X1 PHY_6016 ();
 FILLCELL_X1 PHY_6017 ();
 FILLCELL_X1 PHY_6018 ();
 FILLCELL_X1 PHY_6019 ();
 FILLCELL_X1 PHY_602 ();
 FILLCELL_X1 PHY_6020 ();
 FILLCELL_X1 PHY_6021 ();
 FILLCELL_X1 PHY_6022 ();
 FILLCELL_X1 PHY_6023 ();
 FILLCELL_X1 PHY_6024 ();
 FILLCELL_X1 PHY_6025 ();
 FILLCELL_X1 PHY_6026 ();
 FILLCELL_X1 PHY_6027 ();
 FILLCELL_X1 PHY_6028 ();
 FILLCELL_X1 PHY_6029 ();
 FILLCELL_X1 PHY_603 ();
 FILLCELL_X1 PHY_6030 ();
 FILLCELL_X1 PHY_6031 ();
 FILLCELL_X1 PHY_6032 ();
 FILLCELL_X1 PHY_6033 ();
 FILLCELL_X1 PHY_6034 ();
 FILLCELL_X1 PHY_6035 ();
 FILLCELL_X1 PHY_6036 ();
 FILLCELL_X1 PHY_6037 ();
 FILLCELL_X1 PHY_6038 ();
 FILLCELL_X1 PHY_6039 ();
 FILLCELL_X1 PHY_604 ();
 FILLCELL_X1 PHY_6040 ();
 FILLCELL_X1 PHY_6041 ();
 FILLCELL_X1 PHY_6042 ();
 FILLCELL_X1 PHY_6043 ();
 FILLCELL_X1 PHY_6044 ();
 FILLCELL_X1 PHY_6045 ();
 FILLCELL_X1 PHY_6046 ();
 FILLCELL_X1 PHY_6047 ();
 FILLCELL_X1 PHY_6048 ();
 FILLCELL_X1 PHY_6049 ();
 FILLCELL_X1 PHY_605 ();
 FILLCELL_X1 PHY_6050 ();
 FILLCELL_X1 PHY_6051 ();
 FILLCELL_X1 PHY_6052 ();
 FILLCELL_X1 PHY_6053 ();
 FILLCELL_X1 PHY_6054 ();
 FILLCELL_X1 PHY_6055 ();
 FILLCELL_X1 PHY_6056 ();
 FILLCELL_X1 PHY_6057 ();
 FILLCELL_X1 PHY_6058 ();
 FILLCELL_X1 PHY_6059 ();
 FILLCELL_X1 PHY_606 ();
 FILLCELL_X1 PHY_6060 ();
 FILLCELL_X1 PHY_6061 ();
 FILLCELL_X1 PHY_6062 ();
 FILLCELL_X1 PHY_6063 ();
 FILLCELL_X1 PHY_6064 ();
 FILLCELL_X1 PHY_6065 ();
 FILLCELL_X1 PHY_6066 ();
 FILLCELL_X1 PHY_6067 ();
 FILLCELL_X1 PHY_6068 ();
 FILLCELL_X1 PHY_6069 ();
 FILLCELL_X1 PHY_607 ();
 FILLCELL_X1 PHY_6070 ();
 FILLCELL_X1 PHY_6071 ();
 FILLCELL_X1 PHY_6072 ();
 FILLCELL_X1 PHY_6073 ();
 FILLCELL_X1 PHY_6074 ();
 FILLCELL_X1 PHY_6075 ();
 FILLCELL_X1 PHY_6076 ();
 FILLCELL_X1 PHY_6077 ();
 FILLCELL_X1 PHY_6078 ();
 FILLCELL_X1 PHY_6079 ();
 FILLCELL_X1 PHY_608 ();
 FILLCELL_X1 PHY_6080 ();
 FILLCELL_X1 PHY_6081 ();
 FILLCELL_X1 PHY_6082 ();
 FILLCELL_X1 PHY_6083 ();
 FILLCELL_X1 PHY_6084 ();
 FILLCELL_X1 PHY_6085 ();
 FILLCELL_X1 PHY_6086 ();
 FILLCELL_X1 PHY_6087 ();
 FILLCELL_X1 PHY_6088 ();
 FILLCELL_X1 PHY_6089 ();
 FILLCELL_X1 PHY_609 ();
 FILLCELL_X1 PHY_6090 ();
 FILLCELL_X1 PHY_6091 ();
 FILLCELL_X1 PHY_6092 ();
 FILLCELL_X1 PHY_6093 ();
 FILLCELL_X1 PHY_6094 ();
 FILLCELL_X1 PHY_6095 ();
 FILLCELL_X1 PHY_6096 ();
 FILLCELL_X1 PHY_6097 ();
 FILLCELL_X1 PHY_6098 ();
 FILLCELL_X1 PHY_6099 ();
 FILLCELL_X1 PHY_61 ();
 FILLCELL_X1 PHY_610 ();
 FILLCELL_X1 PHY_6100 ();
 FILLCELL_X1 PHY_6101 ();
 FILLCELL_X1 PHY_6102 ();
 FILLCELL_X1 PHY_6103 ();
 FILLCELL_X1 PHY_6104 ();
 FILLCELL_X1 PHY_6105 ();
 FILLCELL_X1 PHY_6106 ();
 FILLCELL_X1 PHY_6107 ();
 FILLCELL_X1 PHY_6108 ();
 FILLCELL_X1 PHY_6109 ();
 FILLCELL_X1 PHY_611 ();
 FILLCELL_X1 PHY_6110 ();
 FILLCELL_X1 PHY_6111 ();
 FILLCELL_X1 PHY_6112 ();
 FILLCELL_X1 PHY_6113 ();
 FILLCELL_X1 PHY_6114 ();
 FILLCELL_X1 PHY_6115 ();
 FILLCELL_X1 PHY_6116 ();
 FILLCELL_X1 PHY_6117 ();
 FILLCELL_X1 PHY_6118 ();
 FILLCELL_X1 PHY_6119 ();
 FILLCELL_X1 PHY_612 ();
 FILLCELL_X1 PHY_6120 ();
 FILLCELL_X1 PHY_6121 ();
 FILLCELL_X1 PHY_6122 ();
 FILLCELL_X1 PHY_6123 ();
 FILLCELL_X1 PHY_6124 ();
 FILLCELL_X1 PHY_6125 ();
 FILLCELL_X1 PHY_6126 ();
 FILLCELL_X1 PHY_6127 ();
 FILLCELL_X1 PHY_6128 ();
 FILLCELL_X1 PHY_6129 ();
 FILLCELL_X1 PHY_613 ();
 FILLCELL_X1 PHY_6130 ();
 FILLCELL_X1 PHY_6131 ();
 FILLCELL_X1 PHY_6132 ();
 FILLCELL_X1 PHY_6133 ();
 FILLCELL_X1 PHY_6134 ();
 FILLCELL_X1 PHY_6135 ();
 FILLCELL_X1 PHY_6136 ();
 FILLCELL_X1 PHY_6137 ();
 FILLCELL_X1 PHY_6138 ();
 FILLCELL_X1 PHY_6139 ();
 FILLCELL_X1 PHY_614 ();
 FILLCELL_X1 PHY_6140 ();
 FILLCELL_X1 PHY_6141 ();
 FILLCELL_X1 PHY_6142 ();
 FILLCELL_X1 PHY_6143 ();
 FILLCELL_X1 PHY_6144 ();
 FILLCELL_X1 PHY_6145 ();
 FILLCELL_X1 PHY_6146 ();
 FILLCELL_X1 PHY_6147 ();
 FILLCELL_X1 PHY_6148 ();
 FILLCELL_X1 PHY_6149 ();
 FILLCELL_X1 PHY_615 ();
 FILLCELL_X1 PHY_6150 ();
 FILLCELL_X1 PHY_6151 ();
 FILLCELL_X1 PHY_6152 ();
 FILLCELL_X1 PHY_6153 ();
 FILLCELL_X1 PHY_6154 ();
 FILLCELL_X1 PHY_6155 ();
 FILLCELL_X1 PHY_6156 ();
 FILLCELL_X1 PHY_6157 ();
 FILLCELL_X1 PHY_6158 ();
 FILLCELL_X1 PHY_6159 ();
 FILLCELL_X1 PHY_616 ();
 FILLCELL_X1 PHY_6160 ();
 FILLCELL_X1 PHY_6161 ();
 FILLCELL_X1 PHY_6162 ();
 FILLCELL_X1 PHY_6163 ();
 FILLCELL_X1 PHY_6164 ();
 FILLCELL_X1 PHY_6165 ();
 FILLCELL_X1 PHY_6166 ();
 FILLCELL_X1 PHY_6167 ();
 FILLCELL_X1 PHY_6168 ();
 FILLCELL_X1 PHY_6169 ();
 FILLCELL_X1 PHY_617 ();
 FILLCELL_X1 PHY_6170 ();
 FILLCELL_X1 PHY_6171 ();
 FILLCELL_X1 PHY_6172 ();
 FILLCELL_X1 PHY_6173 ();
 FILLCELL_X1 PHY_6174 ();
 FILLCELL_X1 PHY_6175 ();
 FILLCELL_X1 PHY_6176 ();
 FILLCELL_X1 PHY_6177 ();
 FILLCELL_X1 PHY_6178 ();
 FILLCELL_X1 PHY_6179 ();
 FILLCELL_X1 PHY_618 ();
 FILLCELL_X1 PHY_6180 ();
 FILLCELL_X1 PHY_6181 ();
 FILLCELL_X1 PHY_6182 ();
 FILLCELL_X1 PHY_6183 ();
 FILLCELL_X1 PHY_6184 ();
 FILLCELL_X1 PHY_6185 ();
 FILLCELL_X1 PHY_6186 ();
 FILLCELL_X1 PHY_6187 ();
 FILLCELL_X1 PHY_6188 ();
 FILLCELL_X1 PHY_6189 ();
 FILLCELL_X1 PHY_619 ();
 FILLCELL_X1 PHY_6190 ();
 FILLCELL_X1 PHY_6191 ();
 FILLCELL_X1 PHY_6192 ();
 FILLCELL_X1 PHY_6193 ();
 FILLCELL_X1 PHY_6194 ();
 FILLCELL_X1 PHY_6195 ();
 FILLCELL_X1 PHY_6196 ();
 FILLCELL_X1 PHY_6197 ();
 FILLCELL_X1 PHY_6198 ();
 FILLCELL_X1 PHY_6199 ();
 FILLCELL_X1 PHY_62 ();
 FILLCELL_X1 PHY_620 ();
 FILLCELL_X1 PHY_6200 ();
 FILLCELL_X1 PHY_6201 ();
 FILLCELL_X1 PHY_6202 ();
 FILLCELL_X1 PHY_6203 ();
 FILLCELL_X1 PHY_6204 ();
 FILLCELL_X1 PHY_6205 ();
 FILLCELL_X1 PHY_6206 ();
 FILLCELL_X1 PHY_6207 ();
 FILLCELL_X1 PHY_6208 ();
 FILLCELL_X1 PHY_6209 ();
 FILLCELL_X1 PHY_621 ();
 FILLCELL_X1 PHY_6210 ();
 FILLCELL_X1 PHY_6211 ();
 FILLCELL_X1 PHY_6212 ();
 FILLCELL_X1 PHY_6213 ();
 FILLCELL_X1 PHY_6214 ();
 FILLCELL_X1 PHY_6215 ();
 FILLCELL_X1 PHY_6216 ();
 FILLCELL_X1 PHY_6217 ();
 FILLCELL_X1 PHY_6218 ();
 FILLCELL_X1 PHY_6219 ();
 FILLCELL_X1 PHY_622 ();
 FILLCELL_X1 PHY_6220 ();
 FILLCELL_X1 PHY_6221 ();
 FILLCELL_X1 PHY_6222 ();
 FILLCELL_X1 PHY_6223 ();
 FILLCELL_X1 PHY_6224 ();
 FILLCELL_X1 PHY_6225 ();
 FILLCELL_X1 PHY_6226 ();
 FILLCELL_X1 PHY_6227 ();
 FILLCELL_X1 PHY_6228 ();
 FILLCELL_X1 PHY_6229 ();
 FILLCELL_X1 PHY_623 ();
 FILLCELL_X1 PHY_6230 ();
 FILLCELL_X1 PHY_6231 ();
 FILLCELL_X1 PHY_6232 ();
 FILLCELL_X1 PHY_6233 ();
 FILLCELL_X1 PHY_6234 ();
 FILLCELL_X1 PHY_6235 ();
 FILLCELL_X1 PHY_6236 ();
 FILLCELL_X1 PHY_6237 ();
 FILLCELL_X1 PHY_6238 ();
 FILLCELL_X1 PHY_6239 ();
 FILLCELL_X1 PHY_624 ();
 FILLCELL_X1 PHY_6240 ();
 FILLCELL_X1 PHY_6241 ();
 FILLCELL_X1 PHY_6242 ();
 FILLCELL_X1 PHY_6243 ();
 FILLCELL_X1 PHY_6244 ();
 FILLCELL_X1 PHY_6245 ();
 FILLCELL_X1 PHY_6246 ();
 FILLCELL_X1 PHY_6247 ();
 FILLCELL_X1 PHY_6248 ();
 FILLCELL_X1 PHY_6249 ();
 FILLCELL_X1 PHY_625 ();
 FILLCELL_X1 PHY_6250 ();
 FILLCELL_X1 PHY_6251 ();
 FILLCELL_X1 PHY_6252 ();
 FILLCELL_X1 PHY_6253 ();
 FILLCELL_X1 PHY_6254 ();
 FILLCELL_X1 PHY_6255 ();
 FILLCELL_X1 PHY_6256 ();
 FILLCELL_X1 PHY_6257 ();
 FILLCELL_X1 PHY_6258 ();
 FILLCELL_X1 PHY_6259 ();
 FILLCELL_X1 PHY_626 ();
 FILLCELL_X1 PHY_6260 ();
 FILLCELL_X1 PHY_6261 ();
 FILLCELL_X1 PHY_6262 ();
 FILLCELL_X1 PHY_6263 ();
 FILLCELL_X1 PHY_6264 ();
 FILLCELL_X1 PHY_6265 ();
 FILLCELL_X1 PHY_6266 ();
 FILLCELL_X1 PHY_6267 ();
 FILLCELL_X1 PHY_6268 ();
 FILLCELL_X1 PHY_6269 ();
 FILLCELL_X1 PHY_627 ();
 FILLCELL_X1 PHY_6270 ();
 FILLCELL_X1 PHY_6271 ();
 FILLCELL_X1 PHY_6272 ();
 FILLCELL_X1 PHY_6273 ();
 FILLCELL_X1 PHY_6274 ();
 FILLCELL_X1 PHY_6275 ();
 FILLCELL_X1 PHY_6276 ();
 FILLCELL_X1 PHY_6277 ();
 FILLCELL_X1 PHY_6278 ();
 FILLCELL_X1 PHY_6279 ();
 FILLCELL_X1 PHY_628 ();
 FILLCELL_X1 PHY_6280 ();
 FILLCELL_X1 PHY_6281 ();
 FILLCELL_X1 PHY_6282 ();
 FILLCELL_X1 PHY_6283 ();
 FILLCELL_X1 PHY_6284 ();
 FILLCELL_X1 PHY_6285 ();
 FILLCELL_X1 PHY_6286 ();
 FILLCELL_X1 PHY_6287 ();
 FILLCELL_X1 PHY_6288 ();
 FILLCELL_X1 PHY_6289 ();
 FILLCELL_X1 PHY_629 ();
 FILLCELL_X1 PHY_6290 ();
 FILLCELL_X1 PHY_6291 ();
 FILLCELL_X1 PHY_6292 ();
 FILLCELL_X1 PHY_6293 ();
 FILLCELL_X1 PHY_6294 ();
 FILLCELL_X1 PHY_6295 ();
 FILLCELL_X1 PHY_6296 ();
 FILLCELL_X1 PHY_6297 ();
 FILLCELL_X1 PHY_6298 ();
 FILLCELL_X1 PHY_6299 ();
 FILLCELL_X1 PHY_63 ();
 FILLCELL_X1 PHY_630 ();
 FILLCELL_X1 PHY_6300 ();
 FILLCELL_X1 PHY_6301 ();
 FILLCELL_X1 PHY_6302 ();
 FILLCELL_X1 PHY_6303 ();
 FILLCELL_X1 PHY_6304 ();
 FILLCELL_X1 PHY_6305 ();
 FILLCELL_X1 PHY_6306 ();
 FILLCELL_X1 PHY_6307 ();
 FILLCELL_X1 PHY_6308 ();
 FILLCELL_X1 PHY_6309 ();
 FILLCELL_X1 PHY_631 ();
 FILLCELL_X1 PHY_6310 ();
 FILLCELL_X1 PHY_6311 ();
 FILLCELL_X1 PHY_6312 ();
 FILLCELL_X1 PHY_6313 ();
 FILLCELL_X1 PHY_6314 ();
 FILLCELL_X1 PHY_6315 ();
 FILLCELL_X1 PHY_6316 ();
 FILLCELL_X1 PHY_6317 ();
 FILLCELL_X1 PHY_6318 ();
 FILLCELL_X1 PHY_6319 ();
 FILLCELL_X1 PHY_632 ();
 FILLCELL_X1 PHY_6320 ();
 FILLCELL_X1 PHY_6321 ();
 FILLCELL_X1 PHY_6322 ();
 FILLCELL_X1 PHY_6323 ();
 FILLCELL_X1 PHY_6324 ();
 FILLCELL_X1 PHY_6325 ();
 FILLCELL_X1 PHY_6326 ();
 FILLCELL_X1 PHY_6327 ();
 FILLCELL_X1 PHY_6328 ();
 FILLCELL_X1 PHY_6329 ();
 FILLCELL_X1 PHY_633 ();
 FILLCELL_X1 PHY_6330 ();
 FILLCELL_X1 PHY_6331 ();
 FILLCELL_X1 PHY_6332 ();
 FILLCELL_X1 PHY_6333 ();
 FILLCELL_X1 PHY_6334 ();
 FILLCELL_X1 PHY_6335 ();
 FILLCELL_X1 PHY_6336 ();
 FILLCELL_X1 PHY_6337 ();
 FILLCELL_X1 PHY_6338 ();
 FILLCELL_X1 PHY_6339 ();
 FILLCELL_X1 PHY_634 ();
 FILLCELL_X1 PHY_6340 ();
 FILLCELL_X1 PHY_6341 ();
 FILLCELL_X1 PHY_6342 ();
 FILLCELL_X1 PHY_6343 ();
 FILLCELL_X1 PHY_6344 ();
 FILLCELL_X1 PHY_6345 ();
 FILLCELL_X1 PHY_6346 ();
 FILLCELL_X1 PHY_6347 ();
 FILLCELL_X1 PHY_6348 ();
 FILLCELL_X1 PHY_6349 ();
 FILLCELL_X1 PHY_635 ();
 FILLCELL_X1 PHY_6350 ();
 FILLCELL_X1 PHY_6351 ();
 FILLCELL_X1 PHY_6352 ();
 FILLCELL_X1 PHY_6353 ();
 FILLCELL_X1 PHY_6354 ();
 FILLCELL_X1 PHY_6355 ();
 FILLCELL_X1 PHY_6356 ();
 FILLCELL_X1 PHY_6357 ();
 FILLCELL_X1 PHY_6358 ();
 FILLCELL_X1 PHY_6359 ();
 FILLCELL_X1 PHY_636 ();
 FILLCELL_X1 PHY_6360 ();
 FILLCELL_X1 PHY_6361 ();
 FILLCELL_X1 PHY_6362 ();
 FILLCELL_X1 PHY_6363 ();
 FILLCELL_X1 PHY_6364 ();
 FILLCELL_X1 PHY_6365 ();
 FILLCELL_X1 PHY_6366 ();
 FILLCELL_X1 PHY_6367 ();
 FILLCELL_X1 PHY_6368 ();
 FILLCELL_X1 PHY_6369 ();
 FILLCELL_X1 PHY_637 ();
 FILLCELL_X1 PHY_6370 ();
 FILLCELL_X1 PHY_6371 ();
 FILLCELL_X1 PHY_6372 ();
 FILLCELL_X1 PHY_6373 ();
 FILLCELL_X1 PHY_6374 ();
 FILLCELL_X1 PHY_6375 ();
 FILLCELL_X1 PHY_6376 ();
 FILLCELL_X1 PHY_6377 ();
 FILLCELL_X1 PHY_6378 ();
 FILLCELL_X1 PHY_6379 ();
 FILLCELL_X1 PHY_638 ();
 FILLCELL_X1 PHY_6380 ();
 FILLCELL_X1 PHY_6381 ();
 FILLCELL_X1 PHY_6382 ();
 FILLCELL_X1 PHY_6383 ();
 FILLCELL_X1 PHY_6384 ();
 FILLCELL_X1 PHY_6385 ();
 FILLCELL_X1 PHY_6386 ();
 FILLCELL_X1 PHY_6387 ();
 FILLCELL_X1 PHY_6388 ();
 FILLCELL_X1 PHY_6389 ();
 FILLCELL_X1 PHY_639 ();
 FILLCELL_X1 PHY_6390 ();
 FILLCELL_X1 PHY_6391 ();
 FILLCELL_X1 PHY_6392 ();
 FILLCELL_X1 PHY_6393 ();
 FILLCELL_X1 PHY_6394 ();
 FILLCELL_X1 PHY_6395 ();
 FILLCELL_X1 PHY_6396 ();
 FILLCELL_X1 PHY_6397 ();
 FILLCELL_X1 PHY_6398 ();
 FILLCELL_X1 PHY_6399 ();
 FILLCELL_X1 PHY_64 ();
 FILLCELL_X1 PHY_640 ();
 FILLCELL_X1 PHY_6400 ();
 FILLCELL_X1 PHY_6401 ();
 FILLCELL_X1 PHY_6402 ();
 FILLCELL_X1 PHY_6403 ();
 FILLCELL_X1 PHY_6404 ();
 FILLCELL_X1 PHY_6405 ();
 FILLCELL_X1 PHY_6406 ();
 FILLCELL_X1 PHY_6407 ();
 FILLCELL_X1 PHY_6408 ();
 FILLCELL_X1 PHY_6409 ();
 FILLCELL_X1 PHY_641 ();
 FILLCELL_X1 PHY_6410 ();
 FILLCELL_X1 PHY_6411 ();
 FILLCELL_X1 PHY_6412 ();
 FILLCELL_X1 PHY_6413 ();
 FILLCELL_X1 PHY_6414 ();
 FILLCELL_X1 PHY_6415 ();
 FILLCELL_X1 PHY_6416 ();
 FILLCELL_X1 PHY_6417 ();
 FILLCELL_X1 PHY_6418 ();
 FILLCELL_X1 PHY_6419 ();
 FILLCELL_X1 PHY_642 ();
 FILLCELL_X1 PHY_6420 ();
 FILLCELL_X1 PHY_6421 ();
 FILLCELL_X1 PHY_6422 ();
 FILLCELL_X1 PHY_6423 ();
 FILLCELL_X1 PHY_6424 ();
 FILLCELL_X1 PHY_6425 ();
 FILLCELL_X1 PHY_6426 ();
 FILLCELL_X1 PHY_6427 ();
 FILLCELL_X1 PHY_6428 ();
 FILLCELL_X1 PHY_6429 ();
 FILLCELL_X1 PHY_643 ();
 FILLCELL_X1 PHY_6430 ();
 FILLCELL_X1 PHY_6431 ();
 FILLCELL_X1 PHY_6432 ();
 FILLCELL_X1 PHY_6433 ();
 FILLCELL_X1 PHY_6434 ();
 FILLCELL_X1 PHY_6435 ();
 FILLCELL_X1 PHY_6436 ();
 FILLCELL_X1 PHY_6437 ();
 FILLCELL_X1 PHY_6438 ();
 FILLCELL_X1 PHY_6439 ();
 FILLCELL_X1 PHY_644 ();
 FILLCELL_X1 PHY_6440 ();
 FILLCELL_X1 PHY_6441 ();
 FILLCELL_X1 PHY_6442 ();
 FILLCELL_X1 PHY_6443 ();
 FILLCELL_X1 PHY_6444 ();
 FILLCELL_X1 PHY_6445 ();
 FILLCELL_X1 PHY_6446 ();
 FILLCELL_X1 PHY_6447 ();
 FILLCELL_X1 PHY_6448 ();
 FILLCELL_X1 PHY_6449 ();
 FILLCELL_X1 PHY_645 ();
 FILLCELL_X1 PHY_6450 ();
 FILLCELL_X1 PHY_6451 ();
 FILLCELL_X1 PHY_6452 ();
 FILLCELL_X1 PHY_6453 ();
 FILLCELL_X1 PHY_6454 ();
 FILLCELL_X1 PHY_6455 ();
 FILLCELL_X1 PHY_6456 ();
 FILLCELL_X1 PHY_6457 ();
 FILLCELL_X1 PHY_6458 ();
 FILLCELL_X1 PHY_6459 ();
 FILLCELL_X1 PHY_646 ();
 FILLCELL_X1 PHY_6460 ();
 FILLCELL_X1 PHY_6461 ();
 FILLCELL_X1 PHY_6462 ();
 FILLCELL_X1 PHY_6463 ();
 FILLCELL_X1 PHY_6464 ();
 FILLCELL_X1 PHY_6465 ();
 FILLCELL_X1 PHY_6466 ();
 FILLCELL_X1 PHY_6467 ();
 FILLCELL_X1 PHY_6468 ();
 FILLCELL_X1 PHY_6469 ();
 FILLCELL_X1 PHY_647 ();
 FILLCELL_X1 PHY_6470 ();
 FILLCELL_X1 PHY_6471 ();
 FILLCELL_X1 PHY_6472 ();
 FILLCELL_X1 PHY_6473 ();
 FILLCELL_X1 PHY_6474 ();
 FILLCELL_X1 PHY_6475 ();
 FILLCELL_X1 PHY_6476 ();
 FILLCELL_X1 PHY_6477 ();
 FILLCELL_X1 PHY_6478 ();
 FILLCELL_X1 PHY_6479 ();
 FILLCELL_X1 PHY_648 ();
 FILLCELL_X1 PHY_6480 ();
 FILLCELL_X1 PHY_6481 ();
 FILLCELL_X1 PHY_6482 ();
 FILLCELL_X1 PHY_6483 ();
 FILLCELL_X1 PHY_6484 ();
 FILLCELL_X1 PHY_6485 ();
 FILLCELL_X1 PHY_6486 ();
 FILLCELL_X1 PHY_6487 ();
 FILLCELL_X1 PHY_6488 ();
 FILLCELL_X1 PHY_6489 ();
 FILLCELL_X1 PHY_649 ();
 FILLCELL_X1 PHY_6490 ();
 FILLCELL_X1 PHY_6491 ();
 FILLCELL_X1 PHY_6492 ();
 FILLCELL_X1 PHY_6493 ();
 FILLCELL_X1 PHY_6494 ();
 FILLCELL_X1 PHY_6495 ();
 FILLCELL_X1 PHY_6496 ();
 FILLCELL_X1 PHY_6497 ();
 FILLCELL_X1 PHY_6498 ();
 FILLCELL_X1 PHY_6499 ();
 FILLCELL_X1 PHY_65 ();
 FILLCELL_X1 PHY_650 ();
 FILLCELL_X1 PHY_6500 ();
 FILLCELL_X1 PHY_6501 ();
 FILLCELL_X1 PHY_6502 ();
 FILLCELL_X1 PHY_6503 ();
 FILLCELL_X1 PHY_6504 ();
 FILLCELL_X1 PHY_6505 ();
 FILLCELL_X1 PHY_6506 ();
 FILLCELL_X1 PHY_6507 ();
 FILLCELL_X1 PHY_6508 ();
 FILLCELL_X1 PHY_6509 ();
 FILLCELL_X1 PHY_651 ();
 FILLCELL_X1 PHY_6510 ();
 FILLCELL_X1 PHY_6511 ();
 FILLCELL_X1 PHY_6512 ();
 FILLCELL_X1 PHY_6513 ();
 FILLCELL_X1 PHY_6514 ();
 FILLCELL_X1 PHY_6515 ();
 FILLCELL_X1 PHY_6516 ();
 FILLCELL_X1 PHY_6517 ();
 FILLCELL_X1 PHY_6518 ();
 FILLCELL_X1 PHY_6519 ();
 FILLCELL_X1 PHY_652 ();
 FILLCELL_X1 PHY_6520 ();
 FILLCELL_X1 PHY_6521 ();
 FILLCELL_X1 PHY_6522 ();
 FILLCELL_X1 PHY_6523 ();
 FILLCELL_X1 PHY_6524 ();
 FILLCELL_X1 PHY_6525 ();
 FILLCELL_X1 PHY_6526 ();
 FILLCELL_X1 PHY_6527 ();
 FILLCELL_X1 PHY_6528 ();
 FILLCELL_X1 PHY_6529 ();
 FILLCELL_X1 PHY_653 ();
 FILLCELL_X1 PHY_6530 ();
 FILLCELL_X1 PHY_6531 ();
 FILLCELL_X1 PHY_6532 ();
 FILLCELL_X1 PHY_6533 ();
 FILLCELL_X1 PHY_6534 ();
 FILLCELL_X1 PHY_6535 ();
 FILLCELL_X1 PHY_6536 ();
 FILLCELL_X1 PHY_6537 ();
 FILLCELL_X1 PHY_6538 ();
 FILLCELL_X1 PHY_6539 ();
 FILLCELL_X1 PHY_654 ();
 FILLCELL_X1 PHY_6540 ();
 FILLCELL_X1 PHY_6541 ();
 FILLCELL_X1 PHY_6542 ();
 FILLCELL_X1 PHY_6543 ();
 FILLCELL_X1 PHY_6544 ();
 FILLCELL_X1 PHY_6545 ();
 FILLCELL_X1 PHY_6546 ();
 FILLCELL_X1 PHY_6547 ();
 FILLCELL_X1 PHY_6548 ();
 FILLCELL_X1 PHY_6549 ();
 FILLCELL_X1 PHY_655 ();
 FILLCELL_X1 PHY_6550 ();
 FILLCELL_X1 PHY_6551 ();
 FILLCELL_X1 PHY_6552 ();
 FILLCELL_X1 PHY_6553 ();
 FILLCELL_X1 PHY_6554 ();
 FILLCELL_X1 PHY_6555 ();
 FILLCELL_X1 PHY_6556 ();
 FILLCELL_X1 PHY_6557 ();
 FILLCELL_X1 PHY_6558 ();
 FILLCELL_X1 PHY_6559 ();
 FILLCELL_X1 PHY_656 ();
 FILLCELL_X1 PHY_6560 ();
 FILLCELL_X1 PHY_6561 ();
 FILLCELL_X1 PHY_6562 ();
 FILLCELL_X1 PHY_6563 ();
 FILLCELL_X1 PHY_6564 ();
 FILLCELL_X1 PHY_6565 ();
 FILLCELL_X1 PHY_6566 ();
 FILLCELL_X1 PHY_6567 ();
 FILLCELL_X1 PHY_6568 ();
 FILLCELL_X1 PHY_6569 ();
 FILLCELL_X1 PHY_657 ();
 FILLCELL_X1 PHY_6570 ();
 FILLCELL_X1 PHY_6571 ();
 FILLCELL_X1 PHY_6572 ();
 FILLCELL_X1 PHY_6573 ();
 FILLCELL_X1 PHY_6574 ();
 FILLCELL_X1 PHY_6575 ();
 FILLCELL_X1 PHY_6576 ();
 FILLCELL_X1 PHY_6577 ();
 FILLCELL_X1 PHY_6578 ();
 FILLCELL_X1 PHY_6579 ();
 FILLCELL_X1 PHY_658 ();
 FILLCELL_X1 PHY_6580 ();
 FILLCELL_X1 PHY_6581 ();
 FILLCELL_X1 PHY_6582 ();
 FILLCELL_X1 PHY_6583 ();
 FILLCELL_X1 PHY_6584 ();
 FILLCELL_X1 PHY_6585 ();
 FILLCELL_X1 PHY_6586 ();
 FILLCELL_X1 PHY_6587 ();
 FILLCELL_X1 PHY_6588 ();
 FILLCELL_X1 PHY_6589 ();
 FILLCELL_X1 PHY_659 ();
 FILLCELL_X1 PHY_6590 ();
 FILLCELL_X1 PHY_6591 ();
 FILLCELL_X1 PHY_6592 ();
 FILLCELL_X1 PHY_6593 ();
 FILLCELL_X1 PHY_6594 ();
 FILLCELL_X1 PHY_6595 ();
 FILLCELL_X1 PHY_6596 ();
 FILLCELL_X1 PHY_6597 ();
 FILLCELL_X1 PHY_6598 ();
 FILLCELL_X1 PHY_6599 ();
 FILLCELL_X1 PHY_66 ();
 FILLCELL_X1 PHY_660 ();
 FILLCELL_X1 PHY_6600 ();
 FILLCELL_X1 PHY_6601 ();
 FILLCELL_X1 PHY_6602 ();
 FILLCELL_X1 PHY_6603 ();
 FILLCELL_X1 PHY_6604 ();
 FILLCELL_X1 PHY_6605 ();
 FILLCELL_X1 PHY_6606 ();
 FILLCELL_X1 PHY_6607 ();
 FILLCELL_X1 PHY_6608 ();
 FILLCELL_X1 PHY_6609 ();
 FILLCELL_X1 PHY_661 ();
 FILLCELL_X1 PHY_6610 ();
 FILLCELL_X1 PHY_6611 ();
 FILLCELL_X1 PHY_6612 ();
 FILLCELL_X1 PHY_6613 ();
 FILLCELL_X1 PHY_6614 ();
 FILLCELL_X1 PHY_6615 ();
 FILLCELL_X1 PHY_6616 ();
 FILLCELL_X1 PHY_6617 ();
 FILLCELL_X1 PHY_6618 ();
 FILLCELL_X1 PHY_6619 ();
 FILLCELL_X1 PHY_662 ();
 FILLCELL_X1 PHY_6620 ();
 FILLCELL_X1 PHY_6621 ();
 FILLCELL_X1 PHY_6622 ();
 FILLCELL_X1 PHY_6623 ();
 FILLCELL_X1 PHY_6624 ();
 FILLCELL_X1 PHY_6625 ();
 FILLCELL_X1 PHY_6626 ();
 FILLCELL_X1 PHY_6627 ();
 FILLCELL_X1 PHY_6628 ();
 FILLCELL_X1 PHY_6629 ();
 FILLCELL_X1 PHY_663 ();
 FILLCELL_X1 PHY_6630 ();
 FILLCELL_X1 PHY_6631 ();
 FILLCELL_X1 PHY_6632 ();
 FILLCELL_X1 PHY_6633 ();
 FILLCELL_X1 PHY_6634 ();
 FILLCELL_X1 PHY_6635 ();
 FILLCELL_X1 PHY_6636 ();
 FILLCELL_X1 PHY_6637 ();
 FILLCELL_X1 PHY_6638 ();
 FILLCELL_X1 PHY_6639 ();
 FILLCELL_X1 PHY_664 ();
 FILLCELL_X1 PHY_6640 ();
 FILLCELL_X1 PHY_6641 ();
 FILLCELL_X1 PHY_6642 ();
 FILLCELL_X1 PHY_6643 ();
 FILLCELL_X1 PHY_6644 ();
 FILLCELL_X1 PHY_6645 ();
 FILLCELL_X1 PHY_6646 ();
 FILLCELL_X1 PHY_6647 ();
 FILLCELL_X1 PHY_6648 ();
 FILLCELL_X1 PHY_6649 ();
 FILLCELL_X1 PHY_665 ();
 FILLCELL_X1 PHY_6650 ();
 FILLCELL_X1 PHY_6651 ();
 FILLCELL_X1 PHY_6652 ();
 FILLCELL_X1 PHY_6653 ();
 FILLCELL_X1 PHY_6654 ();
 FILLCELL_X1 PHY_6655 ();
 FILLCELL_X1 PHY_6656 ();
 FILLCELL_X1 PHY_6657 ();
 FILLCELL_X1 PHY_6658 ();
 FILLCELL_X1 PHY_6659 ();
 FILLCELL_X1 PHY_666 ();
 FILLCELL_X1 PHY_6660 ();
 FILLCELL_X1 PHY_6661 ();
 FILLCELL_X1 PHY_6662 ();
 FILLCELL_X1 PHY_6663 ();
 FILLCELL_X1 PHY_6664 ();
 FILLCELL_X1 PHY_6665 ();
 FILLCELL_X1 PHY_6666 ();
 FILLCELL_X1 PHY_6667 ();
 FILLCELL_X1 PHY_6668 ();
 FILLCELL_X1 PHY_6669 ();
 FILLCELL_X1 PHY_667 ();
 FILLCELL_X1 PHY_6670 ();
 FILLCELL_X1 PHY_6671 ();
 FILLCELL_X1 PHY_6672 ();
 FILLCELL_X1 PHY_6673 ();
 FILLCELL_X1 PHY_6674 ();
 FILLCELL_X1 PHY_6675 ();
 FILLCELL_X1 PHY_6676 ();
 FILLCELL_X1 PHY_6677 ();
 FILLCELL_X1 PHY_6678 ();
 FILLCELL_X1 PHY_6679 ();
 FILLCELL_X1 PHY_668 ();
 FILLCELL_X1 PHY_6680 ();
 FILLCELL_X1 PHY_6681 ();
 FILLCELL_X1 PHY_6682 ();
 FILLCELL_X1 PHY_6683 ();
 FILLCELL_X1 PHY_6684 ();
 FILLCELL_X1 PHY_6685 ();
 FILLCELL_X1 PHY_6686 ();
 FILLCELL_X1 PHY_6687 ();
 FILLCELL_X1 PHY_6688 ();
 FILLCELL_X1 PHY_6689 ();
 FILLCELL_X1 PHY_669 ();
 FILLCELL_X1 PHY_6690 ();
 FILLCELL_X1 PHY_6691 ();
 FILLCELL_X1 PHY_6692 ();
 FILLCELL_X1 PHY_6693 ();
 FILLCELL_X1 PHY_6694 ();
 FILLCELL_X1 PHY_6695 ();
 FILLCELL_X1 PHY_6696 ();
 FILLCELL_X1 PHY_6697 ();
 FILLCELL_X1 PHY_6698 ();
 FILLCELL_X1 PHY_6699 ();
 FILLCELL_X1 PHY_67 ();
 FILLCELL_X1 PHY_670 ();
 FILLCELL_X1 PHY_6700 ();
 FILLCELL_X1 PHY_6701 ();
 FILLCELL_X1 PHY_6702 ();
 FILLCELL_X1 PHY_6703 ();
 FILLCELL_X1 PHY_6704 ();
 FILLCELL_X1 PHY_6705 ();
 FILLCELL_X1 PHY_6706 ();
 FILLCELL_X1 PHY_6707 ();
 FILLCELL_X1 PHY_6708 ();
 FILLCELL_X1 PHY_6709 ();
 FILLCELL_X1 PHY_671 ();
 FILLCELL_X1 PHY_6710 ();
 FILLCELL_X1 PHY_6711 ();
 FILLCELL_X1 PHY_6712 ();
 FILLCELL_X1 PHY_6713 ();
 FILLCELL_X1 PHY_6714 ();
 FILLCELL_X1 PHY_6715 ();
 FILLCELL_X1 PHY_6716 ();
 FILLCELL_X1 PHY_6717 ();
 FILLCELL_X1 PHY_6718 ();
 FILLCELL_X1 PHY_6719 ();
 FILLCELL_X1 PHY_672 ();
 FILLCELL_X1 PHY_6720 ();
 FILLCELL_X1 PHY_6721 ();
 FILLCELL_X1 PHY_6722 ();
 FILLCELL_X1 PHY_6723 ();
 FILLCELL_X1 PHY_6724 ();
 FILLCELL_X1 PHY_6725 ();
 FILLCELL_X1 PHY_6726 ();
 FILLCELL_X1 PHY_6727 ();
 FILLCELL_X1 PHY_6728 ();
 FILLCELL_X1 PHY_6729 ();
 FILLCELL_X1 PHY_673 ();
 FILLCELL_X1 PHY_6730 ();
 FILLCELL_X1 PHY_6731 ();
 FILLCELL_X1 PHY_6732 ();
 FILLCELL_X1 PHY_6733 ();
 FILLCELL_X1 PHY_6734 ();
 FILLCELL_X1 PHY_6735 ();
 FILLCELL_X1 PHY_6736 ();
 FILLCELL_X1 PHY_6737 ();
 FILLCELL_X1 PHY_6738 ();
 FILLCELL_X1 PHY_6739 ();
 FILLCELL_X1 PHY_674 ();
 FILLCELL_X1 PHY_6740 ();
 FILLCELL_X1 PHY_6741 ();
 FILLCELL_X1 PHY_6742 ();
 FILLCELL_X1 PHY_6743 ();
 FILLCELL_X1 PHY_6744 ();
 FILLCELL_X1 PHY_6745 ();
 FILLCELL_X1 PHY_6746 ();
 FILLCELL_X1 PHY_6747 ();
 FILLCELL_X1 PHY_6748 ();
 FILLCELL_X1 PHY_6749 ();
 FILLCELL_X1 PHY_675 ();
 FILLCELL_X1 PHY_6750 ();
 FILLCELL_X1 PHY_6751 ();
 FILLCELL_X1 PHY_6752 ();
 FILLCELL_X1 PHY_6753 ();
 FILLCELL_X1 PHY_6754 ();
 FILLCELL_X1 PHY_6755 ();
 FILLCELL_X1 PHY_6756 ();
 FILLCELL_X1 PHY_6757 ();
 FILLCELL_X1 PHY_6758 ();
 FILLCELL_X1 PHY_6759 ();
 FILLCELL_X1 PHY_676 ();
 FILLCELL_X1 PHY_6760 ();
 FILLCELL_X1 PHY_6761 ();
 FILLCELL_X1 PHY_6762 ();
 FILLCELL_X1 PHY_6763 ();
 FILLCELL_X1 PHY_6764 ();
 FILLCELL_X1 PHY_6765 ();
 FILLCELL_X1 PHY_6766 ();
 FILLCELL_X1 PHY_6767 ();
 FILLCELL_X1 PHY_6768 ();
 FILLCELL_X1 PHY_6769 ();
 FILLCELL_X1 PHY_677 ();
 FILLCELL_X1 PHY_6770 ();
 FILLCELL_X1 PHY_6771 ();
 FILLCELL_X1 PHY_6772 ();
 FILLCELL_X1 PHY_6773 ();
 FILLCELL_X1 PHY_6774 ();
 FILLCELL_X1 PHY_6775 ();
 FILLCELL_X1 PHY_6776 ();
 FILLCELL_X1 PHY_6777 ();
 FILLCELL_X1 PHY_6778 ();
 FILLCELL_X1 PHY_6779 ();
 FILLCELL_X1 PHY_678 ();
 FILLCELL_X1 PHY_6780 ();
 FILLCELL_X1 PHY_6781 ();
 FILLCELL_X1 PHY_6782 ();
 FILLCELL_X1 PHY_6783 ();
 FILLCELL_X1 PHY_6784 ();
 FILLCELL_X1 PHY_6785 ();
 FILLCELL_X1 PHY_6786 ();
 FILLCELL_X1 PHY_6787 ();
 FILLCELL_X1 PHY_6788 ();
 FILLCELL_X1 PHY_6789 ();
 FILLCELL_X1 PHY_679 ();
 FILLCELL_X1 PHY_6790 ();
 FILLCELL_X1 PHY_6791 ();
 FILLCELL_X1 PHY_6792 ();
 FILLCELL_X1 PHY_6793 ();
 FILLCELL_X1 PHY_6794 ();
 FILLCELL_X1 PHY_6795 ();
 FILLCELL_X1 PHY_6796 ();
 FILLCELL_X1 PHY_6797 ();
 FILLCELL_X1 PHY_6798 ();
 FILLCELL_X1 PHY_6799 ();
 FILLCELL_X1 PHY_68 ();
 FILLCELL_X1 PHY_680 ();
 FILLCELL_X1 PHY_6800 ();
 FILLCELL_X1 PHY_6801 ();
 FILLCELL_X1 PHY_6802 ();
 FILLCELL_X1 PHY_6803 ();
 FILLCELL_X1 PHY_6804 ();
 FILLCELL_X1 PHY_6805 ();
 FILLCELL_X1 PHY_6806 ();
 FILLCELL_X1 PHY_6807 ();
 FILLCELL_X1 PHY_6808 ();
 FILLCELL_X1 PHY_6809 ();
 FILLCELL_X1 PHY_681 ();
 FILLCELL_X1 PHY_6810 ();
 FILLCELL_X1 PHY_6811 ();
 FILLCELL_X1 PHY_6812 ();
 FILLCELL_X1 PHY_6813 ();
 FILLCELL_X1 PHY_6814 ();
 FILLCELL_X1 PHY_6815 ();
 FILLCELL_X1 PHY_6816 ();
 FILLCELL_X1 PHY_6817 ();
 FILLCELL_X1 PHY_6818 ();
 FILLCELL_X1 PHY_6819 ();
 FILLCELL_X1 PHY_682 ();
 FILLCELL_X1 PHY_6820 ();
 FILLCELL_X1 PHY_6821 ();
 FILLCELL_X1 PHY_6822 ();
 FILLCELL_X1 PHY_6823 ();
 FILLCELL_X1 PHY_6824 ();
 FILLCELL_X1 PHY_6825 ();
 FILLCELL_X1 PHY_6826 ();
 FILLCELL_X1 PHY_6827 ();
 FILLCELL_X1 PHY_6828 ();
 FILLCELL_X1 PHY_6829 ();
 FILLCELL_X1 PHY_683 ();
 FILLCELL_X1 PHY_6830 ();
 FILLCELL_X1 PHY_6831 ();
 FILLCELL_X1 PHY_6832 ();
 FILLCELL_X1 PHY_6833 ();
 FILLCELL_X1 PHY_6834 ();
 FILLCELL_X1 PHY_6835 ();
 FILLCELL_X1 PHY_6836 ();
 FILLCELL_X1 PHY_6837 ();
 FILLCELL_X1 PHY_6838 ();
 FILLCELL_X1 PHY_6839 ();
 FILLCELL_X1 PHY_684 ();
 FILLCELL_X1 PHY_6840 ();
 FILLCELL_X1 PHY_6841 ();
 FILLCELL_X1 PHY_6842 ();
 FILLCELL_X1 PHY_6843 ();
 FILLCELL_X1 PHY_6844 ();
 FILLCELL_X1 PHY_6845 ();
 FILLCELL_X1 PHY_6846 ();
 FILLCELL_X1 PHY_6847 ();
 FILLCELL_X1 PHY_6848 ();
 FILLCELL_X1 PHY_6849 ();
 FILLCELL_X1 PHY_685 ();
 FILLCELL_X1 PHY_6850 ();
 FILLCELL_X1 PHY_6851 ();
 FILLCELL_X1 PHY_6852 ();
 FILLCELL_X1 PHY_6853 ();
 FILLCELL_X1 PHY_6854 ();
 FILLCELL_X1 PHY_6855 ();
 FILLCELL_X1 PHY_6856 ();
 FILLCELL_X1 PHY_6857 ();
 FILLCELL_X1 PHY_6858 ();
 FILLCELL_X1 PHY_6859 ();
 FILLCELL_X1 PHY_686 ();
 FILLCELL_X1 PHY_6860 ();
 FILLCELL_X1 PHY_6861 ();
 FILLCELL_X1 PHY_6862 ();
 FILLCELL_X1 PHY_6863 ();
 FILLCELL_X1 PHY_6864 ();
 FILLCELL_X1 PHY_6865 ();
 FILLCELL_X1 PHY_6866 ();
 FILLCELL_X1 PHY_6867 ();
 FILLCELL_X1 PHY_6868 ();
 FILLCELL_X1 PHY_6869 ();
 FILLCELL_X1 PHY_687 ();
 FILLCELL_X1 PHY_6870 ();
 FILLCELL_X1 PHY_6871 ();
 FILLCELL_X1 PHY_6872 ();
 FILLCELL_X1 PHY_6873 ();
 FILLCELL_X1 PHY_6874 ();
 FILLCELL_X1 PHY_6875 ();
 FILLCELL_X1 PHY_6876 ();
 FILLCELL_X1 PHY_6877 ();
 FILLCELL_X1 PHY_6878 ();
 FILLCELL_X1 PHY_6879 ();
 FILLCELL_X1 PHY_688 ();
 FILLCELL_X1 PHY_6880 ();
 FILLCELL_X1 PHY_6881 ();
 FILLCELL_X1 PHY_6882 ();
 FILLCELL_X1 PHY_6883 ();
 FILLCELL_X1 PHY_6884 ();
 FILLCELL_X1 PHY_6885 ();
 FILLCELL_X1 PHY_6886 ();
 FILLCELL_X1 PHY_6887 ();
 FILLCELL_X1 PHY_6888 ();
 FILLCELL_X1 PHY_6889 ();
 FILLCELL_X1 PHY_689 ();
 FILLCELL_X1 PHY_6890 ();
 FILLCELL_X1 PHY_6891 ();
 FILLCELL_X1 PHY_6892 ();
 FILLCELL_X1 PHY_6893 ();
 FILLCELL_X1 PHY_6894 ();
 FILLCELL_X1 PHY_6895 ();
 FILLCELL_X1 PHY_6896 ();
 FILLCELL_X1 PHY_6897 ();
 FILLCELL_X1 PHY_6898 ();
 FILLCELL_X1 PHY_6899 ();
 FILLCELL_X1 PHY_69 ();
 FILLCELL_X1 PHY_690 ();
 FILLCELL_X1 PHY_6900 ();
 FILLCELL_X1 PHY_6901 ();
 FILLCELL_X1 PHY_6902 ();
 FILLCELL_X1 PHY_6903 ();
 FILLCELL_X1 PHY_6904 ();
 FILLCELL_X1 PHY_6905 ();
 FILLCELL_X1 PHY_6906 ();
 FILLCELL_X1 PHY_6907 ();
 FILLCELL_X1 PHY_6908 ();
 FILLCELL_X1 PHY_6909 ();
 FILLCELL_X1 PHY_691 ();
 FILLCELL_X1 PHY_6910 ();
 FILLCELL_X1 PHY_6911 ();
 FILLCELL_X1 PHY_6912 ();
 FILLCELL_X1 PHY_6913 ();
 FILLCELL_X1 PHY_6914 ();
 FILLCELL_X1 PHY_6915 ();
 FILLCELL_X1 PHY_6916 ();
 FILLCELL_X1 PHY_6917 ();
 FILLCELL_X1 PHY_6918 ();
 FILLCELL_X1 PHY_6919 ();
 FILLCELL_X1 PHY_692 ();
 FILLCELL_X1 PHY_6920 ();
 FILLCELL_X1 PHY_6921 ();
 FILLCELL_X1 PHY_6922 ();
 FILLCELL_X1 PHY_6923 ();
 FILLCELL_X1 PHY_6924 ();
 FILLCELL_X1 PHY_6925 ();
 FILLCELL_X1 PHY_6926 ();
 FILLCELL_X1 PHY_6927 ();
 FILLCELL_X1 PHY_6928 ();
 FILLCELL_X1 PHY_6929 ();
 FILLCELL_X1 PHY_693 ();
 FILLCELL_X1 PHY_6930 ();
 FILLCELL_X1 PHY_6931 ();
 FILLCELL_X1 PHY_6932 ();
 FILLCELL_X1 PHY_6933 ();
 FILLCELL_X1 PHY_6934 ();
 FILLCELL_X1 PHY_6935 ();
 FILLCELL_X1 PHY_6936 ();
 FILLCELL_X1 PHY_6937 ();
 FILLCELL_X1 PHY_6938 ();
 FILLCELL_X1 PHY_6939 ();
 FILLCELL_X1 PHY_694 ();
 FILLCELL_X1 PHY_6940 ();
 FILLCELL_X1 PHY_6941 ();
 FILLCELL_X1 PHY_6942 ();
 FILLCELL_X1 PHY_6943 ();
 FILLCELL_X1 PHY_6944 ();
 FILLCELL_X1 PHY_6945 ();
 FILLCELL_X1 PHY_6946 ();
 FILLCELL_X1 PHY_6947 ();
 FILLCELL_X1 PHY_6948 ();
 FILLCELL_X1 PHY_6949 ();
 FILLCELL_X1 PHY_695 ();
 FILLCELL_X1 PHY_6950 ();
 FILLCELL_X1 PHY_6951 ();
 FILLCELL_X1 PHY_6952 ();
 FILLCELL_X1 PHY_6953 ();
 FILLCELL_X1 PHY_6954 ();
 FILLCELL_X1 PHY_6955 ();
 FILLCELL_X1 PHY_6956 ();
 FILLCELL_X1 PHY_6957 ();
 FILLCELL_X1 PHY_6958 ();
 FILLCELL_X1 PHY_6959 ();
 FILLCELL_X1 PHY_696 ();
 FILLCELL_X1 PHY_6960 ();
 FILLCELL_X1 PHY_6961 ();
 FILLCELL_X1 PHY_6962 ();
 FILLCELL_X1 PHY_6963 ();
 FILLCELL_X1 PHY_6964 ();
 FILLCELL_X1 PHY_6965 ();
 FILLCELL_X1 PHY_6966 ();
 FILLCELL_X1 PHY_6967 ();
 FILLCELL_X1 PHY_6968 ();
 FILLCELL_X1 PHY_6969 ();
 FILLCELL_X1 PHY_697 ();
 FILLCELL_X1 PHY_6970 ();
 FILLCELL_X1 PHY_6971 ();
 FILLCELL_X1 PHY_6972 ();
 FILLCELL_X1 PHY_6973 ();
 FILLCELL_X1 PHY_6974 ();
 FILLCELL_X1 PHY_6975 ();
 FILLCELL_X1 PHY_6976 ();
 FILLCELL_X1 PHY_6977 ();
 FILLCELL_X1 PHY_6978 ();
 FILLCELL_X1 PHY_6979 ();
 FILLCELL_X1 PHY_698 ();
 FILLCELL_X1 PHY_6980 ();
 FILLCELL_X1 PHY_6981 ();
 FILLCELL_X1 PHY_6982 ();
 FILLCELL_X1 PHY_6983 ();
 FILLCELL_X1 PHY_6984 ();
 FILLCELL_X1 PHY_6985 ();
 FILLCELL_X1 PHY_6986 ();
 FILLCELL_X1 PHY_6987 ();
 FILLCELL_X1 PHY_6988 ();
 FILLCELL_X1 PHY_6989 ();
 FILLCELL_X1 PHY_699 ();
 FILLCELL_X1 PHY_6990 ();
 FILLCELL_X1 PHY_6991 ();
 FILLCELL_X1 PHY_6992 ();
 FILLCELL_X1 PHY_6993 ();
 FILLCELL_X1 PHY_6994 ();
 FILLCELL_X1 PHY_6995 ();
 FILLCELL_X1 PHY_6996 ();
 FILLCELL_X1 PHY_6997 ();
 FILLCELL_X1 PHY_6998 ();
 FILLCELL_X1 PHY_6999 ();
 FILLCELL_X1 PHY_7 ();
 FILLCELL_X1 PHY_70 ();
 FILLCELL_X1 PHY_700 ();
 FILLCELL_X1 PHY_7000 ();
 FILLCELL_X1 PHY_7001 ();
 FILLCELL_X1 PHY_7002 ();
 FILLCELL_X1 PHY_7003 ();
 FILLCELL_X1 PHY_7004 ();
 FILLCELL_X1 PHY_7005 ();
 FILLCELL_X1 PHY_7006 ();
 FILLCELL_X1 PHY_7007 ();
 FILLCELL_X1 PHY_7008 ();
 FILLCELL_X1 PHY_7009 ();
 FILLCELL_X1 PHY_701 ();
 FILLCELL_X1 PHY_7010 ();
 FILLCELL_X1 PHY_7011 ();
 FILLCELL_X1 PHY_7012 ();
 FILLCELL_X1 PHY_7013 ();
 FILLCELL_X1 PHY_7014 ();
 FILLCELL_X1 PHY_7015 ();
 FILLCELL_X1 PHY_7016 ();
 FILLCELL_X1 PHY_7017 ();
 FILLCELL_X1 PHY_7018 ();
 FILLCELL_X1 PHY_7019 ();
 FILLCELL_X1 PHY_702 ();
 FILLCELL_X1 PHY_7020 ();
 FILLCELL_X1 PHY_7021 ();
 FILLCELL_X1 PHY_7022 ();
 FILLCELL_X1 PHY_7023 ();
 FILLCELL_X1 PHY_7024 ();
 FILLCELL_X1 PHY_7025 ();
 FILLCELL_X1 PHY_7026 ();
 FILLCELL_X1 PHY_7027 ();
 FILLCELL_X1 PHY_7028 ();
 FILLCELL_X1 PHY_7029 ();
 FILLCELL_X1 PHY_703 ();
 FILLCELL_X1 PHY_7030 ();
 FILLCELL_X1 PHY_7031 ();
 FILLCELL_X1 PHY_7032 ();
 FILLCELL_X1 PHY_7033 ();
 FILLCELL_X1 PHY_7034 ();
 FILLCELL_X1 PHY_7035 ();
 FILLCELL_X1 PHY_7036 ();
 FILLCELL_X1 PHY_7037 ();
 FILLCELL_X1 PHY_7038 ();
 FILLCELL_X1 PHY_7039 ();
 FILLCELL_X1 PHY_704 ();
 FILLCELL_X1 PHY_7040 ();
 FILLCELL_X1 PHY_7041 ();
 FILLCELL_X1 PHY_7042 ();
 FILLCELL_X1 PHY_7043 ();
 FILLCELL_X1 PHY_7044 ();
 FILLCELL_X1 PHY_7045 ();
 FILLCELL_X1 PHY_7046 ();
 FILLCELL_X1 PHY_7047 ();
 FILLCELL_X1 PHY_7048 ();
 FILLCELL_X1 PHY_7049 ();
 FILLCELL_X1 PHY_705 ();
 FILLCELL_X1 PHY_7050 ();
 FILLCELL_X1 PHY_7051 ();
 FILLCELL_X1 PHY_7052 ();
 FILLCELL_X1 PHY_7053 ();
 FILLCELL_X1 PHY_7054 ();
 FILLCELL_X1 PHY_7055 ();
 FILLCELL_X1 PHY_7056 ();
 FILLCELL_X1 PHY_7057 ();
 FILLCELL_X1 PHY_7058 ();
 FILLCELL_X1 PHY_7059 ();
 FILLCELL_X1 PHY_706 ();
 FILLCELL_X1 PHY_7060 ();
 FILLCELL_X1 PHY_7061 ();
 FILLCELL_X1 PHY_7062 ();
 FILLCELL_X1 PHY_7063 ();
 FILLCELL_X1 PHY_7064 ();
 FILLCELL_X1 PHY_7065 ();
 FILLCELL_X1 PHY_7066 ();
 FILLCELL_X1 PHY_7067 ();
 FILLCELL_X1 PHY_7068 ();
 FILLCELL_X1 PHY_7069 ();
 FILLCELL_X1 PHY_707 ();
 FILLCELL_X1 PHY_7070 ();
 FILLCELL_X1 PHY_7071 ();
 FILLCELL_X1 PHY_7072 ();
 FILLCELL_X1 PHY_7073 ();
 FILLCELL_X1 PHY_7074 ();
 FILLCELL_X1 PHY_7075 ();
 FILLCELL_X1 PHY_7076 ();
 FILLCELL_X1 PHY_7077 ();
 FILLCELL_X1 PHY_7078 ();
 FILLCELL_X1 PHY_7079 ();
 FILLCELL_X1 PHY_708 ();
 FILLCELL_X1 PHY_7080 ();
 FILLCELL_X1 PHY_7081 ();
 FILLCELL_X1 PHY_7082 ();
 FILLCELL_X1 PHY_7083 ();
 FILLCELL_X1 PHY_7084 ();
 FILLCELL_X1 PHY_7085 ();
 FILLCELL_X1 PHY_7086 ();
 FILLCELL_X1 PHY_7087 ();
 FILLCELL_X1 PHY_7088 ();
 FILLCELL_X1 PHY_7089 ();
 FILLCELL_X1 PHY_709 ();
 FILLCELL_X1 PHY_7090 ();
 FILLCELL_X1 PHY_7091 ();
 FILLCELL_X1 PHY_7092 ();
 FILLCELL_X1 PHY_7093 ();
 FILLCELL_X1 PHY_7094 ();
 FILLCELL_X1 PHY_7095 ();
 FILLCELL_X1 PHY_7096 ();
 FILLCELL_X1 PHY_7097 ();
 FILLCELL_X1 PHY_7098 ();
 FILLCELL_X1 PHY_7099 ();
 FILLCELL_X1 PHY_71 ();
 FILLCELL_X1 PHY_710 ();
 FILLCELL_X1 PHY_7100 ();
 FILLCELL_X1 PHY_7101 ();
 FILLCELL_X1 PHY_7102 ();
 FILLCELL_X1 PHY_7103 ();
 FILLCELL_X1 PHY_7104 ();
 FILLCELL_X1 PHY_7105 ();
 FILLCELL_X1 PHY_7106 ();
 FILLCELL_X1 PHY_7107 ();
 FILLCELL_X1 PHY_7108 ();
 FILLCELL_X1 PHY_7109 ();
 FILLCELL_X1 PHY_711 ();
 FILLCELL_X1 PHY_7110 ();
 FILLCELL_X1 PHY_7111 ();
 FILLCELL_X1 PHY_7112 ();
 FILLCELL_X1 PHY_7113 ();
 FILLCELL_X1 PHY_7114 ();
 FILLCELL_X1 PHY_7115 ();
 FILLCELL_X1 PHY_7116 ();
 FILLCELL_X1 PHY_7117 ();
 FILLCELL_X1 PHY_7118 ();
 FILLCELL_X1 PHY_7119 ();
 FILLCELL_X1 PHY_712 ();
 FILLCELL_X1 PHY_7120 ();
 FILLCELL_X1 PHY_7121 ();
 FILLCELL_X1 PHY_7122 ();
 FILLCELL_X1 PHY_7123 ();
 FILLCELL_X1 PHY_7124 ();
 FILLCELL_X1 PHY_7125 ();
 FILLCELL_X1 PHY_7126 ();
 FILLCELL_X1 PHY_7127 ();
 FILLCELL_X1 PHY_7128 ();
 FILLCELL_X1 PHY_7129 ();
 FILLCELL_X1 PHY_713 ();
 FILLCELL_X1 PHY_7130 ();
 FILLCELL_X1 PHY_7131 ();
 FILLCELL_X1 PHY_7132 ();
 FILLCELL_X1 PHY_7133 ();
 FILLCELL_X1 PHY_7134 ();
 FILLCELL_X1 PHY_7135 ();
 FILLCELL_X1 PHY_7136 ();
 FILLCELL_X1 PHY_7137 ();
 FILLCELL_X1 PHY_7138 ();
 FILLCELL_X1 PHY_7139 ();
 FILLCELL_X1 PHY_714 ();
 FILLCELL_X1 PHY_7140 ();
 FILLCELL_X1 PHY_7141 ();
 FILLCELL_X1 PHY_7142 ();
 FILLCELL_X1 PHY_7143 ();
 FILLCELL_X1 PHY_7144 ();
 FILLCELL_X1 PHY_7145 ();
 FILLCELL_X1 PHY_7146 ();
 FILLCELL_X1 PHY_7147 ();
 FILLCELL_X1 PHY_7148 ();
 FILLCELL_X1 PHY_7149 ();
 FILLCELL_X1 PHY_715 ();
 FILLCELL_X1 PHY_7150 ();
 FILLCELL_X1 PHY_7151 ();
 FILLCELL_X1 PHY_7152 ();
 FILLCELL_X1 PHY_7153 ();
 FILLCELL_X1 PHY_7154 ();
 FILLCELL_X1 PHY_7155 ();
 FILLCELL_X1 PHY_7156 ();
 FILLCELL_X1 PHY_7157 ();
 FILLCELL_X1 PHY_7158 ();
 FILLCELL_X1 PHY_7159 ();
 FILLCELL_X1 PHY_716 ();
 FILLCELL_X1 PHY_7160 ();
 FILLCELL_X1 PHY_7161 ();
 FILLCELL_X1 PHY_7162 ();
 FILLCELL_X1 PHY_7163 ();
 FILLCELL_X1 PHY_7164 ();
 FILLCELL_X1 PHY_7165 ();
 FILLCELL_X1 PHY_7166 ();
 FILLCELL_X1 PHY_7167 ();
 FILLCELL_X1 PHY_7168 ();
 FILLCELL_X1 PHY_7169 ();
 FILLCELL_X1 PHY_717 ();
 FILLCELL_X1 PHY_7170 ();
 FILLCELL_X1 PHY_7171 ();
 FILLCELL_X1 PHY_7172 ();
 FILLCELL_X1 PHY_7173 ();
 FILLCELL_X1 PHY_7174 ();
 FILLCELL_X1 PHY_7175 ();
 FILLCELL_X1 PHY_7176 ();
 FILLCELL_X1 PHY_7177 ();
 FILLCELL_X1 PHY_7178 ();
 FILLCELL_X1 PHY_7179 ();
 FILLCELL_X1 PHY_718 ();
 FILLCELL_X1 PHY_7180 ();
 FILLCELL_X1 PHY_7181 ();
 FILLCELL_X1 PHY_7182 ();
 FILLCELL_X1 PHY_7183 ();
 FILLCELL_X1 PHY_7184 ();
 FILLCELL_X1 PHY_7185 ();
 FILLCELL_X1 PHY_7186 ();
 FILLCELL_X1 PHY_7187 ();
 FILLCELL_X1 PHY_7188 ();
 FILLCELL_X1 PHY_7189 ();
 FILLCELL_X1 PHY_719 ();
 FILLCELL_X1 PHY_7190 ();
 FILLCELL_X1 PHY_7191 ();
 FILLCELL_X1 PHY_7192 ();
 FILLCELL_X1 PHY_7193 ();
 FILLCELL_X1 PHY_7194 ();
 FILLCELL_X1 PHY_7195 ();
 FILLCELL_X1 PHY_7196 ();
 FILLCELL_X1 PHY_7197 ();
 FILLCELL_X1 PHY_7198 ();
 FILLCELL_X1 PHY_7199 ();
 FILLCELL_X1 PHY_72 ();
 FILLCELL_X1 PHY_720 ();
 FILLCELL_X1 PHY_7200 ();
 FILLCELL_X1 PHY_7201 ();
 FILLCELL_X1 PHY_7202 ();
 FILLCELL_X1 PHY_7203 ();
 FILLCELL_X1 PHY_7204 ();
 FILLCELL_X1 PHY_7205 ();
 FILLCELL_X1 PHY_7206 ();
 FILLCELL_X1 PHY_7207 ();
 FILLCELL_X1 PHY_7208 ();
 FILLCELL_X1 PHY_7209 ();
 FILLCELL_X1 PHY_721 ();
 FILLCELL_X1 PHY_7210 ();
 FILLCELL_X1 PHY_7211 ();
 FILLCELL_X1 PHY_7212 ();
 FILLCELL_X1 PHY_7213 ();
 FILLCELL_X1 PHY_7214 ();
 FILLCELL_X1 PHY_7215 ();
 FILLCELL_X1 PHY_7216 ();
 FILLCELL_X1 PHY_7217 ();
 FILLCELL_X1 PHY_7218 ();
 FILLCELL_X1 PHY_7219 ();
 FILLCELL_X1 PHY_722 ();
 FILLCELL_X1 PHY_7220 ();
 FILLCELL_X1 PHY_7221 ();
 FILLCELL_X1 PHY_7222 ();
 FILLCELL_X1 PHY_7223 ();
 FILLCELL_X1 PHY_7224 ();
 FILLCELL_X1 PHY_7225 ();
 FILLCELL_X1 PHY_7226 ();
 FILLCELL_X1 PHY_7227 ();
 FILLCELL_X1 PHY_7228 ();
 FILLCELL_X1 PHY_7229 ();
 FILLCELL_X1 PHY_723 ();
 FILLCELL_X1 PHY_7230 ();
 FILLCELL_X1 PHY_7231 ();
 FILLCELL_X1 PHY_7232 ();
 FILLCELL_X1 PHY_7233 ();
 FILLCELL_X1 PHY_7234 ();
 FILLCELL_X1 PHY_7235 ();
 FILLCELL_X1 PHY_7236 ();
 FILLCELL_X1 PHY_7237 ();
 FILLCELL_X1 PHY_7238 ();
 FILLCELL_X1 PHY_7239 ();
 FILLCELL_X1 PHY_724 ();
 FILLCELL_X1 PHY_7240 ();
 FILLCELL_X1 PHY_7241 ();
 FILLCELL_X1 PHY_7242 ();
 FILLCELL_X1 PHY_7243 ();
 FILLCELL_X1 PHY_7244 ();
 FILLCELL_X1 PHY_7245 ();
 FILLCELL_X1 PHY_7246 ();
 FILLCELL_X1 PHY_7247 ();
 FILLCELL_X1 PHY_7248 ();
 FILLCELL_X1 PHY_7249 ();
 FILLCELL_X1 PHY_725 ();
 FILLCELL_X1 PHY_7250 ();
 FILLCELL_X1 PHY_7251 ();
 FILLCELL_X1 PHY_7252 ();
 FILLCELL_X1 PHY_7253 ();
 FILLCELL_X1 PHY_7254 ();
 FILLCELL_X1 PHY_7255 ();
 FILLCELL_X1 PHY_7256 ();
 FILLCELL_X1 PHY_7257 ();
 FILLCELL_X1 PHY_7258 ();
 FILLCELL_X1 PHY_7259 ();
 FILLCELL_X1 PHY_726 ();
 FILLCELL_X1 PHY_7260 ();
 FILLCELL_X1 PHY_7261 ();
 FILLCELL_X1 PHY_7262 ();
 FILLCELL_X1 PHY_7263 ();
 FILLCELL_X1 PHY_7264 ();
 FILLCELL_X1 PHY_7265 ();
 FILLCELL_X1 PHY_7266 ();
 FILLCELL_X1 PHY_7267 ();
 FILLCELL_X1 PHY_7268 ();
 FILLCELL_X1 PHY_7269 ();
 FILLCELL_X1 PHY_727 ();
 FILLCELL_X1 PHY_7270 ();
 FILLCELL_X1 PHY_7271 ();
 FILLCELL_X1 PHY_7272 ();
 FILLCELL_X1 PHY_7273 ();
 FILLCELL_X1 PHY_7274 ();
 FILLCELL_X1 PHY_7275 ();
 FILLCELL_X1 PHY_7276 ();
 FILLCELL_X1 PHY_7277 ();
 FILLCELL_X1 PHY_7278 ();
 FILLCELL_X1 PHY_7279 ();
 FILLCELL_X1 PHY_728 ();
 FILLCELL_X1 PHY_7280 ();
 FILLCELL_X1 PHY_7281 ();
 FILLCELL_X1 PHY_7282 ();
 FILLCELL_X1 PHY_7283 ();
 FILLCELL_X1 PHY_7284 ();
 FILLCELL_X1 PHY_7285 ();
 FILLCELL_X1 PHY_7286 ();
 FILLCELL_X1 PHY_7287 ();
 FILLCELL_X1 PHY_7288 ();
 FILLCELL_X1 PHY_7289 ();
 FILLCELL_X1 PHY_729 ();
 FILLCELL_X1 PHY_7290 ();
 FILLCELL_X1 PHY_7291 ();
 FILLCELL_X1 PHY_7292 ();
 FILLCELL_X1 PHY_7293 ();
 FILLCELL_X1 PHY_7294 ();
 FILLCELL_X1 PHY_7295 ();
 FILLCELL_X1 PHY_7296 ();
 FILLCELL_X1 PHY_7297 ();
 FILLCELL_X1 PHY_7298 ();
 FILLCELL_X1 PHY_7299 ();
 FILLCELL_X1 PHY_73 ();
 FILLCELL_X1 PHY_730 ();
 FILLCELL_X1 PHY_7300 ();
 FILLCELL_X1 PHY_7301 ();
 FILLCELL_X1 PHY_7302 ();
 FILLCELL_X1 PHY_7303 ();
 FILLCELL_X1 PHY_7304 ();
 FILLCELL_X1 PHY_7305 ();
 FILLCELL_X1 PHY_7306 ();
 FILLCELL_X1 PHY_7307 ();
 FILLCELL_X1 PHY_7308 ();
 FILLCELL_X1 PHY_7309 ();
 FILLCELL_X1 PHY_731 ();
 FILLCELL_X1 PHY_7310 ();
 FILLCELL_X1 PHY_7311 ();
 FILLCELL_X1 PHY_7312 ();
 FILLCELL_X1 PHY_7313 ();
 FILLCELL_X1 PHY_7314 ();
 FILLCELL_X1 PHY_7315 ();
 FILLCELL_X1 PHY_7316 ();
 FILLCELL_X1 PHY_7317 ();
 FILLCELL_X1 PHY_7318 ();
 FILLCELL_X1 PHY_7319 ();
 FILLCELL_X1 PHY_732 ();
 FILLCELL_X1 PHY_7320 ();
 FILLCELL_X1 PHY_7321 ();
 FILLCELL_X1 PHY_7322 ();
 FILLCELL_X1 PHY_7323 ();
 FILLCELL_X1 PHY_7324 ();
 FILLCELL_X1 PHY_7325 ();
 FILLCELL_X1 PHY_7326 ();
 FILLCELL_X1 PHY_7327 ();
 FILLCELL_X1 PHY_7328 ();
 FILLCELL_X1 PHY_7329 ();
 FILLCELL_X1 PHY_733 ();
 FILLCELL_X1 PHY_7330 ();
 FILLCELL_X1 PHY_7331 ();
 FILLCELL_X1 PHY_7332 ();
 FILLCELL_X1 PHY_7333 ();
 FILLCELL_X1 PHY_7334 ();
 FILLCELL_X1 PHY_7335 ();
 FILLCELL_X1 PHY_7336 ();
 FILLCELL_X1 PHY_7337 ();
 FILLCELL_X1 PHY_7338 ();
 FILLCELL_X1 PHY_7339 ();
 FILLCELL_X1 PHY_734 ();
 FILLCELL_X1 PHY_7340 ();
 FILLCELL_X1 PHY_7341 ();
 FILLCELL_X1 PHY_7342 ();
 FILLCELL_X1 PHY_7343 ();
 FILLCELL_X1 PHY_7344 ();
 FILLCELL_X1 PHY_7345 ();
 FILLCELL_X1 PHY_7346 ();
 FILLCELL_X1 PHY_7347 ();
 FILLCELL_X1 PHY_7348 ();
 FILLCELL_X1 PHY_7349 ();
 FILLCELL_X1 PHY_735 ();
 FILLCELL_X1 PHY_7350 ();
 FILLCELL_X1 PHY_7351 ();
 FILLCELL_X1 PHY_7352 ();
 FILLCELL_X1 PHY_7353 ();
 FILLCELL_X1 PHY_7354 ();
 FILLCELL_X1 PHY_7355 ();
 FILLCELL_X1 PHY_7356 ();
 FILLCELL_X1 PHY_7357 ();
 FILLCELL_X1 PHY_7358 ();
 FILLCELL_X1 PHY_7359 ();
 FILLCELL_X1 PHY_736 ();
 FILLCELL_X1 PHY_7360 ();
 FILLCELL_X1 PHY_7361 ();
 FILLCELL_X1 PHY_7362 ();
 FILLCELL_X1 PHY_7363 ();
 FILLCELL_X1 PHY_7364 ();
 FILLCELL_X1 PHY_7365 ();
 FILLCELL_X1 PHY_7366 ();
 FILLCELL_X1 PHY_7367 ();
 FILLCELL_X1 PHY_7368 ();
 FILLCELL_X1 PHY_7369 ();
 FILLCELL_X1 PHY_737 ();
 FILLCELL_X1 PHY_7370 ();
 FILLCELL_X1 PHY_7371 ();
 FILLCELL_X1 PHY_7372 ();
 FILLCELL_X1 PHY_7373 ();
 FILLCELL_X1 PHY_7374 ();
 FILLCELL_X1 PHY_7375 ();
 FILLCELL_X1 PHY_7376 ();
 FILLCELL_X1 PHY_7377 ();
 FILLCELL_X1 PHY_7378 ();
 FILLCELL_X1 PHY_7379 ();
 FILLCELL_X1 PHY_738 ();
 FILLCELL_X1 PHY_7380 ();
 FILLCELL_X1 PHY_7381 ();
 FILLCELL_X1 PHY_7382 ();
 FILLCELL_X1 PHY_7383 ();
 FILLCELL_X1 PHY_7384 ();
 FILLCELL_X1 PHY_7385 ();
 FILLCELL_X1 PHY_7386 ();
 FILLCELL_X1 PHY_7387 ();
 FILLCELL_X1 PHY_7388 ();
 FILLCELL_X1 PHY_7389 ();
 FILLCELL_X1 PHY_739 ();
 FILLCELL_X1 PHY_7390 ();
 FILLCELL_X1 PHY_7391 ();
 FILLCELL_X1 PHY_7392 ();
 FILLCELL_X1 PHY_7393 ();
 FILLCELL_X1 PHY_7394 ();
 FILLCELL_X1 PHY_7395 ();
 FILLCELL_X1 PHY_7396 ();
 FILLCELL_X1 PHY_7397 ();
 FILLCELL_X1 PHY_7398 ();
 FILLCELL_X1 PHY_7399 ();
 FILLCELL_X1 PHY_74 ();
 FILLCELL_X1 PHY_740 ();
 FILLCELL_X1 PHY_7400 ();
 FILLCELL_X1 PHY_7401 ();
 FILLCELL_X1 PHY_7402 ();
 FILLCELL_X1 PHY_7403 ();
 FILLCELL_X1 PHY_7404 ();
 FILLCELL_X1 PHY_7405 ();
 FILLCELL_X1 PHY_7406 ();
 FILLCELL_X1 PHY_7407 ();
 FILLCELL_X1 PHY_7408 ();
 FILLCELL_X1 PHY_7409 ();
 FILLCELL_X1 PHY_741 ();
 FILLCELL_X1 PHY_7410 ();
 FILLCELL_X1 PHY_7411 ();
 FILLCELL_X1 PHY_7412 ();
 FILLCELL_X1 PHY_7413 ();
 FILLCELL_X1 PHY_7414 ();
 FILLCELL_X1 PHY_7415 ();
 FILLCELL_X1 PHY_7416 ();
 FILLCELL_X1 PHY_7417 ();
 FILLCELL_X1 PHY_7418 ();
 FILLCELL_X1 PHY_7419 ();
 FILLCELL_X1 PHY_742 ();
 FILLCELL_X1 PHY_7420 ();
 FILLCELL_X1 PHY_7421 ();
 FILLCELL_X1 PHY_7422 ();
 FILLCELL_X1 PHY_7423 ();
 FILLCELL_X1 PHY_7424 ();
 FILLCELL_X1 PHY_7425 ();
 FILLCELL_X1 PHY_7426 ();
 FILLCELL_X1 PHY_7427 ();
 FILLCELL_X1 PHY_7428 ();
 FILLCELL_X1 PHY_7429 ();
 FILLCELL_X1 PHY_743 ();
 FILLCELL_X1 PHY_7430 ();
 FILLCELL_X1 PHY_7431 ();
 FILLCELL_X1 PHY_7432 ();
 FILLCELL_X1 PHY_7433 ();
 FILLCELL_X1 PHY_7434 ();
 FILLCELL_X1 PHY_7435 ();
 FILLCELL_X1 PHY_7436 ();
 FILLCELL_X1 PHY_7437 ();
 FILLCELL_X1 PHY_7438 ();
 FILLCELL_X1 PHY_7439 ();
 FILLCELL_X1 PHY_744 ();
 FILLCELL_X1 PHY_7440 ();
 FILLCELL_X1 PHY_7441 ();
 FILLCELL_X1 PHY_7442 ();
 FILLCELL_X1 PHY_7443 ();
 FILLCELL_X1 PHY_7444 ();
 FILLCELL_X1 PHY_7445 ();
 FILLCELL_X1 PHY_7446 ();
 FILLCELL_X1 PHY_7447 ();
 FILLCELL_X1 PHY_7448 ();
 FILLCELL_X1 PHY_7449 ();
 FILLCELL_X1 PHY_745 ();
 FILLCELL_X1 PHY_7450 ();
 FILLCELL_X1 PHY_7451 ();
 FILLCELL_X1 PHY_7452 ();
 FILLCELL_X1 PHY_7453 ();
 FILLCELL_X1 PHY_7454 ();
 FILLCELL_X1 PHY_7455 ();
 FILLCELL_X1 PHY_7456 ();
 FILLCELL_X1 PHY_7457 ();
 FILLCELL_X1 PHY_7458 ();
 FILLCELL_X1 PHY_7459 ();
 FILLCELL_X1 PHY_746 ();
 FILLCELL_X1 PHY_7460 ();
 FILLCELL_X1 PHY_7461 ();
 FILLCELL_X1 PHY_7462 ();
 FILLCELL_X1 PHY_7463 ();
 FILLCELL_X1 PHY_7464 ();
 FILLCELL_X1 PHY_7465 ();
 FILLCELL_X1 PHY_7466 ();
 FILLCELL_X1 PHY_7467 ();
 FILLCELL_X1 PHY_7468 ();
 FILLCELL_X1 PHY_7469 ();
 FILLCELL_X1 PHY_747 ();
 FILLCELL_X1 PHY_7470 ();
 FILLCELL_X1 PHY_7471 ();
 FILLCELL_X1 PHY_7472 ();
 FILLCELL_X1 PHY_7473 ();
 FILLCELL_X1 PHY_7474 ();
 FILLCELL_X1 PHY_7475 ();
 FILLCELL_X1 PHY_7476 ();
 FILLCELL_X1 PHY_7477 ();
 FILLCELL_X1 PHY_7478 ();
 FILLCELL_X1 PHY_7479 ();
 FILLCELL_X1 PHY_748 ();
 FILLCELL_X1 PHY_7480 ();
 FILLCELL_X1 PHY_7481 ();
 FILLCELL_X1 PHY_7482 ();
 FILLCELL_X1 PHY_7483 ();
 FILLCELL_X1 PHY_7484 ();
 FILLCELL_X1 PHY_7485 ();
 FILLCELL_X1 PHY_7486 ();
 FILLCELL_X1 PHY_7487 ();
 FILLCELL_X1 PHY_7488 ();
 FILLCELL_X1 PHY_7489 ();
 FILLCELL_X1 PHY_749 ();
 FILLCELL_X1 PHY_7490 ();
 FILLCELL_X1 PHY_7491 ();
 FILLCELL_X1 PHY_7492 ();
 FILLCELL_X1 PHY_7493 ();
 FILLCELL_X1 PHY_7494 ();
 FILLCELL_X1 PHY_7495 ();
 FILLCELL_X1 PHY_7496 ();
 FILLCELL_X1 PHY_7497 ();
 FILLCELL_X1 PHY_7498 ();
 FILLCELL_X1 PHY_7499 ();
 FILLCELL_X1 PHY_75 ();
 FILLCELL_X1 PHY_750 ();
 FILLCELL_X1 PHY_7500 ();
 FILLCELL_X1 PHY_7501 ();
 FILLCELL_X1 PHY_7502 ();
 FILLCELL_X1 PHY_7503 ();
 FILLCELL_X1 PHY_7504 ();
 FILLCELL_X1 PHY_7505 ();
 FILLCELL_X1 PHY_7506 ();
 FILLCELL_X1 PHY_7507 ();
 FILLCELL_X1 PHY_7508 ();
 FILLCELL_X1 PHY_7509 ();
 FILLCELL_X1 PHY_751 ();
 FILLCELL_X1 PHY_7510 ();
 FILLCELL_X1 PHY_7511 ();
 FILLCELL_X1 PHY_7512 ();
 FILLCELL_X1 PHY_7513 ();
 FILLCELL_X1 PHY_7514 ();
 FILLCELL_X1 PHY_7515 ();
 FILLCELL_X1 PHY_7516 ();
 FILLCELL_X1 PHY_7517 ();
 FILLCELL_X1 PHY_7518 ();
 FILLCELL_X1 PHY_7519 ();
 FILLCELL_X1 PHY_752 ();
 FILLCELL_X1 PHY_7520 ();
 FILLCELL_X1 PHY_7521 ();
 FILLCELL_X1 PHY_7522 ();
 FILLCELL_X1 PHY_7523 ();
 FILLCELL_X1 PHY_7524 ();
 FILLCELL_X1 PHY_7525 ();
 FILLCELL_X1 PHY_7526 ();
 FILLCELL_X1 PHY_7527 ();
 FILLCELL_X1 PHY_7528 ();
 FILLCELL_X1 PHY_7529 ();
 FILLCELL_X1 PHY_753 ();
 FILLCELL_X1 PHY_7530 ();
 FILLCELL_X1 PHY_7531 ();
 FILLCELL_X1 PHY_7532 ();
 FILLCELL_X1 PHY_7533 ();
 FILLCELL_X1 PHY_7534 ();
 FILLCELL_X1 PHY_7535 ();
 FILLCELL_X1 PHY_7536 ();
 FILLCELL_X1 PHY_7537 ();
 FILLCELL_X1 PHY_7538 ();
 FILLCELL_X1 PHY_7539 ();
 FILLCELL_X1 PHY_754 ();
 FILLCELL_X1 PHY_7540 ();
 FILLCELL_X1 PHY_7541 ();
 FILLCELL_X1 PHY_7542 ();
 FILLCELL_X1 PHY_7543 ();
 FILLCELL_X1 PHY_7544 ();
 FILLCELL_X1 PHY_7545 ();
 FILLCELL_X1 PHY_7546 ();
 FILLCELL_X1 PHY_7547 ();
 FILLCELL_X1 PHY_7548 ();
 FILLCELL_X1 PHY_7549 ();
 FILLCELL_X1 PHY_755 ();
 FILLCELL_X1 PHY_7550 ();
 FILLCELL_X1 PHY_7551 ();
 FILLCELL_X1 PHY_7552 ();
 FILLCELL_X1 PHY_7553 ();
 FILLCELL_X1 PHY_7554 ();
 FILLCELL_X1 PHY_7555 ();
 FILLCELL_X1 PHY_7556 ();
 FILLCELL_X1 PHY_7557 ();
 FILLCELL_X1 PHY_7558 ();
 FILLCELL_X1 PHY_7559 ();
 FILLCELL_X1 PHY_756 ();
 FILLCELL_X1 PHY_7560 ();
 FILLCELL_X1 PHY_7561 ();
 FILLCELL_X1 PHY_7562 ();
 FILLCELL_X1 PHY_7563 ();
 FILLCELL_X1 PHY_7564 ();
 FILLCELL_X1 PHY_7565 ();
 FILLCELL_X1 PHY_7566 ();
 FILLCELL_X1 PHY_7567 ();
 FILLCELL_X1 PHY_7568 ();
 FILLCELL_X1 PHY_7569 ();
 FILLCELL_X1 PHY_757 ();
 FILLCELL_X1 PHY_7570 ();
 FILLCELL_X1 PHY_7571 ();
 FILLCELL_X1 PHY_7572 ();
 FILLCELL_X1 PHY_7573 ();
 FILLCELL_X1 PHY_7574 ();
 FILLCELL_X1 PHY_7575 ();
 FILLCELL_X1 PHY_7576 ();
 FILLCELL_X1 PHY_7577 ();
 FILLCELL_X1 PHY_7578 ();
 FILLCELL_X1 PHY_7579 ();
 FILLCELL_X1 PHY_758 ();
 FILLCELL_X1 PHY_7580 ();
 FILLCELL_X1 PHY_7581 ();
 FILLCELL_X1 PHY_7582 ();
 FILLCELL_X1 PHY_7583 ();
 FILLCELL_X1 PHY_7584 ();
 FILLCELL_X1 PHY_7585 ();
 FILLCELL_X1 PHY_7586 ();
 FILLCELL_X1 PHY_7587 ();
 FILLCELL_X1 PHY_7588 ();
 FILLCELL_X1 PHY_7589 ();
 FILLCELL_X1 PHY_759 ();
 FILLCELL_X1 PHY_7590 ();
 FILLCELL_X1 PHY_7591 ();
 FILLCELL_X1 PHY_7592 ();
 FILLCELL_X1 PHY_7593 ();
 FILLCELL_X1 PHY_7594 ();
 FILLCELL_X1 PHY_7595 ();
 FILLCELL_X1 PHY_7596 ();
 FILLCELL_X1 PHY_7597 ();
 FILLCELL_X1 PHY_7598 ();
 FILLCELL_X1 PHY_7599 ();
 FILLCELL_X1 PHY_76 ();
 FILLCELL_X1 PHY_760 ();
 FILLCELL_X1 PHY_7600 ();
 FILLCELL_X1 PHY_7601 ();
 FILLCELL_X1 PHY_7602 ();
 FILLCELL_X1 PHY_7603 ();
 FILLCELL_X1 PHY_7604 ();
 FILLCELL_X1 PHY_7605 ();
 FILLCELL_X1 PHY_7606 ();
 FILLCELL_X1 PHY_7607 ();
 FILLCELL_X1 PHY_7608 ();
 FILLCELL_X1 PHY_7609 ();
 FILLCELL_X1 PHY_761 ();
 FILLCELL_X1 PHY_7610 ();
 FILLCELL_X1 PHY_7611 ();
 FILLCELL_X1 PHY_7612 ();
 FILLCELL_X1 PHY_7613 ();
 FILLCELL_X1 PHY_7614 ();
 FILLCELL_X1 PHY_7615 ();
 FILLCELL_X1 PHY_7616 ();
 FILLCELL_X1 PHY_7617 ();
 FILLCELL_X1 PHY_7618 ();
 FILLCELL_X1 PHY_7619 ();
 FILLCELL_X1 PHY_762 ();
 FILLCELL_X1 PHY_7620 ();
 FILLCELL_X1 PHY_7621 ();
 FILLCELL_X1 PHY_7622 ();
 FILLCELL_X1 PHY_7623 ();
 FILLCELL_X1 PHY_7624 ();
 FILLCELL_X1 PHY_7625 ();
 FILLCELL_X1 PHY_7626 ();
 FILLCELL_X1 PHY_7627 ();
 FILLCELL_X1 PHY_7628 ();
 FILLCELL_X1 PHY_7629 ();
 FILLCELL_X1 PHY_763 ();
 FILLCELL_X1 PHY_7630 ();
 FILLCELL_X1 PHY_7631 ();
 FILLCELL_X1 PHY_7632 ();
 FILLCELL_X1 PHY_7633 ();
 FILLCELL_X1 PHY_7634 ();
 FILLCELL_X1 PHY_7635 ();
 FILLCELL_X1 PHY_7636 ();
 FILLCELL_X1 PHY_7637 ();
 FILLCELL_X1 PHY_7638 ();
 FILLCELL_X1 PHY_7639 ();
 FILLCELL_X1 PHY_764 ();
 FILLCELL_X1 PHY_7640 ();
 FILLCELL_X1 PHY_7641 ();
 FILLCELL_X1 PHY_7642 ();
 FILLCELL_X1 PHY_7643 ();
 FILLCELL_X1 PHY_7644 ();
 FILLCELL_X1 PHY_7645 ();
 FILLCELL_X1 PHY_7646 ();
 FILLCELL_X1 PHY_7647 ();
 FILLCELL_X1 PHY_7648 ();
 FILLCELL_X1 PHY_7649 ();
 FILLCELL_X1 PHY_765 ();
 FILLCELL_X1 PHY_7650 ();
 FILLCELL_X1 PHY_7651 ();
 FILLCELL_X1 PHY_7652 ();
 FILLCELL_X1 PHY_7653 ();
 FILLCELL_X1 PHY_7654 ();
 FILLCELL_X1 PHY_7655 ();
 FILLCELL_X1 PHY_7656 ();
 FILLCELL_X1 PHY_7657 ();
 FILLCELL_X1 PHY_7658 ();
 FILLCELL_X1 PHY_7659 ();
 FILLCELL_X1 PHY_766 ();
 FILLCELL_X1 PHY_7660 ();
 FILLCELL_X1 PHY_7661 ();
 FILLCELL_X1 PHY_7662 ();
 FILLCELL_X1 PHY_7663 ();
 FILLCELL_X1 PHY_7664 ();
 FILLCELL_X1 PHY_7665 ();
 FILLCELL_X1 PHY_7666 ();
 FILLCELL_X1 PHY_7667 ();
 FILLCELL_X1 PHY_7668 ();
 FILLCELL_X1 PHY_7669 ();
 FILLCELL_X1 PHY_767 ();
 FILLCELL_X1 PHY_7670 ();
 FILLCELL_X1 PHY_7671 ();
 FILLCELL_X1 PHY_7672 ();
 FILLCELL_X1 PHY_7673 ();
 FILLCELL_X1 PHY_7674 ();
 FILLCELL_X1 PHY_7675 ();
 FILLCELL_X1 PHY_7676 ();
 FILLCELL_X1 PHY_7677 ();
 FILLCELL_X1 PHY_7678 ();
 FILLCELL_X1 PHY_7679 ();
 FILLCELL_X1 PHY_768 ();
 FILLCELL_X1 PHY_7680 ();
 FILLCELL_X1 PHY_7681 ();
 FILLCELL_X1 PHY_7682 ();
 FILLCELL_X1 PHY_7683 ();
 FILLCELL_X1 PHY_7684 ();
 FILLCELL_X1 PHY_7685 ();
 FILLCELL_X1 PHY_7686 ();
 FILLCELL_X1 PHY_7687 ();
 FILLCELL_X1 PHY_7688 ();
 FILLCELL_X1 PHY_7689 ();
 FILLCELL_X1 PHY_769 ();
 FILLCELL_X1 PHY_7690 ();
 FILLCELL_X1 PHY_7691 ();
 FILLCELL_X1 PHY_7692 ();
 FILLCELL_X1 PHY_7693 ();
 FILLCELL_X1 PHY_7694 ();
 FILLCELL_X1 PHY_7695 ();
 FILLCELL_X1 PHY_7696 ();
 FILLCELL_X1 PHY_7697 ();
 FILLCELL_X1 PHY_7698 ();
 FILLCELL_X1 PHY_7699 ();
 FILLCELL_X1 PHY_77 ();
 FILLCELL_X1 PHY_770 ();
 FILLCELL_X1 PHY_7700 ();
 FILLCELL_X1 PHY_7701 ();
 FILLCELL_X1 PHY_7702 ();
 FILLCELL_X1 PHY_7703 ();
 FILLCELL_X1 PHY_7704 ();
 FILLCELL_X1 PHY_7705 ();
 FILLCELL_X1 PHY_7706 ();
 FILLCELL_X1 PHY_7707 ();
 FILLCELL_X1 PHY_7708 ();
 FILLCELL_X1 PHY_7709 ();
 FILLCELL_X1 PHY_771 ();
 FILLCELL_X1 PHY_7710 ();
 FILLCELL_X1 PHY_7711 ();
 FILLCELL_X1 PHY_7712 ();
 FILLCELL_X1 PHY_7713 ();
 FILLCELL_X1 PHY_7714 ();
 FILLCELL_X1 PHY_7715 ();
 FILLCELL_X1 PHY_7716 ();
 FILLCELL_X1 PHY_7717 ();
 FILLCELL_X1 PHY_7718 ();
 FILLCELL_X1 PHY_7719 ();
 FILLCELL_X1 PHY_772 ();
 FILLCELL_X1 PHY_7720 ();
 FILLCELL_X1 PHY_7721 ();
 FILLCELL_X1 PHY_7722 ();
 FILLCELL_X1 PHY_7723 ();
 FILLCELL_X1 PHY_7724 ();
 FILLCELL_X1 PHY_7725 ();
 FILLCELL_X1 PHY_7726 ();
 FILLCELL_X1 PHY_7727 ();
 FILLCELL_X1 PHY_7728 ();
 FILLCELL_X1 PHY_7729 ();
 FILLCELL_X1 PHY_773 ();
 FILLCELL_X1 PHY_7730 ();
 FILLCELL_X1 PHY_7731 ();
 FILLCELL_X1 PHY_7732 ();
 FILLCELL_X1 PHY_7733 ();
 FILLCELL_X1 PHY_7734 ();
 FILLCELL_X1 PHY_7735 ();
 FILLCELL_X1 PHY_7736 ();
 FILLCELL_X1 PHY_7737 ();
 FILLCELL_X1 PHY_7738 ();
 FILLCELL_X1 PHY_7739 ();
 FILLCELL_X1 PHY_774 ();
 FILLCELL_X1 PHY_7740 ();
 FILLCELL_X1 PHY_7741 ();
 FILLCELL_X1 PHY_7742 ();
 FILLCELL_X1 PHY_7743 ();
 FILLCELL_X1 PHY_7744 ();
 FILLCELL_X1 PHY_7745 ();
 FILLCELL_X1 PHY_7746 ();
 FILLCELL_X1 PHY_7747 ();
 FILLCELL_X1 PHY_7748 ();
 FILLCELL_X1 PHY_7749 ();
 FILLCELL_X1 PHY_775 ();
 FILLCELL_X1 PHY_7750 ();
 FILLCELL_X1 PHY_7751 ();
 FILLCELL_X1 PHY_7752 ();
 FILLCELL_X1 PHY_7753 ();
 FILLCELL_X1 PHY_7754 ();
 FILLCELL_X1 PHY_7755 ();
 FILLCELL_X1 PHY_7756 ();
 FILLCELL_X1 PHY_7757 ();
 FILLCELL_X1 PHY_7758 ();
 FILLCELL_X1 PHY_7759 ();
 FILLCELL_X1 PHY_776 ();
 FILLCELL_X1 PHY_7760 ();
 FILLCELL_X1 PHY_7761 ();
 FILLCELL_X1 PHY_7762 ();
 FILLCELL_X1 PHY_7763 ();
 FILLCELL_X1 PHY_7764 ();
 FILLCELL_X1 PHY_7765 ();
 FILLCELL_X1 PHY_7766 ();
 FILLCELL_X1 PHY_7767 ();
 FILLCELL_X1 PHY_7768 ();
 FILLCELL_X1 PHY_7769 ();
 FILLCELL_X1 PHY_777 ();
 FILLCELL_X1 PHY_7770 ();
 FILLCELL_X1 PHY_7771 ();
 FILLCELL_X1 PHY_7772 ();
 FILLCELL_X1 PHY_7773 ();
 FILLCELL_X1 PHY_7774 ();
 FILLCELL_X1 PHY_7775 ();
 FILLCELL_X1 PHY_7776 ();
 FILLCELL_X1 PHY_7777 ();
 FILLCELL_X1 PHY_7778 ();
 FILLCELL_X1 PHY_7779 ();
 FILLCELL_X1 PHY_778 ();
 FILLCELL_X1 PHY_7780 ();
 FILLCELL_X1 PHY_7781 ();
 FILLCELL_X1 PHY_7782 ();
 FILLCELL_X1 PHY_7783 ();
 FILLCELL_X1 PHY_7784 ();
 FILLCELL_X1 PHY_7785 ();
 FILLCELL_X1 PHY_7786 ();
 FILLCELL_X1 PHY_7787 ();
 FILLCELL_X1 PHY_7788 ();
 FILLCELL_X1 PHY_7789 ();
 FILLCELL_X1 PHY_779 ();
 FILLCELL_X1 PHY_7790 ();
 FILLCELL_X1 PHY_7791 ();
 FILLCELL_X1 PHY_7792 ();
 FILLCELL_X1 PHY_7793 ();
 FILLCELL_X1 PHY_7794 ();
 FILLCELL_X1 PHY_7795 ();
 FILLCELL_X1 PHY_7796 ();
 FILLCELL_X1 PHY_7797 ();
 FILLCELL_X1 PHY_7798 ();
 FILLCELL_X1 PHY_7799 ();
 FILLCELL_X1 PHY_78 ();
 FILLCELL_X1 PHY_780 ();
 FILLCELL_X1 PHY_7800 ();
 FILLCELL_X1 PHY_7801 ();
 FILLCELL_X1 PHY_7802 ();
 FILLCELL_X1 PHY_7803 ();
 FILLCELL_X1 PHY_7804 ();
 FILLCELL_X1 PHY_7805 ();
 FILLCELL_X1 PHY_7806 ();
 FILLCELL_X1 PHY_7807 ();
 FILLCELL_X1 PHY_7808 ();
 FILLCELL_X1 PHY_7809 ();
 FILLCELL_X1 PHY_781 ();
 FILLCELL_X1 PHY_7810 ();
 FILLCELL_X1 PHY_7811 ();
 FILLCELL_X1 PHY_7812 ();
 FILLCELL_X1 PHY_7813 ();
 FILLCELL_X1 PHY_7814 ();
 FILLCELL_X1 PHY_7815 ();
 FILLCELL_X1 PHY_7816 ();
 FILLCELL_X1 PHY_7817 ();
 FILLCELL_X1 PHY_7818 ();
 FILLCELL_X1 PHY_7819 ();
 FILLCELL_X1 PHY_782 ();
 FILLCELL_X1 PHY_7820 ();
 FILLCELL_X1 PHY_7821 ();
 FILLCELL_X1 PHY_7822 ();
 FILLCELL_X1 PHY_7823 ();
 FILLCELL_X1 PHY_7824 ();
 FILLCELL_X1 PHY_7825 ();
 FILLCELL_X1 PHY_7826 ();
 FILLCELL_X1 PHY_7827 ();
 FILLCELL_X1 PHY_7828 ();
 FILLCELL_X1 PHY_7829 ();
 FILLCELL_X1 PHY_783 ();
 FILLCELL_X1 PHY_7830 ();
 FILLCELL_X1 PHY_7831 ();
 FILLCELL_X1 PHY_7832 ();
 FILLCELL_X1 PHY_7833 ();
 FILLCELL_X1 PHY_7834 ();
 FILLCELL_X1 PHY_7835 ();
 FILLCELL_X1 PHY_7836 ();
 FILLCELL_X1 PHY_7837 ();
 FILLCELL_X1 PHY_7838 ();
 FILLCELL_X1 PHY_7839 ();
 FILLCELL_X1 PHY_784 ();
 FILLCELL_X1 PHY_7840 ();
 FILLCELL_X1 PHY_7841 ();
 FILLCELL_X1 PHY_7842 ();
 FILLCELL_X1 PHY_7843 ();
 FILLCELL_X1 PHY_7844 ();
 FILLCELL_X1 PHY_7845 ();
 FILLCELL_X1 PHY_7846 ();
 FILLCELL_X1 PHY_7847 ();
 FILLCELL_X1 PHY_7848 ();
 FILLCELL_X1 PHY_7849 ();
 FILLCELL_X1 PHY_785 ();
 FILLCELL_X1 PHY_7850 ();
 FILLCELL_X1 PHY_7851 ();
 FILLCELL_X1 PHY_7852 ();
 FILLCELL_X1 PHY_7853 ();
 FILLCELL_X1 PHY_7854 ();
 FILLCELL_X1 PHY_7855 ();
 FILLCELL_X1 PHY_7856 ();
 FILLCELL_X1 PHY_7857 ();
 FILLCELL_X1 PHY_7858 ();
 FILLCELL_X1 PHY_7859 ();
 FILLCELL_X1 PHY_786 ();
 FILLCELL_X1 PHY_7860 ();
 FILLCELL_X1 PHY_7861 ();
 FILLCELL_X1 PHY_7862 ();
 FILLCELL_X1 PHY_7863 ();
 FILLCELL_X1 PHY_7864 ();
 FILLCELL_X1 PHY_7865 ();
 FILLCELL_X1 PHY_7866 ();
 FILLCELL_X1 PHY_7867 ();
 FILLCELL_X1 PHY_7868 ();
 FILLCELL_X1 PHY_7869 ();
 FILLCELL_X1 PHY_787 ();
 FILLCELL_X1 PHY_7870 ();
 FILLCELL_X1 PHY_7871 ();
 FILLCELL_X1 PHY_7872 ();
 FILLCELL_X1 PHY_7873 ();
 FILLCELL_X1 PHY_7874 ();
 FILLCELL_X1 PHY_7875 ();
 FILLCELL_X1 PHY_7876 ();
 FILLCELL_X1 PHY_7877 ();
 FILLCELL_X1 PHY_7878 ();
 FILLCELL_X1 PHY_7879 ();
 FILLCELL_X1 PHY_788 ();
 FILLCELL_X1 PHY_7880 ();
 FILLCELL_X1 PHY_7881 ();
 FILLCELL_X1 PHY_7882 ();
 FILLCELL_X1 PHY_7883 ();
 FILLCELL_X1 PHY_7884 ();
 FILLCELL_X1 PHY_7885 ();
 FILLCELL_X1 PHY_7886 ();
 FILLCELL_X1 PHY_7887 ();
 FILLCELL_X1 PHY_7888 ();
 FILLCELL_X1 PHY_7889 ();
 FILLCELL_X1 PHY_789 ();
 FILLCELL_X1 PHY_7890 ();
 FILLCELL_X1 PHY_7891 ();
 FILLCELL_X1 PHY_7892 ();
 FILLCELL_X1 PHY_7893 ();
 FILLCELL_X1 PHY_7894 ();
 FILLCELL_X1 PHY_7895 ();
 FILLCELL_X1 PHY_7896 ();
 FILLCELL_X1 PHY_7897 ();
 FILLCELL_X1 PHY_7898 ();
 FILLCELL_X1 PHY_7899 ();
 FILLCELL_X1 PHY_79 ();
 FILLCELL_X1 PHY_790 ();
 FILLCELL_X1 PHY_7900 ();
 FILLCELL_X1 PHY_7901 ();
 FILLCELL_X1 PHY_7902 ();
 FILLCELL_X1 PHY_7903 ();
 FILLCELL_X1 PHY_7904 ();
 FILLCELL_X1 PHY_7905 ();
 FILLCELL_X1 PHY_7906 ();
 FILLCELL_X1 PHY_7907 ();
 FILLCELL_X1 PHY_7908 ();
 FILLCELL_X1 PHY_7909 ();
 FILLCELL_X1 PHY_791 ();
 FILLCELL_X1 PHY_7910 ();
 FILLCELL_X1 PHY_7911 ();
 FILLCELL_X1 PHY_7912 ();
 FILLCELL_X1 PHY_7913 ();
 FILLCELL_X1 PHY_7914 ();
 FILLCELL_X1 PHY_7915 ();
 FILLCELL_X1 PHY_7916 ();
 FILLCELL_X1 PHY_7917 ();
 FILLCELL_X1 PHY_7918 ();
 FILLCELL_X1 PHY_7919 ();
 FILLCELL_X1 PHY_792 ();
 FILLCELL_X1 PHY_7920 ();
 FILLCELL_X1 PHY_7921 ();
 FILLCELL_X1 PHY_7922 ();
 FILLCELL_X1 PHY_7923 ();
 FILLCELL_X1 PHY_7924 ();
 FILLCELL_X1 PHY_7925 ();
 FILLCELL_X1 PHY_7926 ();
 FILLCELL_X1 PHY_7927 ();
 FILLCELL_X1 PHY_7928 ();
 FILLCELL_X1 PHY_7929 ();
 FILLCELL_X1 PHY_793 ();
 FILLCELL_X1 PHY_7930 ();
 FILLCELL_X1 PHY_7931 ();
 FILLCELL_X1 PHY_7932 ();
 FILLCELL_X1 PHY_7933 ();
 FILLCELL_X1 PHY_7934 ();
 FILLCELL_X1 PHY_7935 ();
 FILLCELL_X1 PHY_7936 ();
 FILLCELL_X1 PHY_7937 ();
 FILLCELL_X1 PHY_7938 ();
 FILLCELL_X1 PHY_7939 ();
 FILLCELL_X1 PHY_794 ();
 FILLCELL_X1 PHY_7940 ();
 FILLCELL_X1 PHY_7941 ();
 FILLCELL_X1 PHY_7942 ();
 FILLCELL_X1 PHY_7943 ();
 FILLCELL_X1 PHY_7944 ();
 FILLCELL_X1 PHY_7945 ();
 FILLCELL_X1 PHY_7946 ();
 FILLCELL_X1 PHY_7947 ();
 FILLCELL_X1 PHY_7948 ();
 FILLCELL_X1 PHY_7949 ();
 FILLCELL_X1 PHY_795 ();
 FILLCELL_X1 PHY_7950 ();
 FILLCELL_X1 PHY_7951 ();
 FILLCELL_X1 PHY_7952 ();
 FILLCELL_X1 PHY_7953 ();
 FILLCELL_X1 PHY_7954 ();
 FILLCELL_X1 PHY_7955 ();
 FILLCELL_X1 PHY_7956 ();
 FILLCELL_X1 PHY_7957 ();
 FILLCELL_X1 PHY_7958 ();
 FILLCELL_X1 PHY_7959 ();
 FILLCELL_X1 PHY_796 ();
 FILLCELL_X1 PHY_7960 ();
 FILLCELL_X1 PHY_7961 ();
 FILLCELL_X1 PHY_7962 ();
 FILLCELL_X1 PHY_7963 ();
 FILLCELL_X1 PHY_7964 ();
 FILLCELL_X1 PHY_7965 ();
 FILLCELL_X1 PHY_7966 ();
 FILLCELL_X1 PHY_7967 ();
 FILLCELL_X1 PHY_7968 ();
 FILLCELL_X1 PHY_7969 ();
 FILLCELL_X1 PHY_797 ();
 FILLCELL_X1 PHY_7970 ();
 FILLCELL_X1 PHY_7971 ();
 FILLCELL_X1 PHY_7972 ();
 FILLCELL_X1 PHY_7973 ();
 FILLCELL_X1 PHY_7974 ();
 FILLCELL_X1 PHY_7975 ();
 FILLCELL_X1 PHY_7976 ();
 FILLCELL_X1 PHY_7977 ();
 FILLCELL_X1 PHY_7978 ();
 FILLCELL_X1 PHY_7979 ();
 FILLCELL_X1 PHY_798 ();
 FILLCELL_X1 PHY_7980 ();
 FILLCELL_X1 PHY_7981 ();
 FILLCELL_X1 PHY_7982 ();
 FILLCELL_X1 PHY_7983 ();
 FILLCELL_X1 PHY_7984 ();
 FILLCELL_X1 PHY_7985 ();
 FILLCELL_X1 PHY_7986 ();
 FILLCELL_X1 PHY_7987 ();
 FILLCELL_X1 PHY_7988 ();
 FILLCELL_X1 PHY_7989 ();
 FILLCELL_X1 PHY_799 ();
 FILLCELL_X1 PHY_7990 ();
 FILLCELL_X1 PHY_7991 ();
 FILLCELL_X1 PHY_7992 ();
 FILLCELL_X1 PHY_7993 ();
 FILLCELL_X1 PHY_7994 ();
 FILLCELL_X1 PHY_7995 ();
 FILLCELL_X1 PHY_7996 ();
 FILLCELL_X1 PHY_7997 ();
 FILLCELL_X1 PHY_7998 ();
 FILLCELL_X1 PHY_7999 ();
 FILLCELL_X1 PHY_8 ();
 FILLCELL_X1 PHY_80 ();
 FILLCELL_X1 PHY_800 ();
 FILLCELL_X1 PHY_8000 ();
 FILLCELL_X1 PHY_8001 ();
 FILLCELL_X1 PHY_8002 ();
 FILLCELL_X1 PHY_8003 ();
 FILLCELL_X1 PHY_8004 ();
 FILLCELL_X1 PHY_8005 ();
 FILLCELL_X1 PHY_8006 ();
 FILLCELL_X1 PHY_8007 ();
 FILLCELL_X1 PHY_8008 ();
 FILLCELL_X1 PHY_8009 ();
 FILLCELL_X1 PHY_801 ();
 FILLCELL_X1 PHY_8010 ();
 FILLCELL_X1 PHY_8011 ();
 FILLCELL_X1 PHY_8012 ();
 FILLCELL_X1 PHY_8013 ();
 FILLCELL_X1 PHY_8014 ();
 FILLCELL_X1 PHY_8015 ();
 FILLCELL_X1 PHY_8016 ();
 FILLCELL_X1 PHY_8017 ();
 FILLCELL_X1 PHY_8018 ();
 FILLCELL_X1 PHY_8019 ();
 FILLCELL_X1 PHY_802 ();
 FILLCELL_X1 PHY_8020 ();
 FILLCELL_X1 PHY_8021 ();
 FILLCELL_X1 PHY_8022 ();
 FILLCELL_X1 PHY_8023 ();
 FILLCELL_X1 PHY_8024 ();
 FILLCELL_X1 PHY_8025 ();
 FILLCELL_X1 PHY_8026 ();
 FILLCELL_X1 PHY_8027 ();
 FILLCELL_X1 PHY_8028 ();
 FILLCELL_X1 PHY_8029 ();
 FILLCELL_X1 PHY_803 ();
 FILLCELL_X1 PHY_8030 ();
 FILLCELL_X1 PHY_8031 ();
 FILLCELL_X1 PHY_8032 ();
 FILLCELL_X1 PHY_8033 ();
 FILLCELL_X1 PHY_8034 ();
 FILLCELL_X1 PHY_8035 ();
 FILLCELL_X1 PHY_804 ();
 FILLCELL_X1 PHY_805 ();
 FILLCELL_X1 PHY_806 ();
 FILLCELL_X1 PHY_807 ();
 FILLCELL_X1 PHY_808 ();
 FILLCELL_X1 PHY_809 ();
 FILLCELL_X1 PHY_81 ();
 FILLCELL_X1 PHY_810 ();
 FILLCELL_X1 PHY_811 ();
 FILLCELL_X1 PHY_812 ();
 FILLCELL_X1 PHY_813 ();
 FILLCELL_X1 PHY_814 ();
 FILLCELL_X1 PHY_815 ();
 FILLCELL_X1 PHY_816 ();
 FILLCELL_X1 PHY_817 ();
 FILLCELL_X1 PHY_818 ();
 FILLCELL_X1 PHY_819 ();
 FILLCELL_X1 PHY_82 ();
 FILLCELL_X1 PHY_820 ();
 FILLCELL_X1 PHY_821 ();
 FILLCELL_X1 PHY_822 ();
 FILLCELL_X1 PHY_823 ();
 FILLCELL_X1 PHY_824 ();
 FILLCELL_X1 PHY_825 ();
 FILLCELL_X1 PHY_826 ();
 FILLCELL_X1 PHY_827 ();
 FILLCELL_X1 PHY_828 ();
 FILLCELL_X1 PHY_829 ();
 FILLCELL_X1 PHY_83 ();
 FILLCELL_X1 PHY_830 ();
 FILLCELL_X1 PHY_831 ();
 FILLCELL_X1 PHY_832 ();
 FILLCELL_X1 PHY_833 ();
 FILLCELL_X1 PHY_834 ();
 FILLCELL_X1 PHY_835 ();
 FILLCELL_X1 PHY_836 ();
 FILLCELL_X1 PHY_837 ();
 FILLCELL_X1 PHY_838 ();
 FILLCELL_X1 PHY_839 ();
 FILLCELL_X1 PHY_84 ();
 FILLCELL_X1 PHY_840 ();
 FILLCELL_X1 PHY_841 ();
 FILLCELL_X1 PHY_842 ();
 FILLCELL_X1 PHY_843 ();
 FILLCELL_X1 PHY_844 ();
 FILLCELL_X1 PHY_845 ();
 FILLCELL_X1 PHY_846 ();
 FILLCELL_X1 PHY_847 ();
 FILLCELL_X1 PHY_848 ();
 FILLCELL_X1 PHY_849 ();
 FILLCELL_X1 PHY_85 ();
 FILLCELL_X1 PHY_850 ();
 FILLCELL_X1 PHY_851 ();
 FILLCELL_X1 PHY_852 ();
 FILLCELL_X1 PHY_853 ();
 FILLCELL_X1 PHY_854 ();
 FILLCELL_X1 PHY_855 ();
 FILLCELL_X1 PHY_856 ();
 FILLCELL_X1 PHY_857 ();
 FILLCELL_X1 PHY_858 ();
 FILLCELL_X1 PHY_859 ();
 FILLCELL_X1 PHY_86 ();
 FILLCELL_X1 PHY_860 ();
 FILLCELL_X1 PHY_861 ();
 FILLCELL_X1 PHY_862 ();
 FILLCELL_X1 PHY_863 ();
 FILLCELL_X1 PHY_864 ();
 FILLCELL_X1 PHY_865 ();
 FILLCELL_X1 PHY_866 ();
 FILLCELL_X1 PHY_867 ();
 FILLCELL_X1 PHY_868 ();
 FILLCELL_X1 PHY_869 ();
 FILLCELL_X1 PHY_87 ();
 FILLCELL_X1 PHY_870 ();
 FILLCELL_X1 PHY_871 ();
 FILLCELL_X1 PHY_872 ();
 FILLCELL_X1 PHY_873 ();
 FILLCELL_X1 PHY_874 ();
 FILLCELL_X1 PHY_875 ();
 FILLCELL_X1 PHY_876 ();
 FILLCELL_X1 PHY_877 ();
 FILLCELL_X1 PHY_878 ();
 FILLCELL_X1 PHY_879 ();
 FILLCELL_X1 PHY_88 ();
 FILLCELL_X1 PHY_880 ();
 FILLCELL_X1 PHY_881 ();
 FILLCELL_X1 PHY_882 ();
 FILLCELL_X1 PHY_883 ();
 FILLCELL_X1 PHY_884 ();
 FILLCELL_X1 PHY_885 ();
 FILLCELL_X1 PHY_886 ();
 FILLCELL_X1 PHY_887 ();
 FILLCELL_X1 PHY_888 ();
 FILLCELL_X1 PHY_889 ();
 FILLCELL_X1 PHY_89 ();
 FILLCELL_X1 PHY_890 ();
 FILLCELL_X1 PHY_891 ();
 FILLCELL_X1 PHY_892 ();
 FILLCELL_X1 PHY_893 ();
 FILLCELL_X1 PHY_894 ();
 FILLCELL_X1 PHY_895 ();
 FILLCELL_X1 PHY_896 ();
 FILLCELL_X1 PHY_897 ();
 FILLCELL_X1 PHY_898 ();
 FILLCELL_X1 PHY_899 ();
 FILLCELL_X1 PHY_9 ();
 FILLCELL_X1 PHY_90 ();
 FILLCELL_X1 PHY_900 ();
 FILLCELL_X1 PHY_901 ();
 FILLCELL_X1 PHY_902 ();
 FILLCELL_X1 PHY_903 ();
 FILLCELL_X1 PHY_904 ();
 FILLCELL_X1 PHY_905 ();
 FILLCELL_X1 PHY_906 ();
 FILLCELL_X1 PHY_907 ();
 FILLCELL_X1 PHY_908 ();
 FILLCELL_X1 PHY_909 ();
 FILLCELL_X1 PHY_91 ();
 FILLCELL_X1 PHY_910 ();
 FILLCELL_X1 PHY_911 ();
 FILLCELL_X1 PHY_912 ();
 FILLCELL_X1 PHY_913 ();
 FILLCELL_X1 PHY_914 ();
 FILLCELL_X1 PHY_915 ();
 FILLCELL_X1 PHY_916 ();
 FILLCELL_X1 PHY_917 ();
 FILLCELL_X1 PHY_918 ();
 FILLCELL_X1 PHY_919 ();
 FILLCELL_X1 PHY_92 ();
 FILLCELL_X1 PHY_920 ();
 FILLCELL_X1 PHY_921 ();
 FILLCELL_X1 PHY_922 ();
 FILLCELL_X1 PHY_923 ();
 FILLCELL_X1 PHY_924 ();
 FILLCELL_X1 PHY_925 ();
 FILLCELL_X1 PHY_926 ();
 FILLCELL_X1 PHY_927 ();
 FILLCELL_X1 PHY_928 ();
 FILLCELL_X1 PHY_929 ();
 FILLCELL_X1 PHY_93 ();
 FILLCELL_X1 PHY_930 ();
 FILLCELL_X1 PHY_931 ();
 FILLCELL_X1 PHY_932 ();
 FILLCELL_X1 PHY_933 ();
 FILLCELL_X1 PHY_934 ();
 FILLCELL_X1 PHY_935 ();
 FILLCELL_X1 PHY_936 ();
 FILLCELL_X1 PHY_937 ();
 FILLCELL_X1 PHY_938 ();
 FILLCELL_X1 PHY_939 ();
 FILLCELL_X1 PHY_94 ();
 FILLCELL_X1 PHY_940 ();
 FILLCELL_X1 PHY_941 ();
 FILLCELL_X1 PHY_942 ();
 FILLCELL_X1 PHY_943 ();
 FILLCELL_X1 PHY_944 ();
 FILLCELL_X1 PHY_945 ();
 FILLCELL_X1 PHY_946 ();
 FILLCELL_X1 PHY_947 ();
 FILLCELL_X1 PHY_948 ();
 FILLCELL_X1 PHY_949 ();
 FILLCELL_X1 PHY_95 ();
 FILLCELL_X1 PHY_950 ();
 FILLCELL_X1 PHY_951 ();
 FILLCELL_X1 PHY_952 ();
 FILLCELL_X1 PHY_953 ();
 FILLCELL_X1 PHY_954 ();
 FILLCELL_X1 PHY_955 ();
 FILLCELL_X1 PHY_956 ();
 FILLCELL_X1 PHY_957 ();
 FILLCELL_X1 PHY_958 ();
 FILLCELL_X1 PHY_959 ();
 FILLCELL_X1 PHY_96 ();
 FILLCELL_X1 PHY_960 ();
 FILLCELL_X1 PHY_961 ();
 FILLCELL_X1 PHY_962 ();
 FILLCELL_X1 PHY_963 ();
 FILLCELL_X1 PHY_964 ();
 FILLCELL_X1 PHY_965 ();
 FILLCELL_X1 PHY_966 ();
 FILLCELL_X1 PHY_967 ();
 FILLCELL_X1 PHY_968 ();
 FILLCELL_X1 PHY_969 ();
 FILLCELL_X1 PHY_97 ();
 FILLCELL_X1 PHY_970 ();
 FILLCELL_X1 PHY_971 ();
 FILLCELL_X1 PHY_972 ();
 FILLCELL_X1 PHY_973 ();
 FILLCELL_X1 PHY_974 ();
 FILLCELL_X1 PHY_975 ();
 FILLCELL_X1 PHY_976 ();
 FILLCELL_X1 PHY_977 ();
 FILLCELL_X1 PHY_978 ();
 FILLCELL_X1 PHY_979 ();
 FILLCELL_X1 PHY_98 ();
 FILLCELL_X1 PHY_980 ();
 FILLCELL_X1 PHY_981 ();
 FILLCELL_X1 PHY_982 ();
 FILLCELL_X1 PHY_983 ();
 FILLCELL_X1 PHY_984 ();
 FILLCELL_X1 PHY_985 ();
 FILLCELL_X1 PHY_986 ();
 FILLCELL_X1 PHY_987 ();
 FILLCELL_X1 PHY_988 ();
 FILLCELL_X1 PHY_989 ();
 FILLCELL_X1 PHY_99 ();
 FILLCELL_X1 PHY_990 ();
 FILLCELL_X1 PHY_991 ();
 FILLCELL_X1 PHY_992 ();
 FILLCELL_X1 PHY_993 ();
 FILLCELL_X1 PHY_994 ();
 FILLCELL_X1 PHY_995 ();
 FILLCELL_X1 PHY_996 ();
 FILLCELL_X1 PHY_997 ();
 FILLCELL_X1 PHY_998 ();
 FILLCELL_X1 PHY_999 ();
 BUF_X16 _32514_ (.A(\icache.N10 ),
    .Z(_07048_));
 INV_X2 _32515_ (.A(\icache.addr_tv_r [29]),
    .ZN(_07049_));
 BUF_X16 _32516_ (.A(_07049_),
    .Z(_07050_));
 NOR2_X1 _32517_ (.A1(_07050_),
    .A2(net1279),
    .ZN(_07051_));
 INV_X16 _32518_ (.A(net1371),
    .ZN(_07052_));
 AOI21_X1 _32519_ (.A(_07051_),
    .B1(_07052_),
    .B2(net1298),
    .ZN(_07053_));
 INV_X4 _32520_ (.A(net1353),
    .ZN(_07054_));
 BUF_X8 _32521_ (.A(_07054_),
    .Z(_07055_));
 NAND2_X1 _32522_ (.A1(_07055_),
    .A2(net1289),
    .ZN(_07056_));
 INV_X8 _32523_ (.A(\icache.addr_tv_r [25]),
    .ZN(_07057_));
 NOR2_X1 _32524_ (.A1(_07057_),
    .A2(net1287),
    .ZN(_07058_));
 INV_X8 _32525_ (.A(net1356),
    .ZN(_07059_));
 AND2_X1 _32526_ (.A1(_07059_),
    .A2(net1291),
    .ZN(_07060_));
 NOR2_X1 _32527_ (.A1(_07059_),
    .A2(net1291),
    .ZN(_07061_));
 INV_X2 _32528_ (.A(net1380),
    .ZN(_07062_));
 NOR2_X1 _32529_ (.A1(_07062_),
    .A2(net1302),
    .ZN(_07063_));
 NOR4_X1 _32530_ (.A1(_07058_),
    .A2(_07060_),
    .A3(_07061_),
    .A4(_07063_),
    .ZN(_07064_));
 BUF_X8 _32531_ (.A(_07062_),
    .Z(_07065_));
 NAND2_X1 _32532_ (.A1(_07065_),
    .A2(net1302),
    .ZN(_07066_));
 INV_X8 _32533_ (.A(net1374),
    .ZN(_07067_));
 INV_X8 _32534_ (.A(net1361),
    .ZN(_07068_));
 BUF_X16 _32535_ (.A(_07068_),
    .Z(_07069_));
 AOI22_X1 _32536_ (.A1(_07067_),
    .A2(net1300),
    .B1(_07069_),
    .B2(net1294),
    .ZN(_07070_));
 AND4_X1 _32537_ (.A1(_07056_),
    .A2(_07064_),
    .A3(_07066_),
    .A4(_07070_),
    .ZN(_07071_));
 INV_X8 _32538_ (.A(net1317),
    .ZN(_07072_));
 OR2_X1 _32539_ (.A1(_07072_),
    .A2(net1272),
    .ZN(_07073_));
 INV_X2 _32540_ (.A(net1330),
    .ZN(_07074_));
 AND2_X1 _32541_ (.A1(_07074_),
    .A2(net1275),
    .ZN(_07075_));
 INV_X1 _32542_ (.A(_07075_),
    .ZN(_07076_));
 NAND2_X1 _32543_ (.A1(_07050_),
    .A2(net1279),
    .ZN(_07077_));
 INV_X8 _32544_ (.A(net1325),
    .ZN(_07078_));
 OR2_X1 _32545_ (.A1(_07078_),
    .A2(\icache.tag_tv_r [131]),
    .ZN(_07079_));
 AND4_X1 _32546_ (.A1(_07073_),
    .A2(_07076_),
    .A3(_07077_),
    .A4(_07079_),
    .ZN(_07080_));
 BUF_X16 _32547_ (.A(_07072_),
    .Z(_07081_));
 NAND2_X1 _32548_ (.A1(_07081_),
    .A2(net1272),
    .ZN(_07082_));
 BUF_X16 _32549_ (.A(_07074_),
    .Z(_07083_));
 NOR2_X1 _32550_ (.A1(_07083_),
    .A2(net1275),
    .ZN(_07084_));
 INV_X1 _32551_ (.A(_07084_),
    .ZN(_07085_));
 BUF_X16 _32552_ (.A(_07078_),
    .Z(_07086_));
 NAND2_X1 _32553_ (.A1(_07086_),
    .A2(\icache.tag_tv_r [131]),
    .ZN(_07087_));
 INV_X8 _32554_ (.A(net1335),
    .ZN(_07088_));
 OR2_X1 _32555_ (.A1(_07088_),
    .A2(net1277),
    .ZN(_07089_));
 AND4_X1 _32556_ (.A1(_07082_),
    .A2(_07085_),
    .A3(_07087_),
    .A4(_07089_),
    .ZN(_07090_));
 AND3_X1 _32557_ (.A1(_07071_),
    .A2(_07080_),
    .A3(_07090_),
    .ZN(_07091_));
 BUF_X16 _32558_ (.A(\icache.addr_tv_r [36]),
    .Z(_07092_));
 XNOR2_X1 _32559_ (.A(_07092_),
    .B(net1273),
    .ZN(_07093_));
 NOR2_X4 _32560_ (.A1(\icache.state_tv_r [9]),
    .A2(\icache.state_tv_r [8]),
    .ZN(_07094_));
 INV_X1 _32561_ (.A(_07094_),
    .ZN(_07095_));
 NOR2_X1 _32562_ (.A1(_07067_),
    .A2(net1300),
    .ZN(_07096_));
 INV_X1 _32563_ (.A(_07096_),
    .ZN(_07097_));
 INV_X1 _32564_ (.A(net1349),
    .ZN(_07098_));
 BUF_X8 _32565_ (.A(_07098_),
    .Z(_07099_));
 OR2_X1 _32566_ (.A1(_07099_),
    .A2(net1283),
    .ZN(_07100_));
 BUF_X16 _32567_ (.A(_07088_),
    .Z(_07101_));
 NAND2_X1 _32568_ (.A1(_07101_),
    .A2(net1277),
    .ZN(_07102_));
 AND4_X1 _32569_ (.A1(_07095_),
    .A2(_07097_),
    .A3(_07100_),
    .A4(_07102_),
    .ZN(_07103_));
 AND4_X1 _32570_ (.A1(_07053_),
    .A2(_07091_),
    .A3(_07093_),
    .A4(_07103_),
    .ZN(_07104_));
 BUF_X16 _32571_ (.A(net1351),
    .Z(_07105_));
 INV_X1 _32572_ (.A(net1288),
    .ZN(_07106_));
 BUF_X16 _32573_ (.A(\icache.addr_tv_r [26]),
    .Z(_07107_));
 INV_X16 _32574_ (.A(_07107_),
    .ZN(_07108_));
 AOI22_X2 _32575_ (.A1(_07105_),
    .A2(_07106_),
    .B1(_07108_),
    .B2(net1285),
    .ZN(_07109_));
 INV_X4 _32576_ (.A(net1344),
    .ZN(_07110_));
 BUF_X16 _32577_ (.A(_07110_),
    .Z(_07111_));
 OAI221_X2 _32578_ (.A(_07109_),
    .B1(_07105_),
    .B2(_07106_),
    .C1(_07111_),
    .C2(net1281),
    .ZN(_07112_));
 BUF_X16 _32579_ (.A(net1366),
    .Z(_07113_));
 INV_X1 _32580_ (.A(net1296),
    .ZN(_07114_));
 AOI22_X2 _32581_ (.A1(_07113_),
    .A2(_07114_),
    .B1(_07111_),
    .B2(net1282),
    .ZN(_07115_));
 INV_X16 _32582_ (.A(\icache.addr_tv_r [34]),
    .ZN(_07116_));
 OAI221_X2 _32583_ (.A(_07115_),
    .B1(_07113_),
    .B2(_07114_),
    .C1(_07116_),
    .C2(net1274),
    .ZN(_07117_));
 BUF_X16 _32584_ (.A(\icache.addr_tv_r [22]),
    .Z(_07118_));
 XNOR2_X2 _32585_ (.A(_07118_),
    .B(net1290),
    .ZN(_07119_));
 INV_X8 _32586_ (.A(net1316),
    .ZN(_07120_));
 NAND2_X1 _32587_ (.A1(_07120_),
    .A2(net1271),
    .ZN(_07121_));
 OAI211_X2 _32588_ (.A(_07119_),
    .B(_07121_),
    .C1(_07108_),
    .C2(net1284),
    .ZN(_07122_));
 BUF_X16 _32589_ (.A(\icache.addr_tv_r [16]),
    .Z(_07123_));
 INV_X1 _32590_ (.A(net1299),
    .ZN(_07124_));
 AOI22_X1 _32591_ (.A1(_07123_),
    .A2(_07124_),
    .B1(_07116_),
    .B2(net1274),
    .ZN(_07125_));
 OAI21_X1 _32592_ (.A(_07125_),
    .B1(_07123_),
    .B2(_07124_),
    .ZN(_07126_));
 NOR4_X2 _32593_ (.A1(_07112_),
    .A2(_07117_),
    .A3(_07122_),
    .A4(_07126_),
    .ZN(_07127_));
 BUF_X16 _32594_ (.A(\icache.addr_tv_r [20]),
    .Z(_07128_));
 XNOR2_X2 _32595_ (.A(_07128_),
    .B(net1292),
    .ZN(_07129_));
 BUF_X16 _32596_ (.A(net1340),
    .Z(_07130_));
 INV_X1 _32597_ (.A(net1278),
    .ZN(_07131_));
 OAI221_X1 _32598_ (.A(_07129_),
    .B1(_07130_),
    .B2(_07131_),
    .C1(_07120_),
    .C2(net1271),
    .ZN(_07132_));
 BUF_X16 _32599_ (.A(\icache.addr_tv_r [32]),
    .Z(_07133_));
 XNOR2_X2 _32600_ (.A(_07133_),
    .B(net1276),
    .ZN(_07134_));
 BUF_X16 _32601_ (.A(\icache.addr_tv_r [25]),
    .Z(_07135_));
 INV_X1 _32602_ (.A(net1286),
    .ZN(_07136_));
 OAI221_X2 _32603_ (.A(_07134_),
    .B1(_07052_),
    .B2(net1298),
    .C1(_07135_),
    .C2(_07136_),
    .ZN(_07137_));
 INV_X8 _32604_ (.A(net1378),
    .ZN(_07138_));
 AOI22_X1 _32605_ (.A1(_07138_),
    .A2(net1301),
    .B1(_07131_),
    .B2(_07130_),
    .ZN(_07139_));
 OAI221_X2 _32606_ (.A(_07139_),
    .B1(_07138_),
    .B2(net1301),
    .C1(_07069_),
    .C2(net1295),
    .ZN(_07140_));
 XNOR2_X2 _32607_ (.A(net1387),
    .B(\icache.tag_tv_r [108]),
    .ZN(_07141_));
 OR2_X1 _32608_ (.A1(_07055_),
    .A2(net1289),
    .ZN(_07142_));
 NAND2_X1 _32609_ (.A1(_07099_),
    .A2(net1283),
    .ZN(_07143_));
 NAND3_X1 _32610_ (.A1(_07141_),
    .A2(_07142_),
    .A3(_07143_),
    .ZN(_07144_));
 NOR4_X1 _32611_ (.A1(_07132_),
    .A2(_07137_),
    .A3(_07140_),
    .A4(_07144_),
    .ZN(_07145_));
 AND3_X4 _32612_ (.A1(_07104_),
    .A2(_07127_),
    .A3(_07145_),
    .ZN(_07146_));
 INV_X1 _32613_ (.A(_07146_),
    .ZN(_07147_));
 INV_X8 _32614_ (.A(\icache.addr_tv_r [16]),
    .ZN(_07148_));
 BUF_X16 _32615_ (.A(_07148_),
    .Z(_07149_));
 NOR2_X1 _32616_ (.A1(_07149_),
    .A2(\icache.tag_tv_r [139]),
    .ZN(_07150_));
 AOI21_X1 _32617_ (.A(_07150_),
    .B1(_07138_),
    .B2(net1268),
    .ZN(_07151_));
 INV_X8 _32618_ (.A(net1343),
    .ZN(_07152_));
 NAND2_X1 _32619_ (.A1(_07152_),
    .A2(\icache.tag_tv_r [153]),
    .ZN(_07153_));
 OAI211_X1 _32620_ (.A(_07151_),
    .B(_07153_),
    .C1(_07138_),
    .C2(net1268),
    .ZN(_07154_));
 XNOR2_X2 _32621_ (.A(_07107_),
    .B(\icache.tag_tv_r [149]),
    .ZN(_07155_));
 BUF_X16 _32622_ (.A(\icache.addr_tv_r [34]),
    .Z(_07156_));
 INV_X1 _32623_ (.A(\icache.tag_tv_r [157]),
    .ZN(_07157_));
 OAI221_X2 _32624_ (.A(_07155_),
    .B1(_07152_),
    .B2(\icache.tag_tv_r [153]),
    .C1(_07156_),
    .C2(_07157_),
    .ZN(_07158_));
 INV_X1 _32625_ (.A(\icache.tag_tv_r [161]),
    .ZN(_07159_));
 BUF_X16 _32626_ (.A(net1314),
    .Z(_07160_));
 AOI22_X1 _32627_ (.A1(_07149_),
    .A2(\icache.tag_tv_r [139]),
    .B1(_07159_),
    .B2(_07160_),
    .ZN(_07161_));
 INV_X16 _32628_ (.A(\icache.addr_tv_r [36]),
    .ZN(_07162_));
 OAI221_X1 _32629_ (.A(_07161_),
    .B1(_07162_),
    .B2(\icache.tag_tv_r [159]),
    .C1(_07160_),
    .C2(_07159_),
    .ZN(_07163_));
 INV_X1 _32630_ (.A(\icache.tag_tv_r [145]),
    .ZN(_07164_));
 AOI22_X1 _32631_ (.A1(_07118_),
    .A2(_07164_),
    .B1(_07162_),
    .B2(\icache.tag_tv_r [159]),
    .ZN(_07165_));
 OAI21_X1 _32632_ (.A(_07165_),
    .B1(_07118_),
    .B2(_07164_),
    .ZN(_07166_));
 OR4_X1 _32633_ (.A1(_07154_),
    .A2(_07158_),
    .A3(_07163_),
    .A4(_07166_),
    .ZN(_07167_));
 BUF_X16 _32634_ (.A(_07059_),
    .Z(_07168_));
 AOI22_X2 _32635_ (.A1(_07168_),
    .A2(\icache.tag_tv_r [144]),
    .B1(_07055_),
    .B2(\icache.tag_tv_r [146]),
    .ZN(_07169_));
 INV_X1 _32636_ (.A(\icache.tag_tv_r [142]),
    .ZN(_07170_));
 OAI221_X2 _32637_ (.A(_07169_),
    .B1(net1364),
    .B2(_07170_),
    .C1(_07168_),
    .C2(\icache.tag_tv_r [144]),
    .ZN(_07171_));
 INV_X16 _32638_ (.A(net1366),
    .ZN(_07172_));
 NOR2_X1 _32639_ (.A1(_07172_),
    .A2(\icache.tag_tv_r [141]),
    .ZN(_07173_));
 AOI21_X1 _32640_ (.A(_07173_),
    .B1(_07111_),
    .B2(\icache.tag_tv_r [151]),
    .ZN(_07174_));
 OR2_X1 _32641_ (.A1(_07078_),
    .A2(\icache.tag_tv_r [158]),
    .ZN(_07175_));
 OAI211_X2 _32642_ (.A(_07174_),
    .B(_07175_),
    .C1(_07111_),
    .C2(\icache.tag_tv_r [151]),
    .ZN(_07176_));
 XNOR2_X2 _32643_ (.A(_07105_),
    .B(\icache.tag_tv_r [147]),
    .ZN(_07177_));
 XNOR2_X2 _32644_ (.A(net1372),
    .B(\icache.tag_tv_r [140]),
    .ZN(_07178_));
 XNOR2_X2 _32645_ (.A(_07128_),
    .B(\icache.tag_tv_r [143]),
    .ZN(_07179_));
 AOI22_X2 _32646_ (.A1(_07172_),
    .A2(\icache.tag_tv_r [141]),
    .B1(_07157_),
    .B2(_07156_),
    .ZN(_07180_));
 NAND4_X2 _32647_ (.A1(_07177_),
    .A2(_07178_),
    .A3(_07179_),
    .A4(_07180_),
    .ZN(_07181_));
 NOR4_X2 _32648_ (.A1(_07167_),
    .A2(_07171_),
    .A3(_07176_),
    .A4(_07181_),
    .ZN(_07182_));
 XNOR2_X1 _32649_ (.A(net1382),
    .B(net1269),
    .ZN(_07183_));
 INV_X8 _32650_ (.A(\icache.addr_tv_r [32]),
    .ZN(_07184_));
 NAND2_X1 _32651_ (.A1(_07184_),
    .A2(\icache.tag_tv_r [155]),
    .ZN(_07185_));
 BUF_X16 _32652_ (.A(net1374),
    .Z(_07186_));
 INV_X1 _32653_ (.A(net1267),
    .ZN(_07187_));
 OAI211_X1 _32654_ (.A(_07183_),
    .B(_07185_),
    .C1(_07186_),
    .C2(_07187_),
    .ZN(_07188_));
 INV_X1 _32655_ (.A(\icache.tag_tv_r [150]),
    .ZN(_07189_));
 BUF_X16 _32656_ (.A(net1350),
    .Z(_07190_));
 OAI22_X2 _32657_ (.A1(_07055_),
    .A2(\icache.tag_tv_r [146]),
    .B1(_07189_),
    .B2(_07190_),
    .ZN(_07191_));
 INV_X1 _32658_ (.A(net1270),
    .ZN(_07192_));
 BUF_X8 _32659_ (.A(net1386),
    .Z(_07193_));
 OAI22_X1 _32660_ (.A1(_07184_),
    .A2(\icache.tag_tv_r [155]),
    .B1(_07192_),
    .B2(_07193_),
    .ZN(_07194_));
 OR3_X1 _32661_ (.A1(_07188_),
    .A2(_07191_),
    .A3(_07194_),
    .ZN(_07195_));
 XOR2_X2 _32662_ (.A(_07135_),
    .B(\icache.tag_tv_r [148]),
    .Z(_07196_));
 NOR2_X1 _32663_ (.A1(_07050_),
    .A2(\icache.tag_tv_r [152]),
    .ZN(_07197_));
 NOR2_X4 _32664_ (.A1(\icache.state_tv_r [11]),
    .A2(\icache.state_tv_r [10]),
    .ZN(_07198_));
 NOR3_X2 _32665_ (.A1(_07196_),
    .A2(_07197_),
    .A3(_07198_),
    .ZN(_07199_));
 NOR2_X1 _32666_ (.A1(_07081_),
    .A2(\icache.tag_tv_r [160]),
    .ZN(_07200_));
 AOI21_X2 _32667_ (.A(_07200_),
    .B1(_07101_),
    .B2(\icache.tag_tv_r [154]),
    .ZN(_07201_));
 NAND2_X1 _32668_ (.A1(_07050_),
    .A2(\icache.tag_tv_r [152]),
    .ZN(_07202_));
 NAND2_X1 _32669_ (.A1(_07189_),
    .A2(_07190_),
    .ZN(_07203_));
 NAND4_X4 _32670_ (.A1(_07199_),
    .A2(_07201_),
    .A3(_07202_),
    .A4(_07203_),
    .ZN(_07204_));
 AOI22_X1 _32671_ (.A1(_07083_),
    .A2(\icache.tag_tv_r [156]),
    .B1(_07192_),
    .B2(_07193_),
    .ZN(_07205_));
 NAND2_X1 _32672_ (.A1(_07086_),
    .A2(\icache.tag_tv_r [158]),
    .ZN(_07206_));
 OAI211_X1 _32673_ (.A(_07205_),
    .B(_07206_),
    .C1(_07069_),
    .C2(\icache.tag_tv_r [142]),
    .ZN(_07207_));
 NOR2_X1 _32674_ (.A1(_07101_),
    .A2(\icache.tag_tv_r [154]),
    .ZN(_07208_));
 AOI21_X1 _32675_ (.A(_07208_),
    .B1(_07081_),
    .B2(\icache.tag_tv_r [160]),
    .ZN(_07209_));
 INV_X1 _32676_ (.A(\icache.tag_tv_r [156]),
    .ZN(_07210_));
 NAND2_X1 _32677_ (.A1(_07210_),
    .A2(net1334),
    .ZN(_07211_));
 OAI211_X1 _32678_ (.A(_07209_),
    .B(_07211_),
    .C1(_07067_),
    .C2(net1267),
    .ZN(_07212_));
 NOR4_X2 _32679_ (.A1(_07195_),
    .A2(_07204_),
    .A3(_07207_),
    .A4(_07212_),
    .ZN(_07213_));
 AND2_X4 _32680_ (.A1(_07182_),
    .A2(_07213_),
    .ZN(_07214_));
 INV_X1 _32681_ (.A(_07214_),
    .ZN(_07215_));
 INV_X1 _32682_ (.A(\icache.tag_tv_r [0]),
    .ZN(_07216_));
 NOR2_X1 _32683_ (.A1(_07216_),
    .A2(net1386),
    .ZN(_07217_));
 INV_X1 _32684_ (.A(_07217_),
    .ZN(_07218_));
 INV_X1 _32685_ (.A(\icache.tag_tv_r [13]),
    .ZN(_07219_));
 NOR2_X1 _32686_ (.A1(_07219_),
    .A2(_07135_),
    .ZN(_07220_));
 INV_X1 _32687_ (.A(_07220_),
    .ZN(_07221_));
 NAND2_X1 _32688_ (.A1(_07168_),
    .A2(\icache.tag_tv_r [9]),
    .ZN(_07222_));
 OR2_X1 _32689_ (.A1(_07068_),
    .A2(\icache.tag_tv_r [7]),
    .ZN(_07223_));
 NAND4_X1 _32690_ (.A1(_07218_),
    .A2(_07221_),
    .A3(_07222_),
    .A4(_07223_),
    .ZN(_07224_));
 XNOR2_X2 _32691_ (.A(net1347),
    .B(\icache.tag_tv_r [16]),
    .ZN(_07225_));
 NAND2_X1 _32692_ (.A1(_07074_),
    .A2(\icache.tag_tv_r [21]),
    .ZN(_07226_));
 OAI211_X2 _32693_ (.A(_07225_),
    .B(_07226_),
    .C1(_07148_),
    .C2(\icache.tag_tv_r [4]),
    .ZN(_07227_));
 OR2_X1 _32694_ (.A1(_07054_),
    .A2(\icache.tag_tv_r [11]),
    .ZN(_07228_));
 OR2_X1 _32695_ (.A1(_07098_),
    .A2(\icache.tag_tv_r [15]),
    .ZN(_07229_));
 OR2_X1 _32696_ (.A1(_07074_),
    .A2(\icache.tag_tv_r [21]),
    .ZN(_07230_));
 NAND2_X1 _32697_ (.A1(_07219_),
    .A2(_07135_),
    .ZN(_07231_));
 NAND4_X1 _32698_ (.A1(_07228_),
    .A2(_07229_),
    .A3(_07230_),
    .A4(_07231_),
    .ZN(_07232_));
 OR2_X1 _32699_ (.A1(_07052_),
    .A2(\icache.tag_tv_r [5]),
    .ZN(_07233_));
 OR2_X1 _32700_ (.A1(_07062_),
    .A2(\icache.tag_tv_r [1]),
    .ZN(_07234_));
 NAND2_X1 _32701_ (.A1(_07099_),
    .A2(\icache.tag_tv_r [15]),
    .ZN(_07235_));
 NAND2_X1 _32702_ (.A1(_07052_),
    .A2(\icache.tag_tv_r [5]),
    .ZN(_07236_));
 NAND4_X1 _32703_ (.A1(_07233_),
    .A2(_07234_),
    .A3(_07235_),
    .A4(_07236_),
    .ZN(_07237_));
 NOR4_X1 _32704_ (.A1(_07224_),
    .A2(_07227_),
    .A3(_07232_),
    .A4(_07237_),
    .ZN(_07238_));
 XNOR2_X1 _32705_ (.A(net1366),
    .B(\icache.tag_tv_r [6]),
    .ZN(_07239_));
 XOR2_X2 _32706_ (.A(net1314),
    .B(\icache.tag_tv_r [26]),
    .Z(_07240_));
 INV_X1 _32707_ (.A(_07240_),
    .ZN(_07241_));
 XNOR2_X1 _32708_ (.A(net1375),
    .B(\icache.tag_tv_r [3]),
    .ZN(_07242_));
 XNOR2_X1 _32709_ (.A(net1376),
    .B(\icache.tag_tv_r [2]),
    .ZN(_07243_));
 AND4_X1 _32710_ (.A1(_07239_),
    .A2(_07241_),
    .A3(_07242_),
    .A4(_07243_),
    .ZN(_07244_));
 AND2_X2 _32711_ (.A1(_07238_),
    .A2(_07244_),
    .ZN(_07245_));
 INV_X1 _32712_ (.A(\icache.tag_tv_r [19]),
    .ZN(_07246_));
 NOR2_X1 _32713_ (.A1(_07246_),
    .A2(net1335),
    .ZN(_07247_));
 BUF_X16 _32714_ (.A(\icache.addr_tv_r [29]),
    .Z(_07248_));
 INV_X1 _32715_ (.A(\icache.tag_tv_r [17]),
    .ZN(_07249_));
 AOI21_X1 _32716_ (.A(_07247_),
    .B1(_07248_),
    .B2(_07249_),
    .ZN(_07250_));
 OAI221_X2 _32717_ (.A(_07250_),
    .B1(_07184_),
    .B2(\icache.tag_tv_r [20]),
    .C1(_07081_),
    .C2(\icache.tag_tv_r [25]),
    .ZN(_07251_));
 OR2_X1 _32718_ (.A1(_07168_),
    .A2(\icache.tag_tv_r [9]),
    .ZN(_07252_));
 INV_X4 _32719_ (.A(\icache.addr_tv_r [20]),
    .ZN(_07253_));
 NAND2_X1 _32720_ (.A1(_07253_),
    .A2(\icache.tag_tv_r [8]),
    .ZN(_07254_));
 NOR2_X4 _32721_ (.A1(\icache.state_tv_r [1]),
    .A2(\icache.state_tv_r [0]),
    .ZN(_07255_));
 INV_X1 _32722_ (.A(_07255_),
    .ZN(_07256_));
 NAND2_X1 _32723_ (.A1(_07055_),
    .A2(\icache.tag_tv_r [11]),
    .ZN(_07257_));
 NAND4_X2 _32724_ (.A1(_07252_),
    .A2(_07254_),
    .A3(_07256_),
    .A4(_07257_),
    .ZN(_07258_));
 AOI22_X2 _32725_ (.A1(_07148_),
    .A2(\icache.tag_tv_r [4]),
    .B1(_07184_),
    .B2(\icache.tag_tv_r [20]),
    .ZN(_07259_));
 NAND2_X1 _32726_ (.A1(_07162_),
    .A2(\icache.tag_tv_r [24]),
    .ZN(_07260_));
 OAI211_X2 _32727_ (.A(_07259_),
    .B(_07260_),
    .C1(_07116_),
    .C2(\icache.tag_tv_r [22]),
    .ZN(_07261_));
 OR2_X1 _32728_ (.A1(_07078_),
    .A2(\icache.tag_tv_r [23]),
    .ZN(_07262_));
 NAND2_X1 _32729_ (.A1(_07086_),
    .A2(\icache.tag_tv_r [23]),
    .ZN(_07263_));
 OAI211_X2 _32730_ (.A(_07262_),
    .B(_07263_),
    .C1(_07101_),
    .C2(\icache.tag_tv_r [19]),
    .ZN(_07264_));
 NOR4_X2 _32731_ (.A1(_07251_),
    .A2(_07258_),
    .A3(_07261_),
    .A4(_07264_),
    .ZN(_07265_));
 AOI22_X1 _32732_ (.A1(_07116_),
    .A2(\icache.tag_tv_r [22]),
    .B1(_07216_),
    .B2(_07193_),
    .ZN(_07266_));
 XNOR2_X2 _32733_ (.A(net1341),
    .B(\icache.tag_tv_r [18]),
    .ZN(_07267_));
 OR2_X1 _32734_ (.A1(_07253_),
    .A2(\icache.tag_tv_r [8]),
    .ZN(_07268_));
 OAI211_X1 _32735_ (.A(_07267_),
    .B(_07268_),
    .C1(_07162_),
    .C2(\icache.tag_tv_r [24]),
    .ZN(_07269_));
 XNOR2_X2 _32736_ (.A(_07107_),
    .B(\icache.tag_tv_r [14]),
    .ZN(_07270_));
 XNOR2_X1 _32737_ (.A(net1352),
    .B(\icache.tag_tv_r [12]),
    .ZN(_07271_));
 NAND2_X1 _32738_ (.A1(_07270_),
    .A2(_07271_),
    .ZN(_07272_));
 NOR2_X1 _32739_ (.A1(_07269_),
    .A2(_07272_),
    .ZN(_07273_));
 XNOR2_X1 _32740_ (.A(_07118_),
    .B(\icache.tag_tv_r [10]),
    .ZN(_07274_));
 NAND2_X1 _32741_ (.A1(_07050_),
    .A2(\icache.tag_tv_r [17]),
    .ZN(_07275_));
 INV_X1 _32742_ (.A(\icache.tag_tv_r [25]),
    .ZN(_07276_));
 NOR2_X1 _32743_ (.A1(_07276_),
    .A2(net1322),
    .ZN(_07277_));
 INV_X1 _32744_ (.A(_07277_),
    .ZN(_07278_));
 NAND2_X1 _32745_ (.A1(_07062_),
    .A2(\icache.tag_tv_r [1]),
    .ZN(_07279_));
 NAND2_X1 _32746_ (.A1(_07068_),
    .A2(\icache.tag_tv_r [7]),
    .ZN(_07280_));
 AND4_X1 _32747_ (.A1(_07275_),
    .A2(_07278_),
    .A3(_07279_),
    .A4(_07280_),
    .ZN(_07281_));
 AND4_X1 _32748_ (.A1(_07266_),
    .A2(_07273_),
    .A3(_07274_),
    .A4(_07281_),
    .ZN(_07282_));
 AND3_X4 _32749_ (.A1(_07245_),
    .A2(_07265_),
    .A3(_07282_),
    .ZN(_07283_));
 NAND2_X1 _32750_ (.A1(_07088_),
    .A2(\icache.tag_tv_r [46]),
    .ZN(_07284_));
 INV_X4 _32751_ (.A(net1385),
    .ZN(_07285_));
 OR2_X1 _32752_ (.A1(_07285_),
    .A2(\icache.tag_tv_r [27]),
    .ZN(_07286_));
 AND2_X1 _32753_ (.A1(_07284_),
    .A2(_07286_),
    .ZN(_07287_));
 INV_X1 _32754_ (.A(\icache.tag_tv_r [33]),
    .ZN(_07288_));
 OAI221_X1 _32755_ (.A(_07287_),
    .B1(_07113_),
    .B2(_07288_),
    .C1(_07101_),
    .C2(\icache.tag_tv_r [46]),
    .ZN(_07289_));
 INV_X1 _32756_ (.A(\icache.tag_tv_r [35]),
    .ZN(_07290_));
 AOI22_X1 _32757_ (.A1(_07148_),
    .A2(\icache.tag_tv_r [31]),
    .B1(_07290_),
    .B2(_07128_),
    .ZN(_07291_));
 NAND2_X1 _32758_ (.A1(_07067_),
    .A2(\icache.tag_tv_r [30]),
    .ZN(_07292_));
 OAI211_X1 _32759_ (.A(_07291_),
    .B(_07292_),
    .C1(_07149_),
    .C2(\icache.tag_tv_r [31]),
    .ZN(_07293_));
 NAND2_X1 _32760_ (.A1(_07052_),
    .A2(\icache.tag_tv_r [32]),
    .ZN(_07294_));
 OR2_X1 _32761_ (.A1(_07052_),
    .A2(\icache.tag_tv_r [32]),
    .ZN(_07295_));
 OAI211_X1 _32762_ (.A(_07294_),
    .B(_07295_),
    .C1(_07172_),
    .C2(\icache.tag_tv_r [33]),
    .ZN(_07296_));
 XNOR2_X2 _32763_ (.A(_07105_),
    .B(\icache.tag_tv_r [39]),
    .ZN(_07297_));
 OR2_X1 _32764_ (.A1(_07057_),
    .A2(\icache.tag_tv_r [40]),
    .ZN(_07298_));
 OAI211_X1 _32765_ (.A(_07297_),
    .B(_07298_),
    .C1(_07128_),
    .C2(_07290_),
    .ZN(_07299_));
 NOR4_X1 _32766_ (.A1(_07289_),
    .A2(_07293_),
    .A3(_07296_),
    .A4(_07299_),
    .ZN(_07300_));
 XNOR2_X1 _32767_ (.A(net1345),
    .B(\icache.tag_tv_r [43]),
    .ZN(_07301_));
 XOR2_X1 _32768_ (.A(\icache.addr_tv_r [26]),
    .B(\icache.tag_tv_r [41]),
    .Z(_07302_));
 INV_X1 _32769_ (.A(_07302_),
    .ZN(_07303_));
 XNOR2_X1 _32770_ (.A(net1339),
    .B(\icache.tag_tv_r [45]),
    .ZN(_07304_));
 XNOR2_X1 _32771_ (.A(_07248_),
    .B(\icache.tag_tv_r [44]),
    .ZN(_07305_));
 AND4_X1 _32772_ (.A1(_07301_),
    .A2(_07303_),
    .A3(_07304_),
    .A4(_07305_),
    .ZN(_07306_));
 XNOR2_X1 _32773_ (.A(_07133_),
    .B(\icache.tag_tv_r [47]),
    .ZN(_07307_));
 XOR2_X2 _32774_ (.A(\icache.addr_tv_r [22]),
    .B(\icache.tag_tv_r [37]),
    .Z(_07308_));
 INV_X1 _32775_ (.A(_07308_),
    .ZN(_07309_));
 XNOR2_X2 _32776_ (.A(\icache.addr_tv_r [34]),
    .B(\icache.tag_tv_r [49]),
    .ZN(_07310_));
 XNOR2_X2 _32777_ (.A(\icache.addr_tv_r [36]),
    .B(\icache.tag_tv_r [51]),
    .ZN(_07311_));
 AND4_X1 _32778_ (.A1(_07307_),
    .A2(_07309_),
    .A3(_07310_),
    .A4(_07311_),
    .ZN(_07312_));
 XNOR2_X2 _32779_ (.A(net1332),
    .B(\icache.tag_tv_r [48]),
    .ZN(_07313_));
 XNOR2_X2 _32780_ (.A(net1318),
    .B(\icache.tag_tv_r [52]),
    .ZN(_07314_));
 NAND2_X1 _32781_ (.A1(_07313_),
    .A2(_07314_),
    .ZN(_07315_));
 INV_X1 _32782_ (.A(\icache.tag_tv_r [50]),
    .ZN(_07316_));
 OAI22_X1 _32783_ (.A1(_07138_),
    .A2(\icache.tag_tv_r [29]),
    .B1(_07316_),
    .B2(net1325),
    .ZN(_07317_));
 AND2_X1 _32784_ (.A1(_07138_),
    .A2(\icache.tag_tv_r [29]),
    .ZN(_07318_));
 NOR2_X1 _32785_ (.A1(_07065_),
    .A2(\icache.tag_tv_r [28]),
    .ZN(_07319_));
 NOR4_X1 _32786_ (.A1(_07315_),
    .A2(_07317_),
    .A3(_07318_),
    .A4(_07319_),
    .ZN(_07320_));
 AND3_X1 _32787_ (.A1(_07306_),
    .A2(_07312_),
    .A3(_07320_),
    .ZN(_07321_));
 OR2_X1 _32788_ (.A1(_07099_),
    .A2(\icache.tag_tv_r [42]),
    .ZN(_07322_));
 OR2_X1 _32789_ (.A1(_07068_),
    .A2(\icache.tag_tv_r [34]),
    .ZN(_07323_));
 NAND2_X1 _32790_ (.A1(_07068_),
    .A2(\icache.tag_tv_r [34]),
    .ZN(_07324_));
 INV_X1 _32791_ (.A(\icache.tag_tv_r [53]),
    .ZN(_07325_));
 NAND2_X1 _32792_ (.A1(_07325_),
    .A2(_07160_),
    .ZN(_07326_));
 AND4_X1 _32793_ (.A1(_07322_),
    .A2(_07323_),
    .A3(_07324_),
    .A4(_07326_),
    .ZN(_07327_));
 OAI22_X1 _32794_ (.A1(_07054_),
    .A2(\icache.tag_tv_r [38]),
    .B1(_07078_),
    .B2(\icache.tag_tv_r [50]),
    .ZN(_07328_));
 AOI221_X4 _32795_ (.A(_07328_),
    .B1(_07099_),
    .B2(\icache.tag_tv_r [42]),
    .C1(_07120_),
    .C2(\icache.tag_tv_r [53]),
    .ZN(_07329_));
 NAND2_X1 _32796_ (.A1(_07065_),
    .A2(\icache.tag_tv_r [28]),
    .ZN(_07330_));
 OR2_X1 _32797_ (.A1(_07059_),
    .A2(\icache.tag_tv_r [36]),
    .ZN(_07331_));
 NAND2_X1 _32798_ (.A1(_07057_),
    .A2(\icache.tag_tv_r [40]),
    .ZN(_07332_));
 NOR2_X4 _32799_ (.A1(\icache.state_tv_r [3]),
    .A2(\icache.state_tv_r [2]),
    .ZN(_07333_));
 INV_X1 _32800_ (.A(_07333_),
    .ZN(_07334_));
 AND4_X1 _32801_ (.A1(_07330_),
    .A2(_07331_),
    .A3(_07332_),
    .A4(_07334_),
    .ZN(_07335_));
 NAND2_X1 _32802_ (.A1(_07055_),
    .A2(\icache.tag_tv_r [38]),
    .ZN(_07336_));
 OR2_X1 _32803_ (.A1(_07067_),
    .A2(\icache.tag_tv_r [30]),
    .ZN(_07337_));
 NAND2_X1 _32804_ (.A1(_07168_),
    .A2(\icache.tag_tv_r [36]),
    .ZN(_07338_));
 NAND2_X1 _32805_ (.A1(_07285_),
    .A2(\icache.tag_tv_r [27]),
    .ZN(_07339_));
 AND4_X1 _32806_ (.A1(_07336_),
    .A2(_07337_),
    .A3(_07338_),
    .A4(_07339_),
    .ZN(_07340_));
 AND4_X1 _32807_ (.A1(_07327_),
    .A2(_07329_),
    .A3(_07335_),
    .A4(_07340_),
    .ZN(_07341_));
 AND3_X4 _32808_ (.A1(_07300_),
    .A2(_07321_),
    .A3(_07341_),
    .ZN(_07342_));
 NOR2_X2 _32809_ (.A1(_07283_),
    .A2(_07342_),
    .ZN(_07343_));
 XNOR2_X1 _32810_ (.A(_07105_),
    .B(\icache.tag_tv_r [93]),
    .ZN(_07344_));
 XNOR2_X1 _32811_ (.A(net1315),
    .B(\icache.tag_tv_r [107]),
    .ZN(_07345_));
 XNOR2_X1 _32812_ (.A(_07133_),
    .B(\icache.tag_tv_r [101]),
    .ZN(_07346_));
 XNOR2_X2 _32813_ (.A(_07128_),
    .B(\icache.tag_tv_r [89]),
    .ZN(_07347_));
 AND4_X1 _32814_ (.A1(_07344_),
    .A2(_07345_),
    .A3(_07346_),
    .A4(_07347_),
    .ZN(_07348_));
 NOR2_X1 _32815_ (.A1(_07111_),
    .A2(\icache.tag_tv_r [97]),
    .ZN(_07349_));
 NOR2_X4 _32816_ (.A1(\icache.state_tv_r [7]),
    .A2(\icache.state_tv_r [6]),
    .ZN(_07350_));
 INV_X8 _32817_ (.A(_07350_),
    .ZN(_07351_));
 OAI21_X1 _32818_ (.A(_07351_),
    .B1(_07072_),
    .B2(\icache.tag_tv_r [106]),
    .ZN(_07352_));
 AOI211_X1 _32819_ (.A(_07349_),
    .B(_07352_),
    .C1(_07152_),
    .C2(\icache.tag_tv_r [99]),
    .ZN(_07353_));
 INV_X1 _32820_ (.A(\icache.tag_tv_r [99]),
    .ZN(_07354_));
 AOI22_X1 _32821_ (.A1(_07130_),
    .A2(_07354_),
    .B1(_07083_),
    .B2(\icache.tag_tv_r [102]),
    .ZN(_07355_));
 XNOR2_X1 _32822_ (.A(net1327),
    .B(\icache.tag_tv_r [104]),
    .ZN(_07356_));
 XNOR2_X2 _32823_ (.A(_07118_),
    .B(\icache.tag_tv_r [91]),
    .ZN(_07357_));
 XNOR2_X1 _32824_ (.A(_07156_),
    .B(\icache.tag_tv_r [103]),
    .ZN(_07358_));
 AND4_X1 _32825_ (.A1(_07355_),
    .A2(_07356_),
    .A3(_07357_),
    .A4(_07358_),
    .ZN(_07359_));
 NAND2_X1 _32826_ (.A1(_07110_),
    .A2(\icache.tag_tv_r [97]),
    .ZN(_07360_));
 OAI21_X1 _32827_ (.A(_07360_),
    .B1(_07162_),
    .B2(\icache.tag_tv_r [105]),
    .ZN(_07361_));
 INV_X1 _32828_ (.A(\icache.tag_tv_r [95]),
    .ZN(_07362_));
 AOI221_X4 _32829_ (.A(_07361_),
    .B1(_07107_),
    .B2(_07362_),
    .C1(_07162_),
    .C2(\icache.tag_tv_r [105]),
    .ZN(_07363_));
 AND4_X1 _32830_ (.A1(_07348_),
    .A2(_07353_),
    .A3(_07359_),
    .A4(_07363_),
    .ZN(_07364_));
 NOR2_X1 _32831_ (.A1(_07149_),
    .A2(\icache.tag_tv_r [85]),
    .ZN(_07365_));
 AND2_X1 _32832_ (.A1(_07052_),
    .A2(\icache.tag_tv_r [86]),
    .ZN(_07366_));
 NOR2_X1 _32833_ (.A1(_07067_),
    .A2(\icache.tag_tv_r [84]),
    .ZN(_07367_));
 NOR2_X1 _32834_ (.A1(_07052_),
    .A2(\icache.tag_tv_r [86]),
    .ZN(_07368_));
 OR4_X1 _32835_ (.A1(_07365_),
    .A2(_07366_),
    .A3(_07367_),
    .A4(_07368_),
    .ZN(_07369_));
 BUF_X16 _32836_ (.A(net1376),
    .Z(_07370_));
 INV_X1 _32837_ (.A(\icache.tag_tv_r [83]),
    .ZN(_07371_));
 AOI22_X1 _32838_ (.A1(_07370_),
    .A2(_07371_),
    .B1(_07172_),
    .B2(\icache.tag_tv_r [87]),
    .ZN(_07372_));
 OAI221_X1 _32839_ (.A(_07372_),
    .B1(_07172_),
    .B2(\icache.tag_tv_r [87]),
    .C1(_07107_),
    .C2(_07362_),
    .ZN(_07373_));
 AOI22_X1 _32840_ (.A1(_07065_),
    .A2(\icache.tag_tv_r [82]),
    .B1(_07149_),
    .B2(\icache.tag_tv_r [85]),
    .ZN(_07374_));
 OR2_X1 _32841_ (.A1(_07285_),
    .A2(\icache.tag_tv_r [81]),
    .ZN(_07375_));
 OAI211_X1 _32842_ (.A(_07374_),
    .B(_07375_),
    .C1(_07370_),
    .C2(_07371_),
    .ZN(_07376_));
 NOR2_X1 _32843_ (.A1(_07099_),
    .A2(\icache.tag_tv_r [96]),
    .ZN(_07377_));
 INV_X1 _32844_ (.A(_07377_),
    .ZN(_07378_));
 OR2_X1 _32845_ (.A1(_07055_),
    .A2(\icache.tag_tv_r [92]),
    .ZN(_07379_));
 OR2_X2 _32846_ (.A1(_07050_),
    .A2(\icache.tag_tv_r [98]),
    .ZN(_07380_));
 NAND2_X1 _32847_ (.A1(_07285_),
    .A2(\icache.tag_tv_r [81]),
    .ZN(_07381_));
 NAND4_X1 _32848_ (.A1(_07378_),
    .A2(_07379_),
    .A3(_07380_),
    .A4(_07381_),
    .ZN(_07382_));
 NOR4_X1 _32849_ (.A1(_07369_),
    .A2(_07373_),
    .A3(_07376_),
    .A4(_07382_),
    .ZN(_07383_));
 NOR2_X1 _32850_ (.A1(_07065_),
    .A2(\icache.tag_tv_r [82]),
    .ZN(_07384_));
 AOI21_X1 _32851_ (.A(_07384_),
    .B1(_07168_),
    .B2(\icache.tag_tv_r [90]),
    .ZN(_07385_));
 OR2_X1 _32852_ (.A1(_07069_),
    .A2(\icache.tag_tv_r [88]),
    .ZN(_07386_));
 INV_X1 _32853_ (.A(\icache.tag_tv_r [96]),
    .ZN(_07387_));
 OAI211_X1 _32854_ (.A(_07385_),
    .B(_07386_),
    .C1(_07190_),
    .C2(_07387_),
    .ZN(_07388_));
 INV_X1 _32855_ (.A(\icache.tag_tv_r [84]),
    .ZN(_07389_));
 NOR2_X1 _32856_ (.A1(_07389_),
    .A2(_07186_),
    .ZN(_07390_));
 INV_X1 _32857_ (.A(_07390_),
    .ZN(_07391_));
 NAND2_X1 _32858_ (.A1(_07069_),
    .A2(\icache.tag_tv_r [88]),
    .ZN(_07392_));
 NAND2_X1 _32859_ (.A1(_07101_),
    .A2(\icache.tag_tv_r [100]),
    .ZN(_07393_));
 NAND2_X1 _32860_ (.A1(_07055_),
    .A2(\icache.tag_tv_r [92]),
    .ZN(_07394_));
 NAND4_X1 _32861_ (.A1(_07391_),
    .A2(_07392_),
    .A3(_07393_),
    .A4(_07394_),
    .ZN(_07395_));
 AOI22_X1 _32862_ (.A1(_07057_),
    .A2(\icache.tag_tv_r [94]),
    .B1(_07081_),
    .B2(\icache.tag_tv_r [106]),
    .ZN(_07396_));
 OR2_X1 _32863_ (.A1(_07057_),
    .A2(\icache.tag_tv_r [94]),
    .ZN(_07397_));
 OAI211_X1 _32864_ (.A(_07396_),
    .B(_07397_),
    .C1(_07168_),
    .C2(\icache.tag_tv_r [90]),
    .ZN(_07398_));
 NAND2_X1 _32865_ (.A1(_07050_),
    .A2(\icache.tag_tv_r [98]),
    .ZN(_07399_));
 OAI221_X2 _32866_ (.A(_07399_),
    .B1(_07101_),
    .B2(\icache.tag_tv_r [100]),
    .C1(_07083_),
    .C2(\icache.tag_tv_r [102]),
    .ZN(_07400_));
 NOR4_X1 _32867_ (.A1(_07388_),
    .A2(_07395_),
    .A3(_07398_),
    .A4(_07400_),
    .ZN(_07401_));
 AND3_X4 _32868_ (.A1(_07364_),
    .A2(_07383_),
    .A3(_07401_),
    .ZN(_07402_));
 INV_X1 _32869_ (.A(_07402_),
    .ZN(_07403_));
 XNOR2_X2 _32870_ (.A(net1315),
    .B(\icache.tag_tv_r [80]),
    .ZN(_07404_));
 XOR2_X1 _32871_ (.A(_07128_),
    .B(\icache.tag_tv_r [62]),
    .Z(_07405_));
 INV_X1 _32872_ (.A(_07405_),
    .ZN(_07406_));
 AOI22_X1 _32873_ (.A1(_07108_),
    .A2(\icache.tag_tv_r [68]),
    .B1(_07162_),
    .B2(\icache.tag_tv_r [78]),
    .ZN(_07407_));
 XNOR2_X2 _32874_ (.A(\icache.addr_tv_r [22]),
    .B(\icache.tag_tv_r [64]),
    .ZN(_07408_));
 AND4_X1 _32875_ (.A1(_07404_),
    .A2(_07406_),
    .A3(_07407_),
    .A4(_07408_),
    .ZN(_07409_));
 NOR2_X1 _32876_ (.A1(_07116_),
    .A2(\icache.tag_tv_r [76]),
    .ZN(_07410_));
 AOI21_X1 _32877_ (.A(_07410_),
    .B1(_07152_),
    .B2(\icache.tag_tv_r [72]),
    .ZN(_07411_));
 NOR2_X1 _32878_ (.A1(_07110_),
    .A2(\icache.tag_tv_r [70]),
    .ZN(_07412_));
 INV_X1 _32879_ (.A(\icache.tag_tv_r [60]),
    .ZN(_07413_));
 AOI21_X1 _32880_ (.A(_07412_),
    .B1(net1367),
    .B2(_07413_),
    .ZN(_07414_));
 NOR2_X1 _32881_ (.A1(_07152_),
    .A2(\icache.tag_tv_r [72]),
    .ZN(_07415_));
 AOI21_X1 _32882_ (.A(_07415_),
    .B1(_07110_),
    .B2(\icache.tag_tv_r [70]),
    .ZN(_07416_));
 AOI22_X1 _32883_ (.A1(_07083_),
    .A2(\icache.tag_tv_r [75]),
    .B1(_07116_),
    .B2(\icache.tag_tv_r [76]),
    .ZN(_07417_));
 AND4_X1 _32884_ (.A1(_07411_),
    .A2(_07414_),
    .A3(_07416_),
    .A4(_07417_),
    .ZN(_07418_));
 NOR2_X1 _32885_ (.A1(_07168_),
    .A2(\icache.tag_tv_r [63]),
    .ZN(_07419_));
 AND2_X1 _32886_ (.A1(_07049_),
    .A2(\icache.tag_tv_r [71]),
    .ZN(_07420_));
 NOR2_X1 _32887_ (.A1(_07099_),
    .A2(\icache.tag_tv_r [69]),
    .ZN(_07421_));
 NOR2_X1 _32888_ (.A1(_07086_),
    .A2(\icache.tag_tv_r [77]),
    .ZN(_07422_));
 NOR4_X1 _32889_ (.A1(_07419_),
    .A2(_07420_),
    .A3(_07421_),
    .A4(_07422_),
    .ZN(_07423_));
 OAI22_X1 _32890_ (.A1(_07083_),
    .A2(\icache.tag_tv_r [75]),
    .B1(_07081_),
    .B2(\icache.tag_tv_r [79]),
    .ZN(_07424_));
 NOR2_X4 _32891_ (.A1(\icache.state_tv_r [5]),
    .A2(\icache.state_tv_r [4]),
    .ZN(_07425_));
 NOR2_X1 _32892_ (.A1(_07050_),
    .A2(\icache.tag_tv_r [71]),
    .ZN(_07426_));
 NOR3_X1 _32893_ (.A1(_07424_),
    .A2(_07425_),
    .A3(_07426_),
    .ZN(_07427_));
 AND4_X1 _32894_ (.A1(_07409_),
    .A2(_07418_),
    .A3(_07423_),
    .A4(_07427_),
    .ZN(_07428_));
 XNOR2_X2 _32895_ (.A(_07105_),
    .B(\icache.tag_tv_r [66]),
    .ZN(_07429_));
 OAI221_X2 _32896_ (.A(_07429_),
    .B1(_07113_),
    .B2(_07413_),
    .C1(_07108_),
    .C2(\icache.tag_tv_r [68]),
    .ZN(_07430_));
 AOI22_X2 _32897_ (.A1(_07138_),
    .A2(\icache.tag_tv_r [56]),
    .B1(_07055_),
    .B2(\icache.tag_tv_r [65]),
    .ZN(_07431_));
 OAI221_X2 _32898_ (.A(_07431_),
    .B1(_07138_),
    .B2(\icache.tag_tv_r [56]),
    .C1(_07162_),
    .C2(\icache.tag_tv_r [78]),
    .ZN(_07432_));
 OR2_X1 _32899_ (.A1(_07065_),
    .A2(\icache.tag_tv_r [55]),
    .ZN(_07433_));
 INV_X1 _32900_ (.A(\icache.tag_tv_r [57]),
    .ZN(_07434_));
 INV_X1 _32901_ (.A(\icache.tag_tv_r [63]),
    .ZN(_07435_));
 OAI221_X2 _32902_ (.A(_07433_),
    .B1(_07186_),
    .B2(_07434_),
    .C1(net1356),
    .C2(_07435_),
    .ZN(_07436_));
 XNOR2_X1 _32903_ (.A(net1370),
    .B(\icache.tag_tv_r [59]),
    .ZN(_07437_));
 AOI22_X1 _32904_ (.A1(_07149_),
    .A2(\icache.tag_tv_r [58]),
    .B1(_07184_),
    .B2(\icache.tag_tv_r [74]),
    .ZN(_07438_));
 NAND2_X1 _32905_ (.A1(_07437_),
    .A2(_07438_),
    .ZN(_07439_));
 NOR4_X1 _32906_ (.A1(_07430_),
    .A2(_07432_),
    .A3(_07436_),
    .A4(_07439_),
    .ZN(_07440_));
 OR2_X1 _32907_ (.A1(_07088_),
    .A2(\icache.tag_tv_r [73]),
    .ZN(_07441_));
 NAND2_X1 _32908_ (.A1(_07086_),
    .A2(\icache.tag_tv_r [77]),
    .ZN(_07442_));
 AND2_X1 _32909_ (.A1(_07441_),
    .A2(_07442_),
    .ZN(_07443_));
 OR2_X1 _32910_ (.A1(_07057_),
    .A2(\icache.tag_tv_r [67]),
    .ZN(_07444_));
 OAI211_X2 _32911_ (.A(_07443_),
    .B(_07444_),
    .C1(_07069_),
    .C2(\icache.tag_tv_r [61]),
    .ZN(_07445_));
 INV_X1 _32912_ (.A(\icache.tag_tv_r [54]),
    .ZN(_07446_));
 AOI22_X2 _32913_ (.A1(_07186_),
    .A2(_07434_),
    .B1(_07446_),
    .B2(_07193_),
    .ZN(_07447_));
 OAI221_X2 _32914_ (.A(_07447_),
    .B1(_07149_),
    .B2(\icache.tag_tv_r [58]),
    .C1(_07184_),
    .C2(\icache.tag_tv_r [74]),
    .ZN(_07448_));
 OR2_X1 _32915_ (.A1(_07055_),
    .A2(\icache.tag_tv_r [65]),
    .ZN(_07449_));
 NAND2_X1 _32916_ (.A1(_07065_),
    .A2(\icache.tag_tv_r [55]),
    .ZN(_07450_));
 NAND2_X2 _32917_ (.A1(_07101_),
    .A2(\icache.tag_tv_r [73]),
    .ZN(_07451_));
 NAND2_X1 _32918_ (.A1(_07285_),
    .A2(\icache.tag_tv_r [54]),
    .ZN(_07452_));
 NAND4_X1 _32919_ (.A1(_07449_),
    .A2(_07450_),
    .A3(_07451_),
    .A4(_07452_),
    .ZN(_07453_));
 AOI22_X1 _32920_ (.A1(_07069_),
    .A2(\icache.tag_tv_r [61]),
    .B1(_07072_),
    .B2(\icache.tag_tv_r [79]),
    .ZN(_07454_));
 NAND2_X1 _32921_ (.A1(_07057_),
    .A2(\icache.tag_tv_r [67]),
    .ZN(_07455_));
 INV_X1 _32922_ (.A(\icache.tag_tv_r [69]),
    .ZN(_07456_));
 OAI211_X1 _32923_ (.A(_07454_),
    .B(_07455_),
    .C1(_07190_),
    .C2(_07456_),
    .ZN(_07457_));
 NOR4_X1 _32924_ (.A1(_07445_),
    .A2(_07448_),
    .A3(_07453_),
    .A4(_07457_),
    .ZN(_07458_));
 AND3_X4 _32925_ (.A1(_07428_),
    .A2(_07440_),
    .A3(_07458_),
    .ZN(_07459_));
 INV_X2 _32926_ (.A(_07459_),
    .ZN(_07460_));
 AND3_X2 _32927_ (.A1(_07343_),
    .A2(_07403_),
    .A3(_07460_),
    .ZN(_07461_));
 AND3_X1 _32928_ (.A1(_07147_),
    .A2(_07215_),
    .A3(_07461_),
    .ZN(_07462_));
 XNOR2_X1 _32929_ (.A(_07160_),
    .B(\icache.tag_tv_r [188]),
    .ZN(_07463_));
 XOR2_X1 _32930_ (.A(net1352),
    .B(\icache.tag_tv_r [174]),
    .Z(_07464_));
 INV_X1 _32931_ (.A(_07464_),
    .ZN(_07465_));
 XNOR2_X2 _32932_ (.A(_07133_),
    .B(\icache.tag_tv_r [182]),
    .ZN(_07466_));
 XNOR2_X1 _32933_ (.A(net1372),
    .B(\icache.tag_tv_r [167]),
    .ZN(_07467_));
 AND4_X1 _32934_ (.A1(_07463_),
    .A2(_07465_),
    .A3(_07466_),
    .A4(_07467_),
    .ZN(_07468_));
 XNOR2_X1 _32935_ (.A(net1363),
    .B(\icache.tag_tv_r [169]),
    .ZN(_07469_));
 OR2_X1 _32936_ (.A1(_07108_),
    .A2(\icache.tag_tv_r [176]),
    .ZN(_07470_));
 NAND2_X1 _32937_ (.A1(_07172_),
    .A2(\icache.tag_tv_r [168]),
    .ZN(_07471_));
 AND3_X1 _32938_ (.A1(_07469_),
    .A2(_07470_),
    .A3(_07471_),
    .ZN(_07472_));
 XNOR2_X1 _32939_ (.A(net1355),
    .B(\icache.tag_tv_r [173]),
    .ZN(_07473_));
 XNOR2_X2 _32940_ (.A(net1338),
    .B(\icache.tag_tv_r [181]),
    .ZN(_07474_));
 AND4_X1 _32941_ (.A1(_07468_),
    .A2(_07472_),
    .A3(_07473_),
    .A4(_07474_),
    .ZN(_07475_));
 XNOR2_X1 _32942_ (.A(\icache.tag_tv_r [162]),
    .B(net1388),
    .ZN(_07476_));
 XNOR2_X2 _32943_ (.A(_07092_),
    .B(\icache.tag_tv_r [186]),
    .ZN(_07477_));
 XOR2_X1 _32944_ (.A(net1379),
    .B(\icache.tag_tv_r [164]),
    .Z(_07478_));
 XOR2_X1 _32945_ (.A(net1374),
    .B(\icache.tag_tv_r [165]),
    .Z(_07479_));
 NOR2_X1 _32946_ (.A1(_07478_),
    .A2(_07479_),
    .ZN(_07480_));
 NAND4_X2 _32947_ (.A1(_07475_),
    .A2(_07476_),
    .A3(_07477_),
    .A4(_07480_),
    .ZN(_07481_));
 XNOR2_X2 _32948_ (.A(_07190_),
    .B(\icache.tag_tv_r [177]),
    .ZN(_07482_));
 INV_X1 _32949_ (.A(\icache.tag_tv_r [179]),
    .ZN(_07483_));
 OAI221_X2 _32950_ (.A(_07482_),
    .B1(_07248_),
    .B2(_07483_),
    .C1(_07086_),
    .C2(\icache.tag_tv_r [185]),
    .ZN(_07484_));
 XNOR2_X1 _32951_ (.A(net1360),
    .B(\icache.tag_tv_r [171]),
    .ZN(_07485_));
 INV_X1 _32952_ (.A(_07118_),
    .ZN(_07486_));
 NAND2_X1 _32953_ (.A1(_07486_),
    .A2(\icache.tag_tv_r [172]),
    .ZN(_07487_));
 OAI211_X2 _32954_ (.A(_07485_),
    .B(_07487_),
    .C1(_07081_),
    .C2(\icache.tag_tv_r [187]),
    .ZN(_07488_));
 XNOR2_X2 _32955_ (.A(_07156_),
    .B(\icache.tag_tv_r [184]),
    .ZN(_07489_));
 OR2_X1 _32956_ (.A1(_07065_),
    .A2(\icache.tag_tv_r [163]),
    .ZN(_07490_));
 NAND2_X1 _32957_ (.A1(_07111_),
    .A2(\icache.tag_tv_r [178]),
    .ZN(_07491_));
 NAND3_X1 _32958_ (.A1(_07489_),
    .A2(_07490_),
    .A3(_07491_),
    .ZN(_07492_));
 XNOR2_X1 _32959_ (.A(_07135_),
    .B(\icache.tag_tv_r [175]),
    .ZN(_07493_));
 NAND2_X1 _32960_ (.A1(_07065_),
    .A2(\icache.tag_tv_r [163]),
    .ZN(_07494_));
 OR2_X1 _32961_ (.A1(_07148_),
    .A2(\icache.tag_tv_r [166]),
    .ZN(_07495_));
 NAND3_X1 _32962_ (.A1(_07493_),
    .A2(_07494_),
    .A3(_07495_),
    .ZN(_07496_));
 NOR4_X1 _32963_ (.A1(_07484_),
    .A2(_07488_),
    .A3(_07492_),
    .A4(_07496_),
    .ZN(_07497_));
 OR2_X1 _32964_ (.A1(_07172_),
    .A2(\icache.tag_tv_r [168]),
    .ZN(_07498_));
 OR2_X1 _32965_ (.A1(_07486_),
    .A2(\icache.tag_tv_r [172]),
    .ZN(_07499_));
 NAND2_X1 _32966_ (.A1(_07081_),
    .A2(\icache.tag_tv_r [187]),
    .ZN(_07500_));
 NOR2_X4 _32967_ (.A1(\icache.state_tv_r [13]),
    .A2(\icache.state_tv_r [12]),
    .ZN(_07501_));
 INV_X4 _32968_ (.A(_07501_),
    .ZN(_07502_));
 NAND4_X1 _32969_ (.A1(_07498_),
    .A2(_07499_),
    .A3(_07500_),
    .A4(_07502_),
    .ZN(_07503_));
 XNOR2_X2 _32970_ (.A(_07130_),
    .B(\icache.tag_tv_r [180]),
    .ZN(_07504_));
 NAND2_X1 _32971_ (.A1(_07149_),
    .A2(\icache.tag_tv_r [166]),
    .ZN(_07505_));
 OAI211_X1 _32972_ (.A(_07504_),
    .B(_07505_),
    .C1(_07111_),
    .C2(\icache.tag_tv_r [178]),
    .ZN(_07506_));
 OR2_X1 _32973_ (.A1(_07253_),
    .A2(\icache.tag_tv_r [170]),
    .ZN(_07507_));
 NAND2_X1 _32974_ (.A1(_07253_),
    .A2(\icache.tag_tv_r [170]),
    .ZN(_07508_));
 OAI211_X1 _32975_ (.A(_07507_),
    .B(_07508_),
    .C1(_07083_),
    .C2(\icache.tag_tv_r [183]),
    .ZN(_07509_));
 AOI22_X1 _32976_ (.A1(_07248_),
    .A2(_07483_),
    .B1(_07086_),
    .B2(\icache.tag_tv_r [185]),
    .ZN(_07510_));
 NAND2_X1 _32977_ (.A1(_07108_),
    .A2(\icache.tag_tv_r [176]),
    .ZN(_07511_));
 NAND2_X1 _32978_ (.A1(_07083_),
    .A2(\icache.tag_tv_r [183]),
    .ZN(_07512_));
 NAND3_X1 _32979_ (.A1(_07510_),
    .A2(_07511_),
    .A3(_07512_),
    .ZN(_07513_));
 NOR4_X1 _32980_ (.A1(_07503_),
    .A2(_07506_),
    .A3(_07509_),
    .A4(_07513_),
    .ZN(_07514_));
 NAND2_X2 _32981_ (.A1(_07497_),
    .A2(_07514_),
    .ZN(_07515_));
 NOR2_X4 _32982_ (.A1(_07481_),
    .A2(_07515_),
    .ZN(_07516_));
 INV_X1 _32983_ (.A(\icache.tag_tv_r [190]),
    .ZN(_07517_));
 AOI22_X1 _32984_ (.A1(_07517_),
    .A2(net1384),
    .B1(_07253_),
    .B2(\icache.tag_tv_r [197]),
    .ZN(_07518_));
 INV_X1 _32985_ (.A(\icache.tag_tv_r [213]),
    .ZN(_07519_));
 OAI221_X1 _32986_ (.A(_07518_),
    .B1(\icache.tag_tv_r [196]),
    .B2(_07069_),
    .C1(_07519_),
    .C2(_07092_),
    .ZN(_07520_));
 AOI22_X1 _32987_ (.A1(_07519_),
    .A2(_07092_),
    .B1(_07120_),
    .B2(\icache.tag_tv_r [215]),
    .ZN(_07521_));
 NAND2_X1 _32988_ (.A1(_07116_),
    .A2(\icache.tag_tv_r [211]),
    .ZN(_07522_));
 OAI211_X1 _32989_ (.A(_07521_),
    .B(_07522_),
    .C1(\icache.tag_tv_r [215]),
    .C2(_07120_),
    .ZN(_07523_));
 NOR2_X1 _32990_ (.A1(_07520_),
    .A2(_07523_),
    .ZN(_07524_));
 OAI22_X1 _32991_ (.A1(\icache.tag_tv_r [194]),
    .A2(_07052_),
    .B1(_07116_),
    .B2(\icache.tag_tv_r [211]),
    .ZN(_07525_));
 INV_X1 _32992_ (.A(\icache.tag_tv_r [192]),
    .ZN(_07526_));
 AOI221_X4 _32993_ (.A(_07525_),
    .B1(_07526_),
    .B2(_07186_),
    .C1(\icache.tag_tv_r [204]),
    .C2(_07099_),
    .ZN(_07527_));
 XNOR2_X2 _32994_ (.A(\icache.tag_tv_r [207]),
    .B(_07130_),
    .ZN(_07528_));
 AOI22_X1 _32995_ (.A1(\icache.tag_tv_r [192]),
    .A2(_07067_),
    .B1(_07052_),
    .B2(\icache.tag_tv_r [194]),
    .ZN(_07529_));
 AND4_X1 _32996_ (.A1(_07524_),
    .A2(_07527_),
    .A3(_07528_),
    .A4(_07529_),
    .ZN(_07530_));
 NOR2_X1 _32997_ (.A1(_07083_),
    .A2(\icache.tag_tv_r [210]),
    .ZN(_07531_));
 AOI21_X1 _32998_ (.A(_07531_),
    .B1(\icache.tag_tv_r [212]),
    .B2(_07086_),
    .ZN(_07532_));
 NAND2_X1 _32999_ (.A1(_07069_),
    .A2(\icache.tag_tv_r [196]),
    .ZN(_07533_));
 XNOR2_X2 _33000_ (.A(\icache.tag_tv_r [202]),
    .B(_07135_),
    .ZN(_07534_));
 XNOR2_X2 _33001_ (.A(_07193_),
    .B(\icache.tag_tv_r [189]),
    .ZN(_07535_));
 NAND4_X1 _33002_ (.A1(_07532_),
    .A2(_07533_),
    .A3(_07534_),
    .A4(_07535_),
    .ZN(_07536_));
 XNOR2_X2 _33003_ (.A(\icache.tag_tv_r [209]),
    .B(_07133_),
    .ZN(_07537_));
 INV_X1 _33004_ (.A(\icache.tag_tv_r [200]),
    .ZN(_07538_));
 OAI221_X1 _33005_ (.A(_07537_),
    .B1(_07538_),
    .B2(net1354),
    .C1(\icache.tag_tv_r [204]),
    .C2(_07099_),
    .ZN(_07539_));
 AOI22_X1 _33006_ (.A1(\icache.tag_tv_r [198]),
    .A2(_07168_),
    .B1(_07538_),
    .B2(net1354),
    .ZN(_07540_));
 NAND2_X1 _33007_ (.A1(_07083_),
    .A2(\icache.tag_tv_r [210]),
    .ZN(_07541_));
 OAI211_X1 _33008_ (.A(_07540_),
    .B(_07541_),
    .C1(\icache.tag_tv_r [198]),
    .C2(_07168_),
    .ZN(_07542_));
 NOR3_X1 _33009_ (.A1(_07536_),
    .A2(_07539_),
    .A3(_07542_),
    .ZN(_07543_));
 AND2_X1 _33010_ (.A1(_07530_),
    .A2(_07543_),
    .ZN(_07544_));
 NOR2_X1 _33011_ (.A1(_07108_),
    .A2(\icache.tag_tv_r [203]),
    .ZN(_07545_));
 NOR2_X1 _33012_ (.A1(_07253_),
    .A2(\icache.tag_tv_r [197]),
    .ZN(_07546_));
 NOR2_X1 _33013_ (.A1(_07545_),
    .A2(_07546_),
    .ZN(_07547_));
 INV_X1 _33014_ (.A(_07105_),
    .ZN(_07548_));
 NAND2_X1 _33015_ (.A1(_07548_),
    .A2(\icache.tag_tv_r [201]),
    .ZN(_07549_));
 OAI211_X1 _33016_ (.A(_07547_),
    .B(_07549_),
    .C1(\icache.tag_tv_r [199]),
    .C2(_07486_),
    .ZN(_07550_));
 AND2_X1 _33017_ (.A1(_07149_),
    .A2(\icache.tag_tv_r [193]),
    .ZN(_07551_));
 AND2_X1 _33018_ (.A1(_07108_),
    .A2(\icache.tag_tv_r [203]),
    .ZN(_07552_));
 NAND2_X1 _33019_ (.A1(_07486_),
    .A2(\icache.tag_tv_r [199]),
    .ZN(_07553_));
 OAI21_X1 _33020_ (.A(_07553_),
    .B1(\icache.tag_tv_r [201]),
    .B2(_07548_),
    .ZN(_07554_));
 OR4_X1 _33021_ (.A1(_07550_),
    .A2(_07551_),
    .A3(_07552_),
    .A4(_07554_),
    .ZN(_07555_));
 INV_X1 _33022_ (.A(\icache.tag_tv_r [191]),
    .ZN(_07556_));
 AOI22_X1 _33023_ (.A1(_07556_),
    .A2(_07370_),
    .B1(_07172_),
    .B2(\icache.tag_tv_r [195]),
    .ZN(_07557_));
 OR2_X1 _33024_ (.A1(_07081_),
    .A2(\icache.tag_tv_r [214]),
    .ZN(_07558_));
 OAI211_X1 _33025_ (.A(_07557_),
    .B(_07558_),
    .C1(\icache.tag_tv_r [208]),
    .C2(_07101_),
    .ZN(_07559_));
 OR2_X1 _33026_ (.A1(_07172_),
    .A2(\icache.tag_tv_r [195]),
    .ZN(_07560_));
 OAI21_X1 _33027_ (.A(_07560_),
    .B1(_07556_),
    .B2(_07370_),
    .ZN(_07561_));
 NOR2_X4 _33028_ (.A1(\icache.state_tv_r [15]),
    .A2(\icache.state_tv_r [14]),
    .ZN(_07562_));
 NOR2_X1 _33029_ (.A1(_07149_),
    .A2(\icache.tag_tv_r [193]),
    .ZN(_07563_));
 OR4_X1 _33030_ (.A1(_07559_),
    .A2(_07561_),
    .A3(_07562_),
    .A4(_07563_),
    .ZN(_07564_));
 AOI22_X2 _33031_ (.A1(\icache.tag_tv_r [205]),
    .A2(_07111_),
    .B1(_07050_),
    .B2(\icache.tag_tv_r [206]),
    .ZN(_07565_));
 OAI221_X2 _33032_ (.A(_07565_),
    .B1(_07517_),
    .B2(net1384),
    .C1(\icache.tag_tv_r [206]),
    .C2(_07050_),
    .ZN(_07566_));
 NOR2_X1 _33033_ (.A1(_07086_),
    .A2(\icache.tag_tv_r [212]),
    .ZN(_07567_));
 AOI21_X1 _33034_ (.A(_07567_),
    .B1(\icache.tag_tv_r [208]),
    .B2(_07101_),
    .ZN(_07568_));
 NAND2_X1 _33035_ (.A1(_07081_),
    .A2(\icache.tag_tv_r [214]),
    .ZN(_07569_));
 OAI211_X2 _33036_ (.A(_07568_),
    .B(_07569_),
    .C1(\icache.tag_tv_r [205]),
    .C2(_07111_),
    .ZN(_07570_));
 NOR4_X2 _33037_ (.A1(_07555_),
    .A2(_07564_),
    .A3(_07566_),
    .A4(_07570_),
    .ZN(_07571_));
 AND2_X4 _33038_ (.A1(_07544_),
    .A2(_07571_),
    .ZN(_07572_));
 OAI21_X4 _33039_ (.A(_07462_),
    .B1(net1213),
    .B2(_07572_),
    .ZN(_07573_));
 INV_X1 _33040_ (.A(_07573_),
    .ZN(_07574_));
 NAND3_X2 _33041_ (.A1(_07147_),
    .A2(_07461_),
    .A3(_07214_),
    .ZN(_07575_));
 NOR3_X2 _33042_ (.A1(_07283_),
    .A2(_07459_),
    .A3(_07342_),
    .ZN(_07576_));
 NAND3_X4 _33043_ (.A1(_07146_),
    .A2(_07403_),
    .A3(_07576_),
    .ZN(_07577_));
 AND2_X4 _33044_ (.A1(_07575_),
    .A2(_07577_),
    .ZN(_07578_));
 INV_X1 _33045_ (.A(_07578_),
    .ZN(_07579_));
 OAI21_X4 _33046_ (.A(_07048_),
    .B1(_07574_),
    .B2(_07579_),
    .ZN(\icache.stat_mem.w_mask_i [1]));
 INV_X16 _33047_ (.A(_00000_),
    .ZN(_07580_));
 NAND3_X4 _33048_ (.A1(_07573_),
    .A2(_07580_),
    .A3(_07578_),
    .ZN(\icache.stat_mem.w_mask_i [2]));
 OAI211_X4 _33049_ (.A(_07461_),
    .B(_07048_),
    .C1(_07214_),
    .C2(_07146_),
    .ZN(_07581_));
 INV_X32 _33050_ (.A(_07581_),
    .ZN(\icache.stat_mem.data_i [2]));
 OAI21_X4 _33051_ (.A(_07343_),
    .B1(_07402_),
    .B2(_07459_),
    .ZN(_07582_));
 NAND2_X4 _33052_ (.A1(_07573_),
    .A2(_07582_),
    .ZN(_07583_));
 AOI21_X4 _33053_ (.A(\icache.stat_mem.data_i [2]),
    .B1(_07583_),
    .B2(_07048_),
    .ZN(\icache.stat_mem.w_mask_i [3]));
 NAND2_X4 _33054_ (.A1(_07582_),
    .A2(_07048_),
    .ZN(\icache.stat_mem.w_mask_i [4]));
 NAND3_X4 _33055_ (.A1(_07575_),
    .A2(_07577_),
    .A3(_07048_),
    .ZN(\icache.stat_mem.w_mask_i [5]));
 INV_X1 _33056_ (.A(_07283_),
    .ZN(_07584_));
 INV_X1 _33057_ (.A(_07342_),
    .ZN(_07585_));
 NAND3_X1 _33058_ (.A1(_07584_),
    .A2(_07585_),
    .A3(_07460_),
    .ZN(_07586_));
 NOR3_X2 _33059_ (.A1(_07146_),
    .A2(_07586_),
    .A3(_07402_),
    .ZN(_07587_));
 NAND3_X2 _33060_ (.A1(_07587_),
    .A2(_07215_),
    .A3(net1215),
    .ZN(_07588_));
 INV_X1 _33061_ (.A(net1214),
    .ZN(_07589_));
 NAND3_X2 _33062_ (.A1(_07587_),
    .A2(_07215_),
    .A3(_07589_),
    .ZN(_07590_));
 INV_X1 _33063_ (.A(_07572_),
    .ZN(_07591_));
 OAI211_X4 _33064_ (.A(_07048_),
    .B(_07588_),
    .C1(_07590_),
    .C2(_07591_),
    .ZN(\icache.stat_mem.w_mask_i [6]));
 AND3_X4 _33065_ (.A1(_07573_),
    .A2(_07048_),
    .A3(_07578_),
    .ZN(\icache.stat_mem.data_i [0]));
 NOR2_X4 _33066_ (.A1(_07583_),
    .A2(net1001),
    .ZN(\icache.stat_mem.data_i [1]));
 NOR2_X2 _33067_ (.A1(_07590_),
    .A2(_07591_),
    .ZN(_07592_));
 NAND3_X1 _33068_ (.A1(_07343_),
    .A2(_07402_),
    .A3(_07460_),
    .ZN(_07593_));
 INV_X1 _33069_ (.A(_07245_),
    .ZN(_07594_));
 AND2_X1 _33070_ (.A1(_07265_),
    .A2(_07282_),
    .ZN(_07595_));
 INV_X1 _33071_ (.A(_07595_),
    .ZN(_07596_));
 OAI21_X4 _33072_ (.A(_07342_),
    .B1(_07594_),
    .B2(_07596_),
    .ZN(_07597_));
 NAND2_X1 _33073_ (.A1(_07593_),
    .A2(_07597_),
    .ZN(_07598_));
 AOI21_X1 _33074_ (.A(_07598_),
    .B1(_07587_),
    .B2(_07214_),
    .ZN(_07599_));
 INV_X2 _33075_ (.A(_07599_),
    .ZN(_07600_));
 NOR4_X4 _33076_ (.A1(_07583_),
    .A2(_07592_),
    .A3(\icache.stat_mem.w_mask_i [5]),
    .A4(_07600_),
    .ZN(\icache.stat_mem.data_i [3]));
 INV_X4 _33077_ (.A(_07048_),
    .ZN(_07601_));
 BUF_X16 _33078_ (.A(_07601_),
    .Z(_07602_));
 NOR4_X4 _33079_ (.A1(_07460_),
    .A2(_07283_),
    .A3(_07602_),
    .A4(_07342_),
    .ZN(\icache.stat_mem.data_i [4]));
 AND3_X4 _33080_ (.A1(_07461_),
    .A2(_07048_),
    .A3(_07146_),
    .ZN(\icache.stat_mem.data_i [5]));
 NAND2_X1 _33081_ (.A1(_07461_),
    .A2(_07147_),
    .ZN(_07603_));
 NOR4_X4 _33082_ (.A1(_07603_),
    .A2(_07602_),
    .A3(_07214_),
    .A4(_07589_),
    .ZN(\icache.stat_mem.data_i [6]));
 INV_X2 _33083_ (.A(\icache.lce.lce_cmd_inst.state_r [1]),
    .ZN(_07604_));
 BUF_X4 _33084_ (.A(\icache.lce.lce_cmd_inst.state_r [0]),
    .Z(_07605_));
 NOR2_X4 _33085_ (.A1(_07604_),
    .A2(_07605_),
    .ZN(_07606_));
 BUF_X32 _33086_ (.A(_07606_),
    .Z(_07607_));
 BUF_X32 _33087_ (.A(_07607_),
    .Z(_07608_));
 BUF_X32 _33088_ (.A(_07608_),
    .Z(lce_data_cmd_v_o));
 INV_X1 _33089_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.head_r ),
    .ZN(_07609_));
 NAND2_X1 _33090_ (.A1(_07609_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [50]),
    .ZN(_07610_));
 NAND2_X1 _33091_ (.A1(\icache.lce.lce_cmd_inst.rv_adapter.head_r ),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [103]),
    .ZN(_07611_));
 NAND2_X4 _33092_ (.A1(_07610_),
    .A2(_07611_),
    .ZN(_07612_));
 BUF_X8 _33093_ (.A(_07609_),
    .Z(_07613_));
 NAND2_X2 _33094_ (.A1(_07613_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [49]),
    .ZN(_07614_));
 NAND2_X2 _33095_ (.A1(\icache.lce.lce_cmd_inst.rv_adapter.head_r ),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [102]),
    .ZN(_07615_));
 NAND2_X2 _33096_ (.A1(_07614_),
    .A2(_07615_),
    .ZN(_07616_));
 NOR2_X2 _33097_ (.A1(_07612_),
    .A2(_07616_),
    .ZN(_07617_));
 BUF_X8 _33098_ (.A(_07617_),
    .Z(_07618_));
 NAND2_X2 _33099_ (.A1(_07613_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [48]),
    .ZN(_07619_));
 NAND2_X2 _33100_ (.A1(\icache.lce.lce_cmd_inst.rv_adapter.head_r ),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [101]),
    .ZN(_07620_));
 AOI211_X2 _33101_ (.A(\icache.lce.lce_cmd_inst.state_r [1]),
    .B(\icache.lce.lce_cmd_inst.state_r [0]),
    .C1(_07619_),
    .C2(_07620_),
    .ZN(_07621_));
 BUF_X8 _33102_ (.A(_07613_),
    .Z(_07622_));
 NAND2_X1 _33103_ (.A1(_07622_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [15]),
    .ZN(_07623_));
 BUF_X8 _33104_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.head_r ),
    .Z(_07624_));
 NAND2_X1 _33105_ (.A1(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [68]),
    .A2(_07624_),
    .ZN(_07625_));
 NAND2_X4 _33106_ (.A1(_07623_),
    .A2(_07625_),
    .ZN(_07626_));
 NAND4_X2 _33107_ (.A1(_07618_),
    .A2(net1262),
    .A3(_07602_),
    .A4(_07626_),
    .ZN(_07627_));
 INV_X2 _33108_ (.A(\icache.addr_tv_r [6]),
    .ZN(_07628_));
 OAI21_X4 _33109_ (.A(_07627_),
    .B1(_07602_),
    .B2(_07628_),
    .ZN(\icache.stat_mem.addr_i [0]));
 BUF_X8 _33110_ (.A(_07613_),
    .Z(_07629_));
 NAND2_X1 _33111_ (.A1(_07629_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [16]),
    .ZN(_07630_));
 NAND2_X1 _33112_ (.A1(_07624_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [69]),
    .ZN(_07631_));
 NAND2_X4 _33113_ (.A1(_07630_),
    .A2(_07631_),
    .ZN(_07632_));
 NAND4_X2 _33114_ (.A1(_07618_),
    .A2(net1262),
    .A3(_07602_),
    .A4(_07632_),
    .ZN(_07633_));
 INV_X2 _33115_ (.A(\icache.addr_tv_r [7]),
    .ZN(_07634_));
 OAI21_X4 _33116_ (.A(_07633_),
    .B1(_07602_),
    .B2(_07634_),
    .ZN(\icache.stat_mem.addr_i [1]));
 NOR2_X1 _33117_ (.A1(_07629_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [70]),
    .ZN(_07635_));
 NOR2_X1 _33118_ (.A1(_07624_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [17]),
    .ZN(_07636_));
 NOR2_X4 _33119_ (.A1(_07635_),
    .A2(_07636_),
    .ZN(_07637_));
 NAND4_X2 _33120_ (.A1(_07618_),
    .A2(net1262),
    .A3(_07601_),
    .A4(_07637_),
    .ZN(_07638_));
 INV_X2 _33121_ (.A(\icache.addr_tv_r [8]),
    .ZN(_07639_));
 OAI21_X4 _33122_ (.A(_07638_),
    .B1(_07602_),
    .B2(_07639_),
    .ZN(\icache.stat_mem.addr_i [2]));
 NAND2_X1 _33123_ (.A1(_07629_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [18]),
    .ZN(_07640_));
 NAND2_X1 _33124_ (.A1(_07624_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [71]),
    .ZN(_07641_));
 NAND2_X4 _33125_ (.A1(_07640_),
    .A2(_07641_),
    .ZN(_07642_));
 NAND4_X4 _33126_ (.A1(_07618_),
    .A2(net1262),
    .A3(_07601_),
    .A4(_07642_),
    .ZN(_07643_));
 INV_X2 _33127_ (.A(\icache.addr_tv_r [9]),
    .ZN(_07644_));
 OAI21_X4 _33128_ (.A(_07643_),
    .B1(_07602_),
    .B2(_07644_),
    .ZN(\icache.stat_mem.addr_i [3]));
 NAND2_X1 _33129_ (.A1(_07629_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [19]),
    .ZN(_07645_));
 NAND2_X1 _33130_ (.A1(_07624_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [72]),
    .ZN(_07646_));
 NAND2_X4 _33131_ (.A1(_07645_),
    .A2(_07646_),
    .ZN(_07647_));
 NAND4_X2 _33132_ (.A1(_07618_),
    .A2(net1262),
    .A3(_07601_),
    .A4(_07647_),
    .ZN(_07648_));
 INV_X2 _33133_ (.A(\icache.addr_tv_r [10]),
    .ZN(_07649_));
 OAI21_X4 _33134_ (.A(_07648_),
    .B1(_07602_),
    .B2(_07649_),
    .ZN(\icache.stat_mem.addr_i [4]));
 NOR2_X1 _33135_ (.A1(_07613_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [73]),
    .ZN(_07650_));
 NOR2_X1 _33136_ (.A1(_07624_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [20]),
    .ZN(_07651_));
 NOR2_X4 _33137_ (.A1(_07650_),
    .A2(_07651_),
    .ZN(_07652_));
 NAND4_X4 _33138_ (.A1(_07618_),
    .A2(net1262),
    .A3(_07601_),
    .A4(_07652_),
    .ZN(_07653_));
 INV_X2 _33139_ (.A(\icache.addr_tv_r [11]),
    .ZN(_07654_));
 OAI21_X4 _33140_ (.A(_07653_),
    .B1(_07602_),
    .B2(_07654_),
    .ZN(\icache.stat_mem.addr_i [5]));
 AND2_X2 _33141_ (.A1(_07617_),
    .A2(net1261),
    .ZN(_07655_));
 AND2_X1 _33142_ (.A1(_07655_),
    .A2(_00001_),
    .ZN(_07656_));
 AND3_X1 _33143_ (.A1(_07473_),
    .A2(_07499_),
    .A3(_07487_),
    .ZN(_07657_));
 AND3_X1 _33144_ (.A1(_07469_),
    .A2(_07471_),
    .A3(_07498_),
    .ZN(_07658_));
 AND4_X1 _33145_ (.A1(_07467_),
    .A2(_07658_),
    .A3(_07505_),
    .A4(_07495_),
    .ZN(_07659_));
 AND3_X1 _33146_ (.A1(_07476_),
    .A2(_07490_),
    .A3(_07494_),
    .ZN(_07660_));
 AND3_X1 _33147_ (.A1(_07659_),
    .A2(_07480_),
    .A3(_07660_),
    .ZN(_07661_));
 AND3_X1 _33148_ (.A1(_07485_),
    .A2(_07507_),
    .A3(_07508_),
    .ZN(_07662_));
 AND2_X1 _33149_ (.A1(_07465_),
    .A2(_07493_),
    .ZN(_07663_));
 AND4_X1 _33150_ (.A1(_07470_),
    .A2(_07663_),
    .A3(_07511_),
    .A4(_07482_),
    .ZN(_07664_));
 AND4_X1 _33151_ (.A1(_07657_),
    .A2(_07661_),
    .A3(_07662_),
    .A4(_07664_),
    .ZN(_07665_));
 XNOR2_X1 _33152_ (.A(_07248_),
    .B(\icache.tag_tv_r [179]),
    .ZN(_07666_));
 XNOR2_X1 _33153_ (.A(net1348),
    .B(\icache.tag_tv_r [178]),
    .ZN(_07667_));
 NAND4_X1 _33154_ (.A1(_07474_),
    .A2(_07504_),
    .A3(_07666_),
    .A4(_07667_),
    .ZN(_07668_));
 XNOR2_X1 _33155_ (.A(net1334),
    .B(\icache.tag_tv_r [183]),
    .ZN(_07669_));
 XNOR2_X1 _33156_ (.A(net1329),
    .B(\icache.tag_tv_r [185]),
    .ZN(_07670_));
 NAND4_X1 _33157_ (.A1(_07466_),
    .A2(_07489_),
    .A3(_07669_),
    .A4(_07670_),
    .ZN(_07671_));
 NOR2_X1 _33158_ (.A1(_07668_),
    .A2(_07671_),
    .ZN(_07672_));
 XNOR2_X1 _33159_ (.A(net1323),
    .B(\icache.tag_tv_r [187]),
    .ZN(_07673_));
 AND4_X1 _33160_ (.A1(_07477_),
    .A2(_07672_),
    .A3(_07463_),
    .A4(_07673_),
    .ZN(_07674_));
 NAND3_X2 _33161_ (.A1(_07665_),
    .A2(_07502_),
    .A3(_07674_),
    .ZN(_07675_));
 XNOR2_X1 _33162_ (.A(_07133_),
    .B(\icache.tag_tv_r [155]),
    .ZN(_07676_));
 XNOR2_X1 _33163_ (.A(net1342),
    .B(\icache.tag_tv_r [153]),
    .ZN(_07677_));
 XNOR2_X1 _33164_ (.A(net1345),
    .B(\icache.tag_tv_r [151]),
    .ZN(_07678_));
 XNOR2_X1 _33165_ (.A(net1337),
    .B(\icache.tag_tv_r [154]),
    .ZN(_07679_));
 XNOR2_X1 _33166_ (.A(_07248_),
    .B(\icache.tag_tv_r [152]),
    .ZN(_07680_));
 AND4_X1 _33167_ (.A1(_07677_),
    .A2(_07678_),
    .A3(_07679_),
    .A4(_07680_),
    .ZN(_07681_));
 XNOR2_X1 _33168_ (.A(_07156_),
    .B(\icache.tag_tv_r [157]),
    .ZN(_07682_));
 AND3_X1 _33169_ (.A1(_07682_),
    .A2(_07206_),
    .A3(_07175_),
    .ZN(_07683_));
 XNOR2_X1 _33170_ (.A(net1334),
    .B(\icache.tag_tv_r [156]),
    .ZN(_07684_));
 AND4_X1 _33171_ (.A1(_07676_),
    .A2(_07681_),
    .A3(_07683_),
    .A4(_07684_),
    .ZN(_07685_));
 XNOR2_X1 _33172_ (.A(_07160_),
    .B(\icache.tag_tv_r [161]),
    .ZN(_07686_));
 XNOR2_X1 _33173_ (.A(_07092_),
    .B(\icache.tag_tv_r [159]),
    .ZN(_07687_));
 XNOR2_X1 _33174_ (.A(net1324),
    .B(\icache.tag_tv_r [160]),
    .ZN(_07688_));
 NAND4_X1 _33175_ (.A1(_07685_),
    .A2(_07686_),
    .A3(_07687_),
    .A4(_07688_),
    .ZN(_07689_));
 INV_X1 _33176_ (.A(_07196_),
    .ZN(_07690_));
 XNOR2_X1 _33177_ (.A(_07190_),
    .B(\icache.tag_tv_r [150]),
    .ZN(_07691_));
 AND4_X1 _33178_ (.A1(_07690_),
    .A2(_07155_),
    .A3(_07177_),
    .A4(_07691_),
    .ZN(_07692_));
 XNOR2_X1 _33179_ (.A(_07118_),
    .B(\icache.tag_tv_r [145]),
    .ZN(_07693_));
 XNOR2_X1 _33180_ (.A(net1354),
    .B(\icache.tag_tv_r [146]),
    .ZN(_07694_));
 XNOR2_X1 _33181_ (.A(net1359),
    .B(\icache.tag_tv_r [144]),
    .ZN(_07695_));
 AND4_X1 _33182_ (.A1(_07179_),
    .A2(_07693_),
    .A3(_07694_),
    .A4(_07695_),
    .ZN(_07696_));
 XNOR2_X1 _33183_ (.A(_07113_),
    .B(\icache.tag_tv_r [141]),
    .ZN(_07697_));
 XNOR2_X1 _33184_ (.A(_07123_),
    .B(\icache.tag_tv_r [139]),
    .ZN(_07698_));
 XNOR2_X1 _33185_ (.A(net1365),
    .B(\icache.tag_tv_r [142]),
    .ZN(_07699_));
 AND4_X1 _33186_ (.A1(_07178_),
    .A2(_07697_),
    .A3(_07698_),
    .A4(_07699_),
    .ZN(_07700_));
 XNOR2_X1 _33187_ (.A(net1379),
    .B(net1268),
    .ZN(_07701_));
 XNOR2_X1 _33188_ (.A(_07186_),
    .B(net1267),
    .ZN(_07702_));
 XNOR2_X1 _33189_ (.A(_07193_),
    .B(net1270),
    .ZN(_07703_));
 AND4_X1 _33190_ (.A1(_07183_),
    .A2(_07701_),
    .A3(_07702_),
    .A4(_07703_),
    .ZN(_07704_));
 NAND4_X2 _33191_ (.A1(_07692_),
    .A2(_07696_),
    .A3(_07700_),
    .A4(_07704_),
    .ZN(_07705_));
 NOR3_X1 _33192_ (.A1(_07689_),
    .A2(_07198_),
    .A3(_07705_),
    .ZN(_07706_));
 XNOR2_X1 _33193_ (.A(_07107_),
    .B(net1284),
    .ZN(_07707_));
 NAND3_X1 _33194_ (.A1(_07707_),
    .A2(_07100_),
    .A3(_07143_),
    .ZN(_07708_));
 XOR2_X2 _33195_ (.A(_07105_),
    .B(net1288),
    .Z(_07709_));
 NOR2_X1 _33196_ (.A1(_07136_),
    .A2(_07135_),
    .ZN(_07710_));
 NOR4_X1 _33197_ (.A1(_07708_),
    .A2(_07709_),
    .A3(_07058_),
    .A4(_07710_),
    .ZN(_07711_));
 NAND3_X1 _33198_ (.A1(_07119_),
    .A2(_07056_),
    .A3(_07142_),
    .ZN(_07712_));
 INV_X1 _33199_ (.A(_07129_),
    .ZN(_07713_));
 NOR4_X1 _33200_ (.A1(_07712_),
    .A2(_07713_),
    .A3(_07060_),
    .A4(_07061_),
    .ZN(_07714_));
 XNOR2_X1 _33201_ (.A(net1368),
    .B(net1296),
    .ZN(_07715_));
 XNOR2_X1 _33202_ (.A(_07123_),
    .B(net1299),
    .ZN(_07716_));
 XNOR2_X1 _33203_ (.A(net1365),
    .B(net1293),
    .ZN(_07717_));
 XNOR2_X1 _33204_ (.A(net1373),
    .B(net1297),
    .ZN(_07718_));
 AND4_X1 _33205_ (.A1(_07715_),
    .A2(_07716_),
    .A3(_07717_),
    .A4(_07718_),
    .ZN(_07719_));
 XNOR2_X1 _33206_ (.A(net1377),
    .B(net1301),
    .ZN(_07720_));
 XNOR2_X1 _33207_ (.A(net1374),
    .B(net1300),
    .ZN(_07721_));
 XNOR2_X1 _33208_ (.A(net1380),
    .B(net1302),
    .ZN(_07722_));
 AND4_X1 _33209_ (.A1(_07141_),
    .A2(_07720_),
    .A3(_07721_),
    .A4(_07722_),
    .ZN(_07723_));
 AND4_X1 _33210_ (.A1(_07711_),
    .A2(_07714_),
    .A3(_07719_),
    .A4(_07723_),
    .ZN(_07724_));
 XNOR2_X1 _33211_ (.A(_07156_),
    .B(net1274),
    .ZN(_07725_));
 AND3_X1 _33212_ (.A1(_07725_),
    .A2(_07079_),
    .A3(_07087_),
    .ZN(_07726_));
 NAND4_X1 _33213_ (.A1(_07726_),
    .A2(_07076_),
    .A3(_07085_),
    .A4(_07134_),
    .ZN(_07727_));
 XNOR2_X1 _33214_ (.A(_07160_),
    .B(net1271),
    .ZN(_07728_));
 NAND4_X1 _33215_ (.A1(_07093_),
    .A2(_07728_),
    .A3(_07073_),
    .A4(_07082_),
    .ZN(_07729_));
 XNOR2_X1 _33216_ (.A(_07130_),
    .B(net1278),
    .ZN(_07730_));
 NAND3_X1 _33217_ (.A1(_07730_),
    .A2(_07102_),
    .A3(_07089_),
    .ZN(_07731_));
 XNOR2_X1 _33218_ (.A(net1345),
    .B(net1280),
    .ZN(_07732_));
 INV_X1 _33219_ (.A(_07051_),
    .ZN(_07733_));
 NAND3_X1 _33220_ (.A1(_07732_),
    .A2(_07733_),
    .A3(_07077_),
    .ZN(_07734_));
 NOR4_X1 _33221_ (.A1(_07727_),
    .A2(_07729_),
    .A3(_07731_),
    .A4(_07734_),
    .ZN(_07735_));
 AND3_X1 _33222_ (.A1(_07724_),
    .A2(_07095_),
    .A3(_07735_),
    .ZN(_07736_));
 NOR2_X2 _33223_ (.A1(_07706_),
    .A2(_07736_),
    .ZN(_07737_));
 NAND2_X1 _33224_ (.A1(_07172_),
    .A2(\icache.tag_tv_r [195]),
    .ZN(_07738_));
 OR2_X1 _33225_ (.A1(_07069_),
    .A2(\icache.tag_tv_r [196]),
    .ZN(_07739_));
 NAND4_X1 _33226_ (.A1(_07738_),
    .A2(_07560_),
    .A3(_07533_),
    .A4(_07739_),
    .ZN(_07740_));
 XOR2_X1 _33227_ (.A(\icache.tag_tv_r [194]),
    .B(net1372),
    .Z(_07741_));
 NOR4_X1 _33228_ (.A1(_07740_),
    .A2(_07741_),
    .A3(_07563_),
    .A4(_07551_),
    .ZN(_07742_));
 OR2_X1 _33229_ (.A1(_07548_),
    .A2(\icache.tag_tv_r [201]),
    .ZN(_07743_));
 NAND3_X1 _33230_ (.A1(_07534_),
    .A2(_07549_),
    .A3(_07743_),
    .ZN(_07744_));
 XOR2_X2 _33231_ (.A(\icache.tag_tv_r [204]),
    .B(net1350),
    .Z(_07745_));
 NOR4_X1 _33232_ (.A1(_07744_),
    .A2(_07745_),
    .A3(_07545_),
    .A4(_07552_),
    .ZN(_07746_));
 XNOR2_X1 _33233_ (.A(\icache.tag_tv_r [190]),
    .B(net1383),
    .ZN(_07747_));
 XNOR2_X1 _33234_ (.A(\icache.tag_tv_r [192]),
    .B(_07186_),
    .ZN(_07748_));
 XNOR2_X1 _33235_ (.A(\icache.tag_tv_r [191]),
    .B(_07370_),
    .ZN(_07749_));
 AND4_X1 _33236_ (.A1(_07535_),
    .A2(_07747_),
    .A3(_07748_),
    .A4(_07749_),
    .ZN(_07750_));
 XNOR2_X1 _33237_ (.A(\icache.tag_tv_r [200]),
    .B(net1354),
    .ZN(_07751_));
 XNOR2_X1 _33238_ (.A(\icache.tag_tv_r [197]),
    .B(_07128_),
    .ZN(_07752_));
 XNOR2_X1 _33239_ (.A(\icache.tag_tv_r [198]),
    .B(net1360),
    .ZN(_07753_));
 XNOR2_X1 _33240_ (.A(\icache.tag_tv_r [199]),
    .B(_07118_),
    .ZN(_07754_));
 AND4_X1 _33241_ (.A1(_07751_),
    .A2(_07752_),
    .A3(_07753_),
    .A4(_07754_),
    .ZN(_07755_));
 NAND4_X1 _33242_ (.A1(_07742_),
    .A2(_07746_),
    .A3(_07750_),
    .A4(_07755_),
    .ZN(_07756_));
 XNOR2_X1 _33243_ (.A(\icache.tag_tv_r [211]),
    .B(_07156_),
    .ZN(_07757_));
 XNOR2_X1 _33244_ (.A(\icache.tag_tv_r [212]),
    .B(net1328),
    .ZN(_07758_));
 XNOR2_X1 _33245_ (.A(\icache.tag_tv_r [210]),
    .B(net1334),
    .ZN(_07759_));
 AND4_X1 _33246_ (.A1(_07537_),
    .A2(_07757_),
    .A3(_07758_),
    .A4(_07759_),
    .ZN(_07760_));
 XNOR2_X1 _33247_ (.A(\icache.tag_tv_r [208]),
    .B(net1338),
    .ZN(_07761_));
 XNOR2_X1 _33248_ (.A(\icache.tag_tv_r [206]),
    .B(_07248_),
    .ZN(_07762_));
 XNOR2_X1 _33249_ (.A(\icache.tag_tv_r [205]),
    .B(net1348),
    .ZN(_07763_));
 AND4_X1 _33250_ (.A1(_07528_),
    .A2(_07761_),
    .A3(_07762_),
    .A4(_07763_),
    .ZN(_07764_));
 XNOR2_X1 _33251_ (.A(\icache.tag_tv_r [215]),
    .B(_07160_),
    .ZN(_07765_));
 XNOR2_X1 _33252_ (.A(\icache.tag_tv_r [213]),
    .B(_07092_),
    .ZN(_07766_));
 AND4_X1 _33253_ (.A1(_07558_),
    .A2(_07765_),
    .A3(_07766_),
    .A4(_07569_),
    .ZN(_07767_));
 NAND3_X1 _33254_ (.A1(_07760_),
    .A2(_07764_),
    .A3(_07767_),
    .ZN(_07768_));
 OR3_X2 _33255_ (.A1(_07756_),
    .A2(_07562_),
    .A3(_07768_),
    .ZN(_07769_));
 AND3_X4 _33256_ (.A1(_07675_),
    .A2(_07737_),
    .A3(_07769_),
    .ZN(_07770_));
 XNOR2_X1 _33257_ (.A(_07133_),
    .B(\icache.tag_tv_r [74]),
    .ZN(_07771_));
 AND2_X1 _33258_ (.A1(_07110_),
    .A2(\icache.tag_tv_r [70]),
    .ZN(_07772_));
 NOR4_X1 _33259_ (.A1(_07772_),
    .A2(_07420_),
    .A3(_07412_),
    .A4(_07426_),
    .ZN(_07773_));
 XNOR2_X1 _33260_ (.A(_07130_),
    .B(\icache.tag_tv_r [72]),
    .ZN(_07774_));
 AND4_X1 _33261_ (.A1(_07451_),
    .A2(_07773_),
    .A3(_07441_),
    .A4(_07774_),
    .ZN(_07775_));
 AND2_X1 _33262_ (.A1(_07116_),
    .A2(\icache.tag_tv_r [76]),
    .ZN(_07776_));
 AND2_X1 _33263_ (.A1(_07086_),
    .A2(\icache.tag_tv_r [77]),
    .ZN(_07777_));
 NOR4_X1 _33264_ (.A1(_07776_),
    .A2(_07777_),
    .A3(_07410_),
    .A4(_07422_),
    .ZN(_07778_));
 XNOR2_X1 _33265_ (.A(net1331),
    .B(\icache.tag_tv_r [75]),
    .ZN(_07779_));
 AND4_X1 _33266_ (.A1(_07771_),
    .A2(_07775_),
    .A3(_07778_),
    .A4(_07779_),
    .ZN(_07780_));
 XNOR2_X1 _33267_ (.A(_07092_),
    .B(\icache.tag_tv_r [78]),
    .ZN(_07781_));
 XNOR2_X1 _33268_ (.A(net1320),
    .B(\icache.tag_tv_r [79]),
    .ZN(_07782_));
 NAND4_X2 _33269_ (.A1(_07780_),
    .A2(_07404_),
    .A3(_07781_),
    .A4(_07782_),
    .ZN(_07783_));
 NAND3_X1 _33270_ (.A1(_07429_),
    .A2(_07444_),
    .A3(_07455_),
    .ZN(_07784_));
 XOR2_X1 _33271_ (.A(_07107_),
    .B(\icache.tag_tv_r [68]),
    .Z(_07785_));
 NOR2_X1 _33272_ (.A1(_07456_),
    .A2(_07190_),
    .ZN(_07786_));
 NOR4_X1 _33273_ (.A1(_07784_),
    .A2(_07785_),
    .A3(_07421_),
    .A4(_07786_),
    .ZN(_07787_));
 XNOR2_X1 _33274_ (.A(net1353),
    .B(\icache.tag_tv_r [65]),
    .ZN(_07788_));
 XNOR2_X1 _33275_ (.A(net1357),
    .B(\icache.tag_tv_r [63]),
    .ZN(_07789_));
 AND4_X1 _33276_ (.A1(_07406_),
    .A2(_07408_),
    .A3(_07788_),
    .A4(_07789_),
    .ZN(_07790_));
 XNOR2_X1 _33277_ (.A(_07113_),
    .B(\icache.tag_tv_r [60]),
    .ZN(_07791_));
 XNOR2_X1 _33278_ (.A(_07123_),
    .B(\icache.tag_tv_r [58]),
    .ZN(_07792_));
 XNOR2_X1 _33279_ (.A(net1362),
    .B(\icache.tag_tv_r [61]),
    .ZN(_07793_));
 AND4_X1 _33280_ (.A1(_07437_),
    .A2(_07791_),
    .A3(_07792_),
    .A4(_07793_),
    .ZN(_07794_));
 NAND2_X1 _33281_ (.A1(_07446_),
    .A2(_07193_),
    .ZN(_07795_));
 NAND4_X2 _33282_ (.A1(_07433_),
    .A2(_07450_),
    .A3(_07452_),
    .A4(_07795_),
    .ZN(_07796_));
 XOR2_X1 _33283_ (.A(_07370_),
    .B(\icache.tag_tv_r [56]),
    .Z(_07797_));
 XOR2_X2 _33284_ (.A(_07186_),
    .B(\icache.tag_tv_r [57]),
    .Z(_07798_));
 NOR3_X2 _33285_ (.A1(_07796_),
    .A2(_07797_),
    .A3(_07798_),
    .ZN(_07799_));
 NAND4_X2 _33286_ (.A1(_07787_),
    .A2(_07790_),
    .A3(_07794_),
    .A4(_07799_),
    .ZN(_07800_));
 NOR3_X2 _33287_ (.A1(_07783_),
    .A2(_07425_),
    .A3(_07800_),
    .ZN(_07801_));
 XNOR2_X1 _33288_ (.A(net1331),
    .B(\icache.tag_tv_r [102]),
    .ZN(_07802_));
 NAND4_X1 _33289_ (.A1(_07346_),
    .A2(_07356_),
    .A3(_07358_),
    .A4(_07802_),
    .ZN(_07803_));
 OR2_X1 _33290_ (.A1(_07111_),
    .A2(\icache.tag_tv_r [97]),
    .ZN(_07804_));
 NAND4_X1 _33291_ (.A1(_07804_),
    .A2(_07380_),
    .A3(_07360_),
    .A4(_07399_),
    .ZN(_07805_));
 XOR2_X1 _33292_ (.A(_07130_),
    .B(\icache.tag_tv_r [99]),
    .Z(_07806_));
 XOR2_X1 _33293_ (.A(net1335),
    .B(\icache.tag_tv_r [100]),
    .Z(_07807_));
 NOR4_X1 _33294_ (.A1(_07803_),
    .A2(_07805_),
    .A3(_07806_),
    .A4(_07807_),
    .ZN(_07808_));
 XNOR2_X1 _33295_ (.A(_07092_),
    .B(\icache.tag_tv_r [105]),
    .ZN(_07809_));
 XNOR2_X1 _33296_ (.A(net1320),
    .B(\icache.tag_tv_r [106]),
    .ZN(_07810_));
 AND4_X1 _33297_ (.A1(_07345_),
    .A2(_07808_),
    .A3(_07809_),
    .A4(_07810_),
    .ZN(_07811_));
 XNOR2_X1 _33298_ (.A(_07107_),
    .B(\icache.tag_tv_r [95]),
    .ZN(_07812_));
 XNOR2_X1 _33299_ (.A(_07190_),
    .B(\icache.tag_tv_r [96]),
    .ZN(_07813_));
 XNOR2_X1 _33300_ (.A(_07135_),
    .B(\icache.tag_tv_r [94]),
    .ZN(_07814_));
 AND4_X1 _33301_ (.A1(_07344_),
    .A2(_07812_),
    .A3(_07813_),
    .A4(_07814_),
    .ZN(_07815_));
 XNOR2_X1 _33302_ (.A(net1358),
    .B(\icache.tag_tv_r [90]),
    .ZN(_07816_));
 AND2_X1 _33303_ (.A1(_07347_),
    .A2(_07816_),
    .ZN(_07817_));
 AND4_X1 _33304_ (.A1(_07357_),
    .A2(_07817_),
    .A3(_07394_),
    .A4(_07379_),
    .ZN(_07818_));
 XNOR2_X1 _33305_ (.A(_07113_),
    .B(\icache.tag_tv_r [87]),
    .ZN(_07819_));
 NAND3_X1 _33306_ (.A1(_07819_),
    .A2(_07386_),
    .A3(_07392_),
    .ZN(_07820_));
 XOR2_X1 _33307_ (.A(_07123_),
    .B(\icache.tag_tv_r [85]),
    .Z(_07821_));
 NOR4_X1 _33308_ (.A1(_07820_),
    .A2(_07821_),
    .A3(_07366_),
    .A4(_07368_),
    .ZN(_07822_));
 XNOR2_X1 _33309_ (.A(net1381),
    .B(\icache.tag_tv_r [82]),
    .ZN(_07823_));
 NAND3_X1 _33310_ (.A1(_07823_),
    .A2(_07375_),
    .A3(_07381_),
    .ZN(_07824_));
 XOR2_X1 _33311_ (.A(_07370_),
    .B(\icache.tag_tv_r [83]),
    .Z(_07825_));
 NOR4_X1 _33312_ (.A1(_07824_),
    .A2(_07825_),
    .A3(_07390_),
    .A4(_07367_),
    .ZN(_07826_));
 AND4_X1 _33313_ (.A1(_07815_),
    .A2(_07818_),
    .A3(_07822_),
    .A4(_07826_),
    .ZN(_07827_));
 AND3_X1 _33314_ (.A1(_07811_),
    .A2(_07351_),
    .A3(_07827_),
    .ZN(_07828_));
 NOR2_X4 _33315_ (.A1(_07801_),
    .A2(_07828_),
    .ZN(_07829_));
 XNOR2_X1 _33316_ (.A(_07156_),
    .B(\icache.tag_tv_r [22]),
    .ZN(_07830_));
 AND3_X1 _33317_ (.A1(_07830_),
    .A2(_07262_),
    .A3(_07263_),
    .ZN(_07831_));
 XNOR2_X1 _33318_ (.A(_07133_),
    .B(\icache.tag_tv_r [20]),
    .ZN(_07832_));
 AND4_X1 _33319_ (.A1(_07226_),
    .A2(_07831_),
    .A3(_07230_),
    .A4(_07832_),
    .ZN(_07833_));
 XNOR2_X1 _33320_ (.A(net1335),
    .B(\icache.tag_tv_r [19]),
    .ZN(_07834_));
 NAND2_X1 _33321_ (.A1(_07249_),
    .A2(_07248_),
    .ZN(_07835_));
 AND3_X1 _33322_ (.A1(_07225_),
    .A2(_07835_),
    .A3(_07275_),
    .ZN(_07836_));
 AND4_X1 _33323_ (.A1(_07267_),
    .A2(_07833_),
    .A3(_07834_),
    .A4(_07836_),
    .ZN(_07837_));
 AND3_X1 _33324_ (.A1(_07239_),
    .A2(_07223_),
    .A3(_07280_),
    .ZN(_07838_));
 XNOR2_X1 _33325_ (.A(_07123_),
    .B(\icache.tag_tv_r [4]),
    .ZN(_07839_));
 AND4_X1 _33326_ (.A1(_07233_),
    .A2(_07838_),
    .A3(_07236_),
    .A4(_07839_),
    .ZN(_07840_));
 NAND2_X1 _33327_ (.A1(_07216_),
    .A2(_07193_),
    .ZN(_07841_));
 AND4_X1 _33328_ (.A1(_07234_),
    .A2(_07218_),
    .A3(_07841_),
    .A4(_07279_),
    .ZN(_07842_));
 AND4_X1 _33329_ (.A1(_07242_),
    .A2(_07840_),
    .A3(_07243_),
    .A4(_07842_),
    .ZN(_07843_));
 OR2_X1 _33330_ (.A1(_07162_),
    .A2(\icache.tag_tv_r [24]),
    .ZN(_07844_));
 XNOR2_X1 _33331_ (.A(net1317),
    .B(\icache.tag_tv_r [25]),
    .ZN(_07845_));
 AND4_X1 _33332_ (.A1(_07241_),
    .A2(_07260_),
    .A3(_07844_),
    .A4(_07845_),
    .ZN(_07846_));
 AND3_X1 _33333_ (.A1(_07270_),
    .A2(_07235_),
    .A3(_07229_),
    .ZN(_07847_));
 AND4_X1 _33334_ (.A1(_07222_),
    .A2(_07252_),
    .A3(_07268_),
    .A4(_07254_),
    .ZN(_07848_));
 AND3_X1 _33335_ (.A1(_07271_),
    .A2(_07221_),
    .A3(_07231_),
    .ZN(_07849_));
 AND3_X1 _33336_ (.A1(_07274_),
    .A2(_07228_),
    .A3(_07257_),
    .ZN(_07850_));
 AND4_X1 _33337_ (.A1(_07847_),
    .A2(_07848_),
    .A3(_07849_),
    .A4(_07850_),
    .ZN(_07851_));
 NAND4_X4 _33338_ (.A1(_07837_),
    .A2(_07843_),
    .A3(_07846_),
    .A4(_07851_),
    .ZN(_07852_));
 NOR2_X2 _33339_ (.A1(_07852_),
    .A2(_07255_),
    .ZN(_07853_));
 NAND2_X1 _33340_ (.A1(_07099_),
    .A2(\icache.tag_tv_r [42]),
    .ZN(_07854_));
 AND3_X1 _33341_ (.A1(_07303_),
    .A2(_07322_),
    .A3(_07854_),
    .ZN(_07855_));
 AND4_X1 _33342_ (.A1(_07297_),
    .A2(_07855_),
    .A3(_07298_),
    .A4(_07332_),
    .ZN(_07856_));
 XNOR2_X1 _33343_ (.A(_07128_),
    .B(\icache.tag_tv_r [35]),
    .ZN(_07857_));
 NAND3_X1 _33344_ (.A1(_07857_),
    .A2(_07331_),
    .A3(_07338_),
    .ZN(_07858_));
 XOR2_X1 _33345_ (.A(net1353),
    .B(\icache.tag_tv_r [38]),
    .Z(_07859_));
 NOR3_X1 _33346_ (.A1(_07858_),
    .A2(_07308_),
    .A3(_07859_),
    .ZN(_07860_));
 XNOR2_X1 _33347_ (.A(_07113_),
    .B(\icache.tag_tv_r [33]),
    .ZN(_07861_));
 AND3_X1 _33348_ (.A1(_07861_),
    .A2(_07323_),
    .A3(_07324_),
    .ZN(_07862_));
 XNOR2_X1 _33349_ (.A(_07123_),
    .B(\icache.tag_tv_r [31]),
    .ZN(_07863_));
 AND4_X1 _33350_ (.A1(_07294_),
    .A2(_07862_),
    .A3(_07295_),
    .A4(_07863_),
    .ZN(_07864_));
 OR2_X1 _33351_ (.A1(_07065_),
    .A2(\icache.tag_tv_r [28]),
    .ZN(_07865_));
 AND4_X1 _33352_ (.A1(_07865_),
    .A2(_07286_),
    .A3(_07330_),
    .A4(_07339_),
    .ZN(_07866_));
 XNOR2_X1 _33353_ (.A(_07370_),
    .B(\icache.tag_tv_r [29]),
    .ZN(_07867_));
 AND4_X1 _33354_ (.A1(_07292_),
    .A2(_07866_),
    .A3(_07337_),
    .A4(_07867_),
    .ZN(_07868_));
 NAND4_X2 _33355_ (.A1(_07856_),
    .A2(_07860_),
    .A3(_07864_),
    .A4(_07868_),
    .ZN(_07869_));
 XNOR2_X1 _33356_ (.A(net1327),
    .B(\icache.tag_tv_r [50]),
    .ZN(_07870_));
 NAND4_X1 _33357_ (.A1(_07307_),
    .A2(_07310_),
    .A3(_07313_),
    .A4(_07870_),
    .ZN(_07871_));
 XNOR2_X1 _33358_ (.A(net1335),
    .B(\icache.tag_tv_r [46]),
    .ZN(_07872_));
 NAND4_X1 _33359_ (.A1(_07301_),
    .A2(_07304_),
    .A3(_07305_),
    .A4(_07872_),
    .ZN(_07873_));
 NOR2_X1 _33360_ (.A1(_07871_),
    .A2(_07873_),
    .ZN(_07874_));
 XNOR2_X2 _33361_ (.A(_07160_),
    .B(\icache.tag_tv_r [53]),
    .ZN(_07875_));
 NAND4_X4 _33362_ (.A1(_07874_),
    .A2(_07311_),
    .A3(_07314_),
    .A4(_07875_),
    .ZN(_07876_));
 NOR3_X4 _33363_ (.A1(_07869_),
    .A2(_07333_),
    .A3(_07876_),
    .ZN(_07877_));
 NOR2_X1 _33364_ (.A1(_07853_),
    .A2(_07877_),
    .ZN(_07878_));
 NAND4_X4 _33365_ (.A1(_07770_),
    .A2(_07829_),
    .A3(_07580_),
    .A4(_07878_),
    .ZN(_07879_));
 NOR2_X1 _33366_ (.A1(_07879_),
    .A2(\icache.N8 ),
    .ZN(_07880_));
 INV_X2 _33367_ (.A(_07880_),
    .ZN(_07881_));
 MUX2_X2 _33368_ (.A(_07656_),
    .B(_07881_),
    .S(_07048_),
    .Z(\icache.stat_mem.w_i ));
 INV_X8 _33369_ (.A(_07612_),
    .ZN(_07882_));
 BUF_X8 _33370_ (.A(_07882_),
    .Z(_07883_));
 BUF_X8 _33371_ (.A(_07613_),
    .Z(_07884_));
 NAND2_X1 _33372_ (.A1(_07884_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [21]),
    .ZN(_07885_));
 BUF_X8 _33373_ (.A(_07624_),
    .Z(_07886_));
 NAND2_X1 _33374_ (.A1(_07886_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [74]),
    .ZN(_07887_));
 AND2_X4 _33375_ (.A1(_07885_),
    .A2(_07887_),
    .ZN(_07888_));
 AND2_X4 _33376_ (.A1(_07604_),
    .A2(_07605_),
    .ZN(_07889_));
 INV_X1 _33377_ (.A(_07889_),
    .ZN(_07890_));
 BUF_X8 _33378_ (.A(_07890_),
    .Z(_07891_));
 BUF_X16 _33379_ (.A(_07891_),
    .Z(_07892_));
 BUF_X8 _33380_ (.A(_07892_),
    .Z(_07893_));
 BUF_X8 _33381_ (.A(_07616_),
    .Z(_07894_));
 BUF_X8 _33382_ (.A(_07894_),
    .Z(_07895_));
 NOR4_X4 _33383_ (.A1(_07883_),
    .A2(_07888_),
    .A3(_07893_),
    .A4(_07895_),
    .ZN(\icache.tag_mem.data_i [0]));
 BUF_X8 _33384_ (.A(_07889_),
    .Z(_07896_));
 BUF_X8 _33385_ (.A(_07896_),
    .Z(_07897_));
 NOR2_X4 _33386_ (.A1(_07882_),
    .A2(_07894_),
    .ZN(_07898_));
 BUF_X8 _33387_ (.A(_07898_),
    .Z(_07899_));
 BUF_X8 _33388_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.head_r ),
    .Z(_07900_));
 OR2_X2 _33389_ (.A1(_07900_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [22]),
    .ZN(_07901_));
 OR2_X2 _33390_ (.A1(_07622_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [75]),
    .ZN(_07902_));
 AND4_X4 _33391_ (.A1(_07897_),
    .A2(_07899_),
    .A3(_07901_),
    .A4(_07902_),
    .ZN(\icache.tag_mem.data_i [117]));
 NAND2_X1 _33392_ (.A1(_07884_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [23]),
    .ZN(_07903_));
 NAND2_X1 _33393_ (.A1(_07886_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [76]),
    .ZN(_07904_));
 AND2_X4 _33394_ (.A1(_07903_),
    .A2(_07904_),
    .ZN(_07905_));
 NOR4_X4 _33395_ (.A1(_07883_),
    .A2(_07905_),
    .A3(_07893_),
    .A4(_07895_),
    .ZN(\icache.tag_mem.data_i [118]));
 BUF_X4 _33396_ (.A(_07624_),
    .Z(_07906_));
 OR2_X2 _33397_ (.A1(_07906_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [24]),
    .ZN(_07907_));
 OR2_X2 _33398_ (.A1(_07622_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [77]),
    .ZN(_07908_));
 AND4_X4 _33399_ (.A1(_07897_),
    .A2(_07899_),
    .A3(_07907_),
    .A4(_07908_),
    .ZN(\icache.tag_mem.data_i [119]));
 OR2_X2 _33400_ (.A1(_07906_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [25]),
    .ZN(_07909_));
 OR2_X2 _33401_ (.A1(_07622_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [78]),
    .ZN(_07910_));
 AND4_X4 _33402_ (.A1(_07897_),
    .A2(_07899_),
    .A3(_07909_),
    .A4(_07910_),
    .ZN(\icache.tag_mem.data_i [120]));
 OR2_X2 _33403_ (.A1(_07906_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [26]),
    .ZN(_07911_));
 OR2_X2 _33404_ (.A1(_07622_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [79]),
    .ZN(_07912_));
 AND4_X4 _33405_ (.A1(_07897_),
    .A2(_07899_),
    .A3(_07911_),
    .A4(_07912_),
    .ZN(\icache.tag_mem.data_i [121]));
 BUF_X8 _33406_ (.A(_07613_),
    .Z(_07913_));
 NAND2_X1 _33407_ (.A1(_07913_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [27]),
    .ZN(_07914_));
 NAND2_X1 _33408_ (.A1(_07886_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [80]),
    .ZN(_07915_));
 AND2_X4 _33409_ (.A1(_07914_),
    .A2(_07915_),
    .ZN(_07916_));
 NOR4_X4 _33410_ (.A1(_07883_),
    .A2(_07916_),
    .A3(_07893_),
    .A4(_07895_),
    .ZN(\icache.tag_mem.data_i [122]));
 NAND2_X1 _33411_ (.A1(_07913_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [28]),
    .ZN(_07917_));
 NAND2_X1 _33412_ (.A1(_07886_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [81]),
    .ZN(_07918_));
 AND2_X4 _33413_ (.A1(_07917_),
    .A2(_07918_),
    .ZN(_07919_));
 NOR4_X4 _33414_ (.A1(_07883_),
    .A2(_07919_),
    .A3(_07893_),
    .A4(_07895_),
    .ZN(\icache.tag_mem.data_i [123]));
 OR2_X1 _33415_ (.A1(_07906_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [29]),
    .ZN(_07920_));
 OR2_X1 _33416_ (.A1(_07622_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [82]),
    .ZN(_07921_));
 AND4_X4 _33417_ (.A1(_07897_),
    .A2(_07899_),
    .A3(_07920_),
    .A4(_07921_),
    .ZN(\icache.tag_mem.data_i [124]));
 OR2_X1 _33418_ (.A1(_07906_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [30]),
    .ZN(_07922_));
 OR2_X2 _33419_ (.A1(_07622_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [83]),
    .ZN(_07923_));
 AND4_X4 _33420_ (.A1(_07897_),
    .A2(_07899_),
    .A3(_07922_),
    .A4(_07923_),
    .ZN(\icache.tag_mem.data_i [125]));
 NAND2_X1 _33421_ (.A1(_07913_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [31]),
    .ZN(_07924_));
 NAND2_X1 _33422_ (.A1(_07886_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [84]),
    .ZN(_07925_));
 AND2_X4 _33423_ (.A1(_07924_),
    .A2(_07925_),
    .ZN(_07926_));
 NOR4_X4 _33424_ (.A1(_07883_),
    .A2(_07926_),
    .A3(_07893_),
    .A4(_07895_),
    .ZN(\icache.tag_mem.data_i [10]));
 OR2_X1 _33425_ (.A1(_07906_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [32]),
    .ZN(_07927_));
 OR2_X2 _33426_ (.A1(_07629_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [85]),
    .ZN(_07928_));
 AND4_X4 _33427_ (.A1(_07897_),
    .A2(_07899_),
    .A3(_07927_),
    .A4(_07928_),
    .ZN(\icache.tag_mem.data_i [11]));
 OR2_X2 _33428_ (.A1(_07906_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [33]),
    .ZN(_07929_));
 OR2_X2 _33429_ (.A1(_07629_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [86]),
    .ZN(_07930_));
 AND4_X4 _33430_ (.A1(_07897_),
    .A2(_07899_),
    .A3(_07929_),
    .A4(_07930_),
    .ZN(\icache.tag_mem.data_i [128]));
 NAND2_X1 _33431_ (.A1(_07913_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [34]),
    .ZN(_07931_));
 NAND2_X1 _33432_ (.A1(_07886_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [87]),
    .ZN(_07932_));
 AND2_X4 _33433_ (.A1(_07931_),
    .A2(_07932_),
    .ZN(_07933_));
 NOR4_X4 _33434_ (.A1(_07883_),
    .A2(_07933_),
    .A3(_07893_),
    .A4(_07895_),
    .ZN(\icache.tag_mem.data_i [100]));
 NAND2_X1 _33435_ (.A1(_07913_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [35]),
    .ZN(_07934_));
 NAND2_X1 _33436_ (.A1(_07900_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [88]),
    .ZN(_07935_));
 AND2_X4 _33437_ (.A1(_07934_),
    .A2(_07935_),
    .ZN(_07936_));
 NOR4_X4 _33438_ (.A1(_07883_),
    .A2(_07936_),
    .A3(_07893_),
    .A4(_07895_),
    .ZN(\icache.tag_mem.data_i [101]));
 OR2_X2 _33439_ (.A1(_07906_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [36]),
    .ZN(_07937_));
 OR2_X2 _33440_ (.A1(_07629_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [89]),
    .ZN(_07938_));
 AND4_X4 _33441_ (.A1(_07897_),
    .A2(_07899_),
    .A3(_07937_),
    .A4(_07938_),
    .ZN(\icache.tag_mem.data_i [102]));
 BUF_X8 _33442_ (.A(_07896_),
    .Z(_07939_));
 OR2_X2 _33443_ (.A1(_07906_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [37]),
    .ZN(_07940_));
 OR2_X2 _33444_ (.A1(_07629_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [90]),
    .ZN(_07941_));
 AND4_X4 _33445_ (.A1(_07939_),
    .A2(_07899_),
    .A3(_07940_),
    .A4(_07941_),
    .ZN(\icache.tag_mem.data_i [103]));
 NAND2_X1 _33446_ (.A1(_07913_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [38]),
    .ZN(_07942_));
 NAND2_X1 _33447_ (.A1(_07900_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [91]),
    .ZN(_07943_));
 AND2_X4 _33448_ (.A1(_07942_),
    .A2(_07943_),
    .ZN(_07944_));
 NOR4_X4 _33449_ (.A1(_07883_),
    .A2(_07944_),
    .A3(_07893_),
    .A4(_07895_),
    .ZN(\icache.tag_mem.data_i [104]));
 OR2_X2 _33450_ (.A1(_07906_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [39]),
    .ZN(_07945_));
 OR2_X2 _33451_ (.A1(_07629_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [92]),
    .ZN(_07946_));
 AND4_X4 _33452_ (.A1(_07939_),
    .A2(_07898_),
    .A3(_07945_),
    .A4(_07946_),
    .ZN(\icache.tag_mem.data_i [105]));
 NAND2_X1 _33453_ (.A1(_07913_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [40]),
    .ZN(_07947_));
 NAND2_X1 _33454_ (.A1(_07900_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [93]),
    .ZN(_07948_));
 AND2_X4 _33455_ (.A1(_07947_),
    .A2(_07948_),
    .ZN(_07949_));
 NOR4_X4 _33456_ (.A1(_07883_),
    .A2(_07949_),
    .A3(_07893_),
    .A4(_07895_),
    .ZN(\icache.tag_mem.data_i [106]));
 NAND2_X1 _33457_ (.A1(_07913_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [41]),
    .ZN(_07950_));
 NAND2_X1 _33458_ (.A1(_07900_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [94]),
    .ZN(_07951_));
 AND2_X4 _33459_ (.A1(_07950_),
    .A2(_07951_),
    .ZN(_07952_));
 NOR4_X4 _33460_ (.A1(_07883_),
    .A2(_07952_),
    .A3(_07893_),
    .A4(_07895_),
    .ZN(\icache.tag_mem.data_i [107]));
 NAND2_X1 _33461_ (.A1(_07913_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [42]),
    .ZN(_07953_));
 NAND2_X1 _33462_ (.A1(_07900_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [95]),
    .ZN(_07954_));
 AND2_X4 _33463_ (.A1(_07953_),
    .A2(_07954_),
    .ZN(_07955_));
 NOR4_X4 _33464_ (.A1(_07882_),
    .A2(_07955_),
    .A3(_07892_),
    .A4(_07894_),
    .ZN(\icache.tag_mem.data_i [108]));
 NAND2_X1 _33465_ (.A1(_07913_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [43]),
    .ZN(_07956_));
 NAND2_X1 _33466_ (.A1(_07900_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [96]),
    .ZN(_07957_));
 AND2_X4 _33467_ (.A1(_07956_),
    .A2(_07957_),
    .ZN(_07958_));
 NOR4_X4 _33468_ (.A1(_07882_),
    .A2(_07958_),
    .A3(_07892_),
    .A4(_07894_),
    .ZN(\icache.tag_mem.data_i [109]));
 NAND2_X1 _33469_ (.A1(_07622_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [44]),
    .ZN(_07959_));
 NAND2_X1 _33470_ (.A1(_07900_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [97]),
    .ZN(_07960_));
 AND2_X4 _33471_ (.A1(_07959_),
    .A2(_07960_),
    .ZN(_07961_));
 NOR4_X4 _33472_ (.A1(_07882_),
    .A2(_07961_),
    .A3(_07892_),
    .A4(_07894_),
    .ZN(\icache.tag_mem.data_i [110]));
 OR2_X2 _33473_ (.A1(_07624_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [45]),
    .ZN(_07962_));
 OR2_X2 _33474_ (.A1(_07629_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [98]),
    .ZN(_07963_));
 AND4_X4 _33475_ (.A1(_07939_),
    .A2(_07898_),
    .A3(_07962_),
    .A4(_07963_),
    .ZN(\icache.tag_mem.data_i [111]));
 NAND2_X1 _33476_ (.A1(_07622_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [46]),
    .ZN(_07964_));
 NAND2_X1 _33477_ (.A1(_07900_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [99]),
    .ZN(_07965_));
 AND2_X4 _33478_ (.A1(_07964_),
    .A2(_07965_),
    .ZN(_07966_));
 NOR4_X4 _33479_ (.A1(_07882_),
    .A2(_07966_),
    .A3(_07892_),
    .A4(_07894_),
    .ZN(\icache.tag_mem.data_i [112]));
 NAND2_X1 _33480_ (.A1(_07622_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [47]),
    .ZN(_07967_));
 NAND2_X1 _33481_ (.A1(_07900_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [100]),
    .ZN(_07968_));
 AND2_X4 _33482_ (.A1(_07967_),
    .A2(_07968_),
    .ZN(_07969_));
 NOR4_X4 _33483_ (.A1(_07882_),
    .A2(_07969_),
    .A3(_07892_),
    .A4(_07894_),
    .ZN(\icache.tag_mem.data_i [113]));
 INV_X1 _33484_ (.A(_07894_),
    .ZN(_07970_));
 BUF_X4 _33485_ (.A(_07889_),
    .Z(_07971_));
 BUF_X8 _33486_ (.A(_07971_),
    .Z(_07972_));
 BUF_X16 _33487_ (.A(_07624_),
    .Z(_07973_));
 MUX2_X2 _33488_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [4]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [57]),
    .S(_07973_),
    .Z(_07974_));
 AND4_X4 _33489_ (.A1(_07612_),
    .A2(_07970_),
    .A3(_07972_),
    .A4(_07974_),
    .ZN(\icache.tag_mem.data_i [114]));
 MUX2_X2 _33490_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [5]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [58]),
    .S(_07973_),
    .Z(_07975_));
 AND4_X4 _33491_ (.A1(_07612_),
    .A2(_07970_),
    .A3(_07972_),
    .A4(_07975_),
    .ZN(\icache.tag_mem.data_i [115]));
 AND2_X2 _33492_ (.A1(_07612_),
    .A2(_07894_),
    .ZN(_07976_));
 NAND2_X4 _33493_ (.A1(_07619_),
    .A2(_07620_),
    .ZN(_07977_));
 INV_X4 _33494_ (.A(_07977_),
    .ZN(_07978_));
 AND2_X4 _33495_ (.A1(_07976_),
    .A2(_07978_),
    .ZN(_07979_));
 AND2_X4 _33496_ (.A1(_07979_),
    .A2(_07889_),
    .ZN(_07980_));
 BUF_X32 _33497_ (.A(_07980_),
    .Z(_07981_));
 AND2_X4 _33498_ (.A1(_07898_),
    .A2(_07889_),
    .ZN(_07982_));
 OR2_X2 _33499_ (.A1(_07981_),
    .A2(_07982_),
    .ZN(_07983_));
 BUF_X16 _33500_ (.A(_07983_),
    .Z(_07984_));
 NAND2_X1 _33501_ (.A1(_07613_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [8]),
    .ZN(_07985_));
 NAND2_X1 _33502_ (.A1(\icache.lce.lce_cmd_inst.rv_adapter.head_r ),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [61]),
    .ZN(_07986_));
 NAND2_X4 _33503_ (.A1(_07985_),
    .A2(_07986_),
    .ZN(_07987_));
 AND2_X2 _33504_ (.A1(_07984_),
    .A2(_07987_),
    .ZN(_07988_));
 NAND2_X1 _33505_ (.A1(_07613_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [7]),
    .ZN(_07989_));
 NAND2_X1 _33506_ (.A1(\icache.lce.lce_cmd_inst.rv_adapter.head_r ),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [60]),
    .ZN(_07990_));
 NAND2_X4 _33507_ (.A1(_07989_),
    .A2(_07990_),
    .ZN(_07991_));
 AND2_X4 _33508_ (.A1(_07983_),
    .A2(_07991_),
    .ZN(_07992_));
 NAND2_X1 _33509_ (.A1(_07613_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [6]),
    .ZN(_07993_));
 NAND2_X1 _33510_ (.A1(\icache.lce.lce_cmd_inst.rv_adapter.head_r ),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [59]),
    .ZN(_07994_));
 NAND2_X4 _33511_ (.A1(_07993_),
    .A2(_07994_),
    .ZN(_07995_));
 AND2_X4 _33512_ (.A1(_07984_),
    .A2(_07995_),
    .ZN(_07996_));
 NOR3_X4 _33513_ (.A1(_07988_),
    .A2(_07992_),
    .A3(_07996_),
    .ZN(\icache.tag_mem.w_mask_i [27]));
 NOR4_X4 _33514_ (.A1(net989),
    .A2(_07882_),
    .A3(_07894_),
    .A4(_07892_),
    .ZN(_07997_));
 NOR2_X4 _33515_ (.A1(net958),
    .A2(_07981_),
    .ZN(\icache.tag_mem.w_mask_i [0]));
 INV_X2 _33516_ (.A(_07988_),
    .ZN(_07998_));
 INV_X2 _33517_ (.A(_07992_),
    .ZN(_07999_));
 NAND3_X4 _33518_ (.A1(_07998_),
    .A2(_07999_),
    .A3(_07996_),
    .ZN(_08000_));
 AOI21_X4 _33519_ (.A(_07981_),
    .B1(_08000_),
    .B2(_07982_),
    .ZN(\icache.tag_mem.w_mask_i [29]));
 NAND2_X4 _33520_ (.A1(_08000_),
    .A2(_07984_),
    .ZN(\icache.tag_mem.w_mask_i [56]));
 INV_X2 _33521_ (.A(_07995_),
    .ZN(_08001_));
 NAND3_X4 _33522_ (.A1(_07998_),
    .A2(_07992_),
    .A3(_08001_),
    .ZN(_08002_));
 AOI21_X4 _33523_ (.A(_07981_),
    .B1(_08002_),
    .B2(_07982_),
    .ZN(\icache.tag_mem.w_mask_i [58]));
 NAND2_X4 _33524_ (.A1(_08002_),
    .A2(_07984_),
    .ZN(\icache.tag_mem.w_mask_i [85]));
 NAND3_X4 _33525_ (.A1(_07998_),
    .A2(_07992_),
    .A3(_07996_),
    .ZN(_08003_));
 AOI21_X4 _33526_ (.A(_07981_),
    .B1(_08003_),
    .B2(_07982_),
    .ZN(\icache.tag_mem.w_mask_i [100]));
 NAND2_X4 _33527_ (.A1(_08003_),
    .A2(_07984_),
    .ZN(\icache.tag_mem.w_mask_i [114]));
 INV_X1 _33528_ (.A(_07996_),
    .ZN(_08004_));
 NAND3_X4 _33529_ (.A1(_07999_),
    .A2(_08004_),
    .A3(_07988_),
    .ZN(_08005_));
 AOI21_X4 _33530_ (.A(_07981_),
    .B1(_08005_),
    .B2(_07982_),
    .ZN(\icache.tag_mem.w_mask_i [116]));
 NAND2_X4 _33531_ (.A1(_08005_),
    .A2(_07984_),
    .ZN(\icache.tag_mem.w_mask_i [143]));
 NAND3_X4 _33532_ (.A1(_07999_),
    .A2(_07987_),
    .A3(_07996_),
    .ZN(_08006_));
 AOI21_X4 _33533_ (.A(_07981_),
    .B1(_08006_),
    .B2(_07982_),
    .ZN(\icache.tag_mem.w_mask_i [145]));
 NAND2_X4 _33534_ (.A1(_08006_),
    .A2(_07984_),
    .ZN(\icache.tag_mem.w_mask_i [172]));
 NAND3_X4 _33535_ (.A1(_07992_),
    .A2(_07987_),
    .A3(_08001_),
    .ZN(_08007_));
 AOI21_X4 _33536_ (.A(_07981_),
    .B1(_08007_),
    .B2(_07982_),
    .ZN(\icache.tag_mem.w_mask_i [174]));
 NAND2_X4 _33537_ (.A1(_08007_),
    .A2(_07984_),
    .ZN(\icache.tag_mem.w_mask_i [201]));
 NAND3_X4 _33538_ (.A1(_07996_),
    .A2(_07987_),
    .A3(_07991_),
    .ZN(_08008_));
 AOI21_X4 _33539_ (.A(_07981_),
    .B1(_08008_),
    .B2(_07982_),
    .ZN(\icache.tag_mem.w_mask_i [203]));
 NAND2_X4 _33540_ (.A1(_08008_),
    .A2(_07984_),
    .ZN(\icache.tag_mem.w_mask_i [230]));
 NOR2_X4 _33541_ (.A1(\icache.lce.lce_cmd_inst.state_r [1]),
    .A2(_07605_),
    .ZN(_08009_));
 NAND2_X1 _33542_ (.A1(_08009_),
    .A2(\icache.N7 ),
    .ZN(_08010_));
 INV_X1 _33543_ (.A(freeze_i),
    .ZN(_08011_));
 NAND3_X1 _33544_ (.A1(\icache.N10 ),
    .A2(\icache.N8 ),
    .A3(_00003_),
    .ZN(_08012_));
 AND2_X1 _33545_ (.A1(_07881_),
    .A2(_08012_),
    .ZN(_08013_));
 NOR2_X2 _33546_ (.A1(\icache.lce.lce_req_inst.state_r [2]),
    .A2(\icache.lce.lce_req_inst.state_r [1]),
    .ZN(_08014_));
 INV_X1 _33547_ (.A(\icache.lce.lce_req_inst.state_r [0]),
    .ZN(_08015_));
 AND2_X4 _33548_ (.A1(_08014_),
    .A2(_08015_),
    .ZN(_08016_));
 AND2_X2 _33549_ (.A1(_08013_),
    .A2(_08016_),
    .ZN(_08017_));
 INV_X1 _33550_ (.A(_00002_),
    .ZN(_08018_));
 AND2_X1 _33551_ (.A1(_08014_),
    .A2(_08018_),
    .ZN(_08019_));
 INV_X1 _33552_ (.A(\icache.lce.lce_req_inst.state_r [2]),
    .ZN(_08020_));
 NOR2_X2 _33553_ (.A1(_08020_),
    .A2(\icache.lce.lce_req_inst.state_r [1]),
    .ZN(_08021_));
 INV_X1 _33554_ (.A(\icache.lce.lce_req_inst.state_r [1]),
    .ZN(_08022_));
 NOR2_X4 _33555_ (.A1(_08022_),
    .A2(\icache.lce.lce_req_inst.state_r [2]),
    .ZN(_08023_));
 NOR4_X4 _33556_ (.A1(_08016_),
    .A2(_08019_),
    .A3(_08021_),
    .A4(_08023_),
    .ZN(_08024_));
 OAI221_X2 _33557_ (.A(_08010_),
    .B1(_08011_),
    .B2(\icache.N7 ),
    .C1(_08017_),
    .C2(_08024_),
    .ZN(_08025_));
 BUF_X16 _33558_ (.A(_08025_),
    .Z(_08026_));
 INV_X1 _33559_ (.A(fe_cmd_i[75]),
    .ZN(_08027_));
 NOR2_X1 _33560_ (.A1(_08027_),
    .A2(fe_cmd_i[74]),
    .ZN(_08028_));
 AND3_X2 _33561_ (.A1(_08028_),
    .A2(fe_cmd_v_i),
    .A3(fe_cmd_i[73]),
    .ZN(_08029_));
 AND2_X1 _33562_ (.A1(_08029_),
    .A2(_00004_),
    .ZN(_08030_));
 BUF_X8 _33563_ (.A(_08030_),
    .Z(_08031_));
 INV_X4 _33564_ (.A(_08031_),
    .ZN(_08032_));
 NOR2_X1 _33565_ (.A1(\bp_fe_pc_gen_1.state_r [0]),
    .A2(\bp_fe_pc_gen_1.state_r [1]),
    .ZN(_08033_));
 INV_X1 _33566_ (.A(_08033_),
    .ZN(_08034_));
 NAND3_X4 _33567_ (.A1(_08032_),
    .A2(fe_queue_ready_i),
    .A3(_08034_),
    .ZN(_08035_));
 NOR2_X4 _33568_ (.A1(_08026_),
    .A2(_08035_),
    .ZN(_08036_));
 BUF_X16 _33569_ (.A(_08036_),
    .Z(_08037_));
 BUF_X16 _33570_ (.A(_08037_),
    .Z(_08038_));
 XOR2_X2 _33571_ (.A(\bp_fe_pc_gen_1.btb.r_tag_r [2]),
    .B(net1401),
    .Z(_08039_));
 INV_X1 _33572_ (.A(\bp_fe_pc_gen_1.btb.r_tag_r [5]),
    .ZN(_08040_));
 INV_X1 _33573_ (.A(net1398),
    .ZN(_08041_));
 AOI22_X1 _33574_ (.A1(_08040_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.data_o [44]),
    .B1(_08041_),
    .B2(\bp_fe_pc_gen_1.btb.r_tag_r [7]),
    .ZN(_08042_));
 INV_X2 _33575_ (.A(net1400),
    .ZN(_08043_));
 OR2_X1 _33576_ (.A1(_08043_),
    .A2(\bp_fe_pc_gen_1.btb.r_tag_r [3]),
    .ZN(_08044_));
 OAI211_X1 _33577_ (.A(_08042_),
    .B(_08044_),
    .C1(_08040_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.data_o [44]),
    .ZN(_08045_));
 INV_X2 _33578_ (.A(\bp_fe_pc_gen_1.btb.r_tag_r [0]),
    .ZN(_08046_));
 AOI211_X1 _33579_ (.A(_08039_),
    .B(_08045_),
    .C1(_08046_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.data_o [39]),
    .ZN(_08047_));
 NOR3_X4 _33580_ (.A1(\bp_fe_pc_gen_1.btb.r_idx_r [2]),
    .A2(\bp_fe_pc_gen_1.btb.r_idx_r [0]),
    .A3(\bp_fe_pc_gen_1.btb.r_idx_r [1]),
    .ZN(_08048_));
 INV_X1 _33581_ (.A(\bp_fe_pc_gen_1.btb.r_idx_r [4]),
    .ZN(_08049_));
 BUF_X2 _33582_ (.A(_08049_),
    .Z(_08050_));
 BUF_X4 _33583_ (.A(_08050_),
    .Z(_08051_));
 INV_X1 _33584_ (.A(\bp_fe_pc_gen_1.btb.r_idx_r [3]),
    .ZN(_08052_));
 BUF_X4 _33585_ (.A(_08052_),
    .Z(_08053_));
 AND3_X4 _33586_ (.A1(_08048_),
    .A2(_08051_),
    .A3(_08053_),
    .ZN(_08054_));
 BUF_X4 _33587_ (.A(_00072_),
    .Z(_08055_));
 BUF_X4 _33588_ (.A(_08055_),
    .Z(_08056_));
 BUF_X2 _33589_ (.A(_08056_),
    .Z(_08057_));
 BUF_X4 _33590_ (.A(_08057_),
    .Z(_08058_));
 NAND3_X4 _33591_ (.A1(_08054_),
    .A2(_08058_),
    .A3(_00006_),
    .ZN(_08059_));
 NOR2_X1 _33592_ (.A1(_08046_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.data_o [39]),
    .ZN(_08060_));
 INV_X1 _33593_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.data_o [40]),
    .ZN(_08061_));
 AOI21_X1 _33594_ (.A(_08060_),
    .B1(\bp_fe_pc_gen_1.btb.r_tag_r [1]),
    .B2(_08061_),
    .ZN(_08062_));
 NAND2_X1 _33595_ (.A1(_08043_),
    .A2(\bp_fe_pc_gen_1.btb.r_tag_r [3]),
    .ZN(_08063_));
 OAI211_X1 _33596_ (.A(_08062_),
    .B(_08063_),
    .C1(\bp_fe_pc_gen_1.btb.r_tag_r [1]),
    .C2(_08061_),
    .ZN(_08064_));
 XOR2_X1 _33597_ (.A(\bp_fe_pc_gen_1.btb.r_tag_r [6]),
    .B(net1399),
    .Z(_08065_));
 XOR2_X1 _33598_ (.A(\bp_fe_pc_gen_1.btb.r_tag_r [4]),
    .B(\bp_fe_pc_gen_1.btb.tag_mem.data_o [43]),
    .Z(_08066_));
 NOR3_X1 _33599_ (.A1(_08064_),
    .A2(_08065_),
    .A3(_08066_),
    .ZN(_08067_));
 XOR2_X2 _33600_ (.A(\bp_fe_pc_gen_1.btb.r_tag_r [8]),
    .B(\bp_fe_pc_gen_1.btb.tag_mem.data_o [47]),
    .Z(_08068_));
 INV_X1 _33601_ (.A(\bp_fe_pc_gen_1.btb.r_tag_r [9]),
    .ZN(_08069_));
 OAI22_X1 _33602_ (.A1(\bp_fe_pc_gen_1.btb.r_tag_r [7]),
    .A2(_08041_),
    .B1(_08069_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.data_o [48]),
    .ZN(_08070_));
 AND2_X1 _33603_ (.A1(_08069_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.data_o [48]),
    .ZN(_08071_));
 INV_X1 _33604_ (.A(\bp_fe_pc_gen_1.btb.r_v_r ),
    .ZN(_08072_));
 NOR4_X2 _33605_ (.A1(_08068_),
    .A2(_08070_),
    .A3(_08071_),
    .A4(_08072_),
    .ZN(_08073_));
 NAND4_X2 _33606_ (.A1(_08047_),
    .A2(_08059_),
    .A3(_08067_),
    .A4(_08073_),
    .ZN(_08074_));
 INV_X2 _33607_ (.A(\bp_fe_pc_gen_1.btb.r_idx_r [1]),
    .ZN(_08075_));
 NOR3_X4 _33608_ (.A1(_08075_),
    .A2(\bp_fe_pc_gen_1.btb.r_idx_r [2]),
    .A3(\bp_fe_pc_gen_1.btb.r_idx_r [0]),
    .ZN(_08076_));
 AND3_X2 _33609_ (.A1(_08076_),
    .A2(_08051_),
    .A3(_08053_),
    .ZN(_08077_));
 NAND3_X1 _33610_ (.A1(_08077_),
    .A2(_08058_),
    .A3(_00008_),
    .ZN(_08078_));
 AND2_X1 _33611_ (.A1(\bp_fe_pc_gen_1.btb.r_idx_r [0]),
    .A2(\bp_fe_pc_gen_1.btb.r_idx_r [1]),
    .ZN(_08079_));
 INV_X1 _33612_ (.A(_00071_),
    .ZN(_08080_));
 AND3_X2 _33613_ (.A1(_08079_),
    .A2(_08052_),
    .A3(_08080_),
    .ZN(_08081_));
 INV_X1 _33614_ (.A(_08081_),
    .ZN(_08082_));
 INV_X4 _33615_ (.A(_00072_),
    .ZN(_08083_));
 NOR4_X1 _33616_ (.A1(_08082_),
    .A2(\bp_fe_pc_gen_1.btb.r_idx_r [4]),
    .A3(_08083_),
    .A4(_00013_),
    .ZN(_08084_));
 NOR3_X4 _33617_ (.A1(_08075_),
    .A2(\bp_fe_pc_gen_1.btb.r_idx_r [0]),
    .A3(_00071_),
    .ZN(_08085_));
 AND3_X2 _33618_ (.A1(_08085_),
    .A2(_08050_),
    .A3(_08053_),
    .ZN(_08086_));
 AOI21_X1 _33619_ (.A(_08084_),
    .B1(_08058_),
    .B2(_08086_),
    .ZN(_08087_));
 INV_X2 _33620_ (.A(\bp_fe_pc_gen_1.btb.r_idx_r [2]),
    .ZN(_08088_));
 NAND3_X4 _33621_ (.A1(_08088_),
    .A2(_08075_),
    .A3(\bp_fe_pc_gen_1.btb.r_idx_r [0]),
    .ZN(_08089_));
 NOR3_X2 _33622_ (.A1(_08089_),
    .A2(\bp_fe_pc_gen_1.btb.r_idx_r [4]),
    .A3(_00070_),
    .ZN(_08090_));
 AND2_X1 _33623_ (.A1(_08090_),
    .A2(_08057_),
    .ZN(_08091_));
 INV_X1 _33624_ (.A(_08091_),
    .ZN(_08092_));
 NOR2_X1 _33625_ (.A1(_08092_),
    .A2(_00015_),
    .ZN(_08093_));
 NOR2_X1 _33626_ (.A1(\bp_fe_pc_gen_1.btb.r_idx_r [0]),
    .A2(\bp_fe_pc_gen_1.btb.r_idx_r [1]),
    .ZN(_08094_));
 INV_X1 _33627_ (.A(_00070_),
    .ZN(_08095_));
 BUF_X4 _33628_ (.A(_08095_),
    .Z(_08096_));
 AND3_X2 _33629_ (.A1(_08094_),
    .A2(_08088_),
    .A3(_08096_),
    .ZN(_08097_));
 AND3_X1 _33630_ (.A1(_08097_),
    .A2(_08051_),
    .A3(_08057_),
    .ZN(_08098_));
 OR2_X1 _33631_ (.A1(_08093_),
    .A2(_08098_),
    .ZN(_08099_));
 AND3_X1 _33632_ (.A1(_08076_),
    .A2(_08050_),
    .A3(_08096_),
    .ZN(_08100_));
 AND3_X1 _33633_ (.A1(_08100_),
    .A2(_08057_),
    .A3(_00016_),
    .ZN(_08101_));
 NOR3_X4 _33634_ (.A1(\bp_fe_pc_gen_1.btb.r_idx_r [0]),
    .A2(\bp_fe_pc_gen_1.btb.r_idx_r [1]),
    .A3(_00071_),
    .ZN(_08102_));
 AND3_X1 _33635_ (.A1(_08102_),
    .A2(_08050_),
    .A3(_08096_),
    .ZN(_08103_));
 NAND3_X1 _33636_ (.A1(_08103_),
    .A2(_08057_),
    .A3(_00018_),
    .ZN(_08104_));
 AND3_X2 _33637_ (.A1(_08075_),
    .A2(_08080_),
    .A3(\bp_fe_pc_gen_1.btb.r_idx_r [0]),
    .ZN(_08105_));
 AND3_X1 _33638_ (.A1(_08105_),
    .A2(_08050_),
    .A3(_08096_),
    .ZN(_08106_));
 AND2_X1 _33639_ (.A1(_08106_),
    .A2(_08056_),
    .ZN(_08107_));
 INV_X1 _33640_ (.A(_08107_),
    .ZN(_08108_));
 AND3_X2 _33641_ (.A1(_08085_),
    .A2(_08050_),
    .A3(_08096_),
    .ZN(_08109_));
 NAND3_X1 _33642_ (.A1(_08109_),
    .A2(_08056_),
    .A3(_00020_),
    .ZN(_08110_));
 NAND2_X1 _33643_ (.A1(_08108_),
    .A2(_08110_),
    .ZN(_08111_));
 NOR3_X2 _33644_ (.A1(_08089_),
    .A2(\bp_fe_pc_gen_1.btb.r_idx_r [3]),
    .A3(_00069_),
    .ZN(_08112_));
 NAND3_X1 _33645_ (.A1(_08112_),
    .A2(_08056_),
    .A3(_00023_),
    .ZN(_08113_));
 INV_X2 _33646_ (.A(_00069_),
    .ZN(_08114_));
 BUF_X2 _33647_ (.A(_08114_),
    .Z(_08115_));
 BUF_X2 _33648_ (.A(_08115_),
    .Z(_08116_));
 AND3_X1 _33649_ (.A1(_08076_),
    .A2(_08053_),
    .A3(_08116_),
    .ZN(_08117_));
 AND2_X1 _33650_ (.A1(_08117_),
    .A2(_08056_),
    .ZN(_08118_));
 NAND3_X4 _33651_ (.A1(_08088_),
    .A2(\bp_fe_pc_gen_1.btb.r_idx_r [0]),
    .A3(\bp_fe_pc_gen_1.btb.r_idx_r [1]),
    .ZN(_08119_));
 NOR2_X4 _33652_ (.A1(_08119_),
    .A2(\bp_fe_pc_gen_1.btb.r_idx_r [3]),
    .ZN(_08120_));
 AND4_X1 _33653_ (.A1(_08116_),
    .A2(_08120_),
    .A3(_08056_),
    .A4(_00025_),
    .ZN(_08121_));
 AND3_X2 _33654_ (.A1(_08080_),
    .A2(\bp_fe_pc_gen_1.btb.r_idx_r [0]),
    .A3(\bp_fe_pc_gen_1.btb.r_idx_r [1]),
    .ZN(_08122_));
 AND3_X2 _33655_ (.A1(_08122_),
    .A2(_08052_),
    .A3(_08115_),
    .ZN(_08123_));
 AND2_X1 _33656_ (.A1(_08123_),
    .A2(_08055_),
    .ZN(_08124_));
 AND3_X2 _33657_ (.A1(_08048_),
    .A2(_08096_),
    .A3(_08115_),
    .ZN(_08125_));
 AND3_X1 _33658_ (.A1(_08125_),
    .A2(_08055_),
    .A3(_00030_),
    .ZN(_08126_));
 NOR2_X4 _33659_ (.A1(_08119_),
    .A2(_00070_),
    .ZN(_08127_));
 NAND2_X1 _33660_ (.A1(_08127_),
    .A2(_08116_),
    .ZN(_08128_));
 NOR3_X1 _33661_ (.A1(_08128_),
    .A2(_08083_),
    .A3(_00033_),
    .ZN(_08129_));
 AND3_X2 _33662_ (.A1(_08094_),
    .A2(_08080_),
    .A3(_08096_),
    .ZN(_08130_));
 AND3_X1 _33663_ (.A1(_08130_),
    .A2(_08116_),
    .A3(_00072_),
    .ZN(_08131_));
 INV_X1 _33664_ (.A(_08131_),
    .ZN(_08132_));
 AND3_X2 _33665_ (.A1(_08085_),
    .A2(_08095_),
    .A3(_08114_),
    .ZN(_08133_));
 AND2_X1 _33666_ (.A1(_08133_),
    .A2(_00072_),
    .ZN(_08134_));
 INV_X1 _33667_ (.A(_08134_),
    .ZN(_08135_));
 NOR2_X1 _33668_ (.A1(_08135_),
    .A2(_00036_),
    .ZN(_08136_));
 AND2_X2 _33669_ (.A1(_08105_),
    .A2(_08095_),
    .ZN(_08137_));
 AND2_X1 _33670_ (.A1(_08137_),
    .A2(_08116_),
    .ZN(_08138_));
 INV_X1 _33671_ (.A(_08054_),
    .ZN(_08139_));
 BUF_X2 _33672_ (.A(\bp_fe_pc_gen_1.btb.r_idx_r [5]),
    .Z(_08140_));
 BUF_X4 _33673_ (.A(_08140_),
    .Z(_08141_));
 INV_X2 _33674_ (.A(_08141_),
    .ZN(_08142_));
 NOR3_X1 _33675_ (.A1(_08139_),
    .A2(_08142_),
    .A3(_00038_),
    .ZN(_08143_));
 AND3_X2 _33676_ (.A1(_08079_),
    .A2(_08080_),
    .A3(_08095_),
    .ZN(_08144_));
 AND3_X1 _33677_ (.A1(_08144_),
    .A2(_08116_),
    .A3(_00072_),
    .ZN(_08145_));
 NOR2_X1 _33678_ (.A1(_08143_),
    .A2(_08145_),
    .ZN(_08146_));
 BUF_X2 _33679_ (.A(_08141_),
    .Z(_08147_));
 BUF_X2 _33680_ (.A(_08147_),
    .Z(_08148_));
 AND3_X1 _33681_ (.A1(_08120_),
    .A2(_08051_),
    .A3(_08148_),
    .ZN(_08149_));
 AOI22_X1 _33682_ (.A1(_08149_),
    .A2(_00041_),
    .B1(_08148_),
    .B2(_08077_),
    .ZN(_08150_));
 AND3_X2 _33683_ (.A1(_08105_),
    .A2(_08050_),
    .A3(_08053_),
    .ZN(_08151_));
 AND3_X1 _33684_ (.A1(_08151_),
    .A2(_08148_),
    .A3(_00043_),
    .ZN(_08152_));
 AND3_X2 _33685_ (.A1(_08102_),
    .A2(_08051_),
    .A3(_08053_),
    .ZN(_08153_));
 AND3_X1 _33686_ (.A1(_08081_),
    .A2(_08050_),
    .A3(_08147_),
    .ZN(_08154_));
 AOI22_X1 _33687_ (.A1(_08154_),
    .A2(_00045_),
    .B1(_08148_),
    .B2(_08086_),
    .ZN(_08155_));
 AND3_X1 _33688_ (.A1(_08090_),
    .A2(_08147_),
    .A3(_00047_),
    .ZN(_08156_));
 AND3_X1 _33689_ (.A1(_08048_),
    .A2(_08050_),
    .A3(_08096_),
    .ZN(_08157_));
 AND2_X1 _33690_ (.A1(_08157_),
    .A2(_08147_),
    .ZN(_08158_));
 OR2_X1 _33691_ (.A1(_08156_),
    .A2(_08158_),
    .ZN(_08159_));
 AND2_X2 _33692_ (.A1(_08076_),
    .A2(_08096_),
    .ZN(_08160_));
 NAND4_X1 _33693_ (.A1(_08160_),
    .A2(_08051_),
    .A3(_08147_),
    .A4(_00048_),
    .ZN(_08161_));
 AND3_X1 _33694_ (.A1(_08106_),
    .A2(_08147_),
    .A3(_00051_),
    .ZN(_08162_));
 AND2_X1 _33695_ (.A1(_08103_),
    .A2(_08141_),
    .ZN(_08163_));
 NOR2_X1 _33696_ (.A1(_08162_),
    .A2(_08163_),
    .ZN(_08164_));
 NAND3_X1 _33697_ (.A1(_08122_),
    .A2(_08049_),
    .A3(_08096_),
    .ZN(_08165_));
 NOR2_X1 _33698_ (.A1(_08165_),
    .A2(_08142_),
    .ZN(_08166_));
 AND2_X1 _33699_ (.A1(_08166_),
    .A2(_00053_),
    .ZN(_08167_));
 NAND3_X1 _33700_ (.A1(_08112_),
    .A2(_08141_),
    .A3(_00055_),
    .ZN(_08168_));
 AND3_X1 _33701_ (.A1(_08048_),
    .A2(_08053_),
    .A3(_08116_),
    .ZN(_08169_));
 NAND2_X1 _33702_ (.A1(_08169_),
    .A2(_08141_),
    .ZN(_08170_));
 AND2_X1 _33703_ (.A1(_08168_),
    .A2(_08170_),
    .ZN(_08171_));
 NOR3_X2 _33704_ (.A1(_08119_),
    .A2(\bp_fe_pc_gen_1.btb.r_idx_r [3]),
    .A3(_00069_),
    .ZN(_08172_));
 NAND2_X1 _33705_ (.A1(_08172_),
    .A2(_08141_),
    .ZN(_08173_));
 AND3_X1 _33706_ (.A1(_08102_),
    .A2(_08053_),
    .A3(_08116_),
    .ZN(_08174_));
 NAND3_X1 _33707_ (.A1(_08174_),
    .A2(_08141_),
    .A3(_00058_),
    .ZN(_08175_));
 AND3_X2 _33708_ (.A1(_08085_),
    .A2(_08052_),
    .A3(_08115_),
    .ZN(_08176_));
 AND3_X1 _33709_ (.A1(_08176_),
    .A2(_08140_),
    .A3(_00060_),
    .ZN(_08177_));
 AND3_X2 _33710_ (.A1(_08105_),
    .A2(_08053_),
    .A3(_08115_),
    .ZN(_08178_));
 NAND3_X1 _33711_ (.A1(_08123_),
    .A2(_08140_),
    .A3(_00061_),
    .ZN(_08179_));
 NOR3_X4 _33712_ (.A1(_08089_),
    .A2(_00070_),
    .A3(_00069_),
    .ZN(_08180_));
 AND3_X1 _33713_ (.A1(_08180_),
    .A2(\bp_fe_pc_gen_1.btb.r_idx_r [5]),
    .A3(_00063_),
    .ZN(_08181_));
 NAND4_X1 _33714_ (.A1(_08144_),
    .A2(_08114_),
    .A3(\bp_fe_pc_gen_1.btb.r_idx_r [5]),
    .A4(\bp_fe_pc_gen_1.btb.v_r [63]),
    .ZN(_08182_));
 NAND2_X1 _33715_ (.A1(_08133_),
    .A2(\bp_fe_pc_gen_1.btb.r_idx_r [5]),
    .ZN(_08183_));
 MUX2_X1 _33716_ (.A(_00068_),
    .B(_08182_),
    .S(_08183_),
    .Z(_08184_));
 NAND3_X1 _33717_ (.A1(_08137_),
    .A2(_08114_),
    .A3(\bp_fe_pc_gen_1.btb.r_idx_r [5]),
    .ZN(_08185_));
 MUX2_X1 _33718_ (.A(_00067_),
    .B(_08184_),
    .S(_08185_),
    .Z(_08186_));
 NAND3_X1 _33719_ (.A1(_08130_),
    .A2(_08115_),
    .A3(\bp_fe_pc_gen_1.btb.r_idx_r [5]),
    .ZN(_08187_));
 MUX2_X1 _33720_ (.A(_00066_),
    .B(_08186_),
    .S(_08187_),
    .Z(_08188_));
 NAND3_X1 _33721_ (.A1(_08127_),
    .A2(_08115_),
    .A3(\bp_fe_pc_gen_1.btb.r_idx_r [5]),
    .ZN(_08189_));
 MUX2_X1 _33722_ (.A(_00065_),
    .B(_08188_),
    .S(_08189_),
    .Z(_08190_));
 AND2_X1 _33723_ (.A1(_08160_),
    .A2(_08115_),
    .ZN(_08191_));
 NAND2_X1 _33724_ (.A1(_08191_),
    .A2(\bp_fe_pc_gen_1.btb.r_idx_r [5]),
    .ZN(_08192_));
 MUX2_X1 _33725_ (.A(_00064_),
    .B(_08190_),
    .S(_08192_),
    .Z(_08193_));
 NOR2_X2 _33726_ (.A1(_08089_),
    .A2(_00070_),
    .ZN(_08194_));
 AND3_X1 _33727_ (.A1(_08194_),
    .A2(_08115_),
    .A3(\bp_fe_pc_gen_1.btb.r_idx_r [5]),
    .ZN(_08195_));
 INV_X1 _33728_ (.A(_08195_),
    .ZN(_08196_));
 AOI221_X1 _33729_ (.A(_08181_),
    .B1(_08140_),
    .B2(_08125_),
    .C1(_08193_),
    .C2(_08196_),
    .ZN(_08197_));
 NAND2_X1 _33730_ (.A1(_08125_),
    .A2(_08140_),
    .ZN(_08198_));
 NOR2_X1 _33731_ (.A1(_08198_),
    .A2(_00062_),
    .ZN(_08199_));
 AND3_X1 _33732_ (.A1(_08081_),
    .A2(_08115_),
    .A3(_08140_),
    .ZN(_08200_));
 OR2_X1 _33733_ (.A1(_08199_),
    .A2(_08200_),
    .ZN(_08201_));
 OAI21_X1 _33734_ (.A(_08179_),
    .B1(_08197_),
    .B2(_08201_),
    .ZN(_08202_));
 NAND2_X1 _33735_ (.A1(_08176_),
    .A2(_08140_),
    .ZN(_08203_));
 AOI221_X2 _33736_ (.A(_08177_),
    .B1(_08140_),
    .B2(_08178_),
    .C1(_08202_),
    .C2(_08203_),
    .ZN(_08204_));
 NAND2_X1 _33737_ (.A1(_08178_),
    .A2(_08140_),
    .ZN(_08205_));
 NOR2_X1 _33738_ (.A1(_08205_),
    .A2(_00059_),
    .ZN(_08206_));
 AND2_X1 _33739_ (.A1(_08174_),
    .A2(_08140_),
    .ZN(_08207_));
 OR2_X1 _33740_ (.A1(_08206_),
    .A2(_08207_),
    .ZN(_08208_));
 OAI211_X1 _33741_ (.A(_08173_),
    .B(_08175_),
    .C1(_08204_),
    .C2(_08208_),
    .ZN(_08209_));
 OR2_X1 _33742_ (.A1(_08173_),
    .A2(_00057_),
    .ZN(_08210_));
 AOI22_X1 _33743_ (.A1(_08209_),
    .A2(_08210_),
    .B1(_08141_),
    .B2(_08117_),
    .ZN(_08211_));
 NAND2_X1 _33744_ (.A1(_08117_),
    .A2(_08141_),
    .ZN(_08212_));
 INV_X1 _33745_ (.A(_08112_),
    .ZN(_08213_));
 OAI22_X1 _33746_ (.A1(_08212_),
    .A2(_00056_),
    .B1(_08142_),
    .B2(_08213_),
    .ZN(_08214_));
 OAI21_X1 _33747_ (.A(_08171_),
    .B1(_08211_),
    .B2(_08214_),
    .ZN(_08215_));
 NOR2_X1 _33748_ (.A1(_08170_),
    .A2(_00054_),
    .ZN(_08216_));
 NOR2_X1 _33749_ (.A1(_08216_),
    .A2(_08166_),
    .ZN(_08217_));
 AOI221_X2 _33750_ (.A(_08167_),
    .B1(_08141_),
    .B2(_08109_),
    .C1(_08215_),
    .C2(_08217_),
    .ZN(_08218_));
 NAND2_X1 _33751_ (.A1(_08106_),
    .A2(_08147_),
    .ZN(_08219_));
 NAND2_X1 _33752_ (.A1(_08109_),
    .A2(_08147_),
    .ZN(_08220_));
 OAI21_X1 _33753_ (.A(_08219_),
    .B1(_08220_),
    .B2(_00052_),
    .ZN(_08221_));
 OAI21_X1 _33754_ (.A(_08164_),
    .B1(_08218_),
    .B2(_08221_),
    .ZN(_08222_));
 INV_X1 _33755_ (.A(_08163_),
    .ZN(_08223_));
 NOR2_X1 _33756_ (.A1(_08223_),
    .A2(_00050_),
    .ZN(_08224_));
 AND3_X1 _33757_ (.A1(_08127_),
    .A2(_08050_),
    .A3(_08147_),
    .ZN(_08225_));
 NOR2_X1 _33758_ (.A1(_08224_),
    .A2(_08225_),
    .ZN(_08226_));
 AOI22_X2 _33759_ (.A1(_08222_),
    .A2(_08226_),
    .B1(_00049_),
    .B2(_08225_),
    .ZN(_08227_));
 AND2_X1 _33760_ (.A1(_08100_),
    .A2(_08147_),
    .ZN(_08228_));
 OAI21_X1 _33761_ (.A(_08161_),
    .B1(_08227_),
    .B2(_08228_),
    .ZN(_08229_));
 NAND3_X1 _33762_ (.A1(_08194_),
    .A2(_08051_),
    .A3(_08148_),
    .ZN(_08230_));
 AOI21_X1 _33763_ (.A(_08159_),
    .B1(_08229_),
    .B2(_08230_),
    .ZN(_08231_));
 INV_X1 _33764_ (.A(_08154_),
    .ZN(_08232_));
 INV_X1 _33765_ (.A(_08158_),
    .ZN(_08233_));
 OAI21_X1 _33766_ (.A(_08232_),
    .B1(_08233_),
    .B2(_00046_),
    .ZN(_08234_));
 OAI21_X1 _33767_ (.A(_08155_),
    .B1(_08231_),
    .B2(_08234_),
    .ZN(_08235_));
 INV_X1 _33768_ (.A(_08086_),
    .ZN(_08236_));
 NOR3_X1 _33769_ (.A1(_08236_),
    .A2(_08142_),
    .A3(_00044_),
    .ZN(_08237_));
 AOI21_X1 _33770_ (.A(_08237_),
    .B1(_08148_),
    .B2(_08151_),
    .ZN(_08238_));
 AOI221_X2 _33771_ (.A(_08152_),
    .B1(_08148_),
    .B2(_08153_),
    .C1(_08235_),
    .C2(_08238_),
    .ZN(_08239_));
 INV_X1 _33772_ (.A(_08149_),
    .ZN(_08240_));
 NAND2_X1 _33773_ (.A1(_08153_),
    .A2(_08148_),
    .ZN(_08241_));
 OAI21_X1 _33774_ (.A(_08240_),
    .B1(_08241_),
    .B2(_00042_),
    .ZN(_08242_));
 OAI21_X1 _33775_ (.A(_08150_),
    .B1(_08239_),
    .B2(_08242_),
    .ZN(_08243_));
 AND2_X1 _33776_ (.A1(_08077_),
    .A2(_08148_),
    .ZN(_08244_));
 INV_X1 _33777_ (.A(_08244_),
    .ZN(_08245_));
 NOR2_X1 _33778_ (.A1(_08245_),
    .A2(_00040_),
    .ZN(_08246_));
 OR3_X2 _33779_ (.A1(_08089_),
    .A2(\bp_fe_pc_gen_1.btb.r_idx_r [4]),
    .A3(\bp_fe_pc_gen_1.btb.r_idx_r [3]),
    .ZN(_08247_));
 NOR2_X1 _33780_ (.A1(_08247_),
    .A2(_08142_),
    .ZN(_08248_));
 NOR2_X1 _33781_ (.A1(_08246_),
    .A2(_08248_),
    .ZN(_08249_));
 AND2_X1 _33782_ (.A1(_08243_),
    .A2(_08249_),
    .ZN(_08250_));
 AND2_X1 _33783_ (.A1(_08248_),
    .A2(_00039_),
    .ZN(_08251_));
 AND2_X1 _33784_ (.A1(_08054_),
    .A2(_08148_),
    .ZN(_08252_));
 OR2_X1 _33785_ (.A1(_08251_),
    .A2(_08252_),
    .ZN(_08253_));
 OAI21_X2 _33786_ (.A(_08146_),
    .B1(_08250_),
    .B2(_08253_),
    .ZN(_08254_));
 AOI22_X2 _33787_ (.A1(_08145_),
    .A2(_00037_),
    .B1(_00072_),
    .B2(_08133_),
    .ZN(_08255_));
 AOI221_X2 _33788_ (.A(_08136_),
    .B1(_00072_),
    .B2(_08138_),
    .C1(_08254_),
    .C2(_08255_),
    .ZN(_08256_));
 AND4_X1 _33789_ (.A1(_08116_),
    .A2(_08137_),
    .A3(_08055_),
    .A4(_00035_),
    .ZN(_08257_));
 OAI21_X1 _33790_ (.A(_08132_),
    .B1(_08256_),
    .B2(_08257_),
    .ZN(_08258_));
 NOR2_X1 _33791_ (.A1(_08128_),
    .A2(_08083_),
    .ZN(_08259_));
 AOI21_X1 _33792_ (.A(_08259_),
    .B1(_08131_),
    .B2(_00034_),
    .ZN(_08260_));
 AOI21_X1 _33793_ (.A(_08129_),
    .B1(_08258_),
    .B2(_08260_),
    .ZN(_08261_));
 NAND2_X1 _33794_ (.A1(_08191_),
    .A2(_08055_),
    .ZN(_08262_));
 MUX2_X1 _33795_ (.A(_00032_),
    .B(_08261_),
    .S(_08262_),
    .Z(_08263_));
 NAND2_X1 _33796_ (.A1(_08180_),
    .A2(_08055_),
    .ZN(_08264_));
 MUX2_X1 _33797_ (.A(_00031_),
    .B(_08263_),
    .S(_08264_),
    .Z(_08265_));
 NAND3_X1 _33798_ (.A1(_08097_),
    .A2(_08116_),
    .A3(_08055_),
    .ZN(_08266_));
 AOI211_X1 _33799_ (.A(_08124_),
    .B(_08126_),
    .C1(_08265_),
    .C2(_08266_),
    .ZN(_08267_));
 AND2_X1 _33800_ (.A1(_08176_),
    .A2(_08055_),
    .ZN(_08268_));
 INV_X1 _33801_ (.A(_08124_),
    .ZN(_08269_));
 NOR2_X1 _33802_ (.A1(_08269_),
    .A2(_00029_),
    .ZN(_08270_));
 OR3_X1 _33803_ (.A1(_08267_),
    .A2(_08268_),
    .A3(_08270_),
    .ZN(_08271_));
 NAND3_X1 _33804_ (.A1(_08176_),
    .A2(_08055_),
    .A3(_00028_),
    .ZN(_08272_));
 NAND2_X1 _33805_ (.A1(_08271_),
    .A2(_08272_),
    .ZN(_08273_));
 AND2_X1 _33806_ (.A1(_08178_),
    .A2(_08055_),
    .ZN(_08274_));
 MUX2_X1 _33807_ (.A(_08273_),
    .B(_00027_),
    .S(_08274_),
    .Z(_08275_));
 NAND2_X1 _33808_ (.A1(_08174_),
    .A2(_08056_),
    .ZN(_08276_));
 MUX2_X1 _33809_ (.A(_00026_),
    .B(_08275_),
    .S(_08276_),
    .Z(_08277_));
 NAND2_X1 _33810_ (.A1(_08172_),
    .A2(_08056_),
    .ZN(_08278_));
 AOI211_X1 _33811_ (.A(_08118_),
    .B(_08121_),
    .C1(_08277_),
    .C2(_08278_),
    .ZN(_08279_));
 INV_X1 _33812_ (.A(_08118_),
    .ZN(_08280_));
 OAI22_X1 _33813_ (.A1(_08280_),
    .A2(_00024_),
    .B1(_08083_),
    .B2(_08213_),
    .ZN(_08281_));
 OAI21_X1 _33814_ (.A(_08113_),
    .B1(_08279_),
    .B2(_08281_),
    .ZN(_08282_));
 NAND2_X1 _33815_ (.A1(_08169_),
    .A2(_08056_),
    .ZN(_08283_));
 MUX2_X1 _33816_ (.A(_00022_),
    .B(_08282_),
    .S(_08283_),
    .Z(_08284_));
 OR2_X1 _33817_ (.A1(_08165_),
    .A2(_08083_),
    .ZN(_08285_));
 MUX2_X1 _33818_ (.A(_00021_),
    .B(_08284_),
    .S(_08285_),
    .Z(_08286_));
 NAND2_X1 _33819_ (.A1(_08109_),
    .A2(_08057_),
    .ZN(_08287_));
 AOI21_X1 _33820_ (.A(_08111_),
    .B1(_08286_),
    .B2(_08287_),
    .ZN(_08288_));
 NAND3_X1 _33821_ (.A1(_08130_),
    .A2(_08051_),
    .A3(_08056_),
    .ZN(_08289_));
 OAI21_X1 _33822_ (.A(_08289_),
    .B1(_08108_),
    .B2(_00019_),
    .ZN(_08290_));
 OAI21_X1 _33823_ (.A(_08104_),
    .B1(_08288_),
    .B2(_08290_),
    .ZN(_08291_));
 NOR3_X1 _33824_ (.A1(_08119_),
    .A2(\bp_fe_pc_gen_1.btb.r_idx_r [4]),
    .A3(_00070_),
    .ZN(_08292_));
 NAND2_X1 _33825_ (.A1(_08292_),
    .A2(_08057_),
    .ZN(_08293_));
 MUX2_X1 _33826_ (.A(_00017_),
    .B(_08291_),
    .S(_08293_),
    .Z(_08294_));
 NAND2_X1 _33827_ (.A1(_08100_),
    .A2(_08057_),
    .ZN(_08295_));
 AOI21_X1 _33828_ (.A(_08101_),
    .B1(_08294_),
    .B2(_08295_),
    .ZN(_08296_));
 AOI21_X1 _33829_ (.A(_08099_),
    .B1(_08296_),
    .B2(_08092_),
    .ZN(_08297_));
 AND3_X1 _33830_ (.A1(_08122_),
    .A2(_08051_),
    .A3(_08053_),
    .ZN(_08298_));
 AND2_X1 _33831_ (.A1(_08298_),
    .A2(_08057_),
    .ZN(_08299_));
 AND3_X1 _33832_ (.A1(_08157_),
    .A2(_08057_),
    .A3(_00014_),
    .ZN(_08300_));
 OR2_X1 _33833_ (.A1(_08299_),
    .A2(_08300_),
    .ZN(_08301_));
 OAI21_X1 _33834_ (.A(_08087_),
    .B1(_08297_),
    .B2(_08301_),
    .ZN(_08302_));
 NAND3_X1 _33835_ (.A1(_08086_),
    .A2(_08058_),
    .A3(_00012_),
    .ZN(_08303_));
 AOI22_X1 _33836_ (.A1(_08302_),
    .A2(_08303_),
    .B1(_08058_),
    .B2(_08151_),
    .ZN(_08304_));
 AND2_X1 _33837_ (.A1(_08153_),
    .A2(_08058_),
    .ZN(_08305_));
 AND3_X1 _33838_ (.A1(_08151_),
    .A2(_08058_),
    .A3(_00011_),
    .ZN(_08306_));
 OR3_X1 _33839_ (.A1(_08304_),
    .A2(_08305_),
    .A3(_08306_),
    .ZN(_08307_));
 INV_X1 _33840_ (.A(_08305_),
    .ZN(_08308_));
 NOR2_X1 _33841_ (.A1(_08308_),
    .A2(_00010_),
    .ZN(_08309_));
 AND3_X1 _33842_ (.A1(_08120_),
    .A2(_08051_),
    .A3(_08058_),
    .ZN(_08310_));
 NOR2_X1 _33843_ (.A1(_08309_),
    .A2(_08310_),
    .ZN(_08311_));
 AOI22_X1 _33844_ (.A1(_08307_),
    .A2(_08311_),
    .B1(_00009_),
    .B2(_08310_),
    .ZN(_08312_));
 AND2_X1 _33845_ (.A1(_08077_),
    .A2(_08058_),
    .ZN(_08313_));
 OAI21_X1 _33846_ (.A(_08078_),
    .B1(_08312_),
    .B2(_08313_),
    .ZN(_08314_));
 OR2_X2 _33847_ (.A1(_08247_),
    .A2(_08083_),
    .ZN(_08315_));
 MUX2_X2 _33848_ (.A(_00007_),
    .B(_08314_),
    .S(_08315_),
    .Z(_08316_));
 NAND2_X4 _33849_ (.A1(_08054_),
    .A2(_08058_),
    .ZN(_08317_));
 AOI21_X4 _33850_ (.A(_08074_),
    .B1(_08316_),
    .B2(_08317_),
    .ZN(_08318_));
 BUF_X8 _33851_ (.A(_08318_),
    .Z(_08319_));
 BUF_X8 _33852_ (.A(_08319_),
    .Z(_08320_));
 BUF_X8 _33853_ (.A(_08320_),
    .Z(_08321_));
 INV_X2 _33854_ (.A(fe_cmd_v_i),
    .ZN(_08322_));
 NAND2_X1 _33855_ (.A1(_08027_),
    .A2(fe_cmd_i[73]),
    .ZN(_08323_));
 NOR2_X1 _33856_ (.A1(fe_cmd_i[32]),
    .A2(fe_cmd_i[31]),
    .ZN(_08324_));
 NAND2_X1 _33857_ (.A1(_08324_),
    .A2(fe_cmd_i[33]),
    .ZN(_08325_));
 INV_X1 _33858_ (.A(fe_cmd_i[74]),
    .ZN(_08326_));
 AOI211_X2 _33859_ (.A(_08322_),
    .B(_08323_),
    .C1(_08325_),
    .C2(_08326_),
    .ZN(_08327_));
 NOR2_X1 _33860_ (.A1(_08322_),
    .A2(fe_cmd_i[73]),
    .ZN(_08328_));
 AND3_X4 _33861_ (.A1(_08328_),
    .A2(fe_cmd_i[74]),
    .A3(fe_cmd_i[75]),
    .ZN(_08329_));
 NOR2_X2 _33862_ (.A1(_08327_),
    .A2(_08329_),
    .ZN(_08330_));
 INV_X8 _33863_ (.A(_08330_),
    .ZN(_08331_));
 OR3_X2 _33864_ (.A1(fe_cmd_i[73]),
    .A2(fe_cmd_i[74]),
    .A3(fe_cmd_i[75]),
    .ZN(_08332_));
 NOR2_X4 _33865_ (.A1(_08332_),
    .A2(_08322_),
    .ZN(_08333_));
 NOR2_X4 _33866_ (.A1(_08331_),
    .A2(_08333_),
    .ZN(_08334_));
 INV_X1 _33867_ (.A(\bp_fe_pc_gen_1.state_r [1]),
    .ZN(_08335_));
 AND2_X1 _33868_ (.A1(_08335_),
    .A2(\bp_fe_pc_gen_1.state_r [0]),
    .ZN(_08336_));
 BUF_X8 _33869_ (.A(_08336_),
    .Z(_08337_));
 AND2_X4 _33870_ (.A1(_08334_),
    .A2(_08337_),
    .ZN(_08338_));
 BUF_X8 _33871_ (.A(_08338_),
    .Z(_08339_));
 BUF_X8 _33872_ (.A(_08339_),
    .Z(_08340_));
 BUF_X4 _33873_ (.A(_08340_),
    .Z(_08341_));
 NAND3_X2 _33874_ (.A1(_08321_),
    .A2(\bp_fe_pc_gen_1.btb.br_tgt_o [6]),
    .A3(_08341_),
    .ZN(_08342_));
 INV_X1 _33875_ (.A(\bp_fe_pc_gen_1.pc_resume_r [6]),
    .ZN(_08343_));
 INV_X4 _33876_ (.A(_08337_),
    .ZN(_08344_));
 AND2_X4 _33877_ (.A1(_08334_),
    .A2(_08344_),
    .ZN(_08345_));
 INV_X8 _33878_ (.A(_08345_),
    .ZN(_08346_));
 BUF_X8 _33879_ (.A(_08346_),
    .Z(_08347_));
 BUF_X8 _33880_ (.A(_08347_),
    .Z(_08348_));
 INV_X1 _33881_ (.A(fe_cmd_i[40]),
    .ZN(_08349_));
 BUF_X4 _33882_ (.A(_08334_),
    .Z(_08350_));
 OAI221_X2 _33883_ (.A(_08342_),
    .B1(_08343_),
    .B2(_08348_),
    .C1(_08349_),
    .C2(_08350_),
    .ZN(_08351_));
 INV_X8 _33884_ (.A(_08338_),
    .ZN(_08352_));
 BUF_X8 _33885_ (.A(_08352_),
    .Z(_08353_));
 BUF_X8 _33886_ (.A(_08353_),
    .Z(_08354_));
 AND3_X2 _33887_ (.A1(\bp_fe_pc_gen_1.pc_if1_r [4]),
    .A2(\bp_fe_pc_gen_1.pc_if1_r [3]),
    .A3(\bp_fe_pc_gen_1.pc_if1_r [2]),
    .ZN(_08355_));
 AND2_X2 _33888_ (.A1(_08355_),
    .A2(\bp_fe_pc_gen_1.pc_if1_r [5]),
    .ZN(_08356_));
 XOR2_X2 _33889_ (.A(_08356_),
    .B(_00005_),
    .Z(_08357_));
 NOR3_X4 _33890_ (.A1(_08321_),
    .A2(_08354_),
    .A3(_08357_),
    .ZN(_08358_));
 OAI21_X4 _33891_ (.A(_08038_),
    .B1(_08351_),
    .B2(_08358_),
    .ZN(_08359_));
 OR2_X4 _33892_ (.A1(_07984_),
    .A2(_07655_),
    .ZN(_08360_));
 OAI211_X2 _33893_ (.A(_07626_),
    .B(_08360_),
    .C1(_08026_),
    .C2(_08035_),
    .ZN(_08361_));
 NAND2_X4 _33894_ (.A1(_08359_),
    .A2(_08361_),
    .ZN(\icache.tag_mem.addr_i [0]));
 NAND3_X1 _33895_ (.A1(_08321_),
    .A2(\bp_fe_pc_gen_1.btb.br_tgt_o [7]),
    .A3(_08341_),
    .ZN(_08362_));
 INV_X1 _33896_ (.A(\bp_fe_pc_gen_1.pc_resume_r [7]),
    .ZN(_08363_));
 INV_X1 _33897_ (.A(fe_cmd_i[41]),
    .ZN(_08364_));
 OAI221_X2 _33898_ (.A(_08362_),
    .B1(_08363_),
    .B2(_08348_),
    .C1(_08364_),
    .C2(_08350_),
    .ZN(_08365_));
 AND3_X2 _33899_ (.A1(_08355_),
    .A2(\bp_fe_pc_gen_1.pc_if1_r [6]),
    .A3(\bp_fe_pc_gen_1.pc_if1_r [5]),
    .ZN(_08366_));
 XNOR2_X2 _33900_ (.A(_08366_),
    .B(\bp_fe_pc_gen_1.pc_if1_r [7]),
    .ZN(_08367_));
 NOR3_X4 _33901_ (.A1(_08321_),
    .A2(_08354_),
    .A3(_08367_),
    .ZN(_08368_));
 OAI21_X4 _33902_ (.A(_08038_),
    .B1(_08365_),
    .B2(_08368_),
    .ZN(_08369_));
 OAI211_X2 _33903_ (.A(_07632_),
    .B(_08360_),
    .C1(_08026_),
    .C2(_08035_),
    .ZN(_08370_));
 NAND2_X4 _33904_ (.A1(_08369_),
    .A2(_08370_),
    .ZN(\icache.tag_mem.addr_i [1]));
 BUF_X8 _33905_ (.A(_08321_),
    .Z(_08371_));
 NAND3_X1 _33906_ (.A1(_08371_),
    .A2(\bp_fe_pc_gen_1.btb.br_tgt_o [8]),
    .A3(_08341_),
    .ZN(_08372_));
 INV_X1 _33907_ (.A(\bp_fe_pc_gen_1.pc_resume_r [8]),
    .ZN(_08373_));
 INV_X1 _33908_ (.A(fe_cmd_i[42]),
    .ZN(_08374_));
 OAI221_X2 _33909_ (.A(_08372_),
    .B1(_08373_),
    .B2(_08348_),
    .C1(_08374_),
    .C2(_08350_),
    .ZN(_08375_));
 NAND2_X1 _33910_ (.A1(_08366_),
    .A2(\bp_fe_pc_gen_1.pc_if1_r [7]),
    .ZN(_08376_));
 XNOR2_X1 _33911_ (.A(_08376_),
    .B(_00073_),
    .ZN(_08377_));
 NOR3_X2 _33912_ (.A1(_08371_),
    .A2(_08354_),
    .A3(_08377_),
    .ZN(_08378_));
 OAI21_X4 _33913_ (.A(_08038_),
    .B1(_08375_),
    .B2(_08378_),
    .ZN(_08379_));
 OAI211_X2 _33914_ (.A(_07637_),
    .B(_08360_),
    .C1(_08026_),
    .C2(_08035_),
    .ZN(_08380_));
 NAND2_X4 _33915_ (.A1(_08379_),
    .A2(_08380_),
    .ZN(\icache.tag_mem.addr_i [2]));
 NAND3_X1 _33916_ (.A1(_08371_),
    .A2(net1414),
    .A3(_08341_),
    .ZN(_08381_));
 INV_X1 _33917_ (.A(\bp_fe_pc_gen_1.pc_resume_r [9]),
    .ZN(_08382_));
 INV_X1 _33918_ (.A(fe_cmd_i[43]),
    .ZN(_08383_));
 OAI221_X2 _33919_ (.A(_08381_),
    .B1(_08382_),
    .B2(_08348_),
    .C1(_08383_),
    .C2(_08350_),
    .ZN(_08384_));
 NAND3_X2 _33920_ (.A1(_08366_),
    .A2(\bp_fe_pc_gen_1.pc_if1_r [7]),
    .A3(\bp_fe_pc_gen_1.pc_if1_r [8]),
    .ZN(_08385_));
 INV_X2 _33921_ (.A(\bp_fe_pc_gen_1.pc_if1_r [9]),
    .ZN(_08386_));
 XNOR2_X2 _33922_ (.A(_08385_),
    .B(_08386_),
    .ZN(_08387_));
 NOR3_X4 _33923_ (.A1(_08371_),
    .A2(_08354_),
    .A3(_08387_),
    .ZN(_08388_));
 OAI21_X4 _33924_ (.A(_08038_),
    .B1(_08384_),
    .B2(_08388_),
    .ZN(_08389_));
 OAI211_X2 _33925_ (.A(_07642_),
    .B(_08360_),
    .C1(_08026_),
    .C2(_08035_),
    .ZN(_08390_));
 NAND2_X4 _33926_ (.A1(_08389_),
    .A2(_08390_),
    .ZN(\icache.tag_mem.addr_i [3]));
 NAND3_X1 _33927_ (.A1(_08371_),
    .A2(net1413),
    .A3(_08341_),
    .ZN(_08391_));
 INV_X1 _33928_ (.A(\bp_fe_pc_gen_1.pc_resume_r [10]),
    .ZN(_08392_));
 INV_X2 _33929_ (.A(fe_cmd_i[44]),
    .ZN(_08393_));
 OAI221_X2 _33930_ (.A(_08391_),
    .B1(_08392_),
    .B2(_08348_),
    .C1(_08393_),
    .C2(_08350_),
    .ZN(_08394_));
 NOR2_X1 _33931_ (.A1(_08385_),
    .A2(_08386_),
    .ZN(_08395_));
 XOR2_X2 _33932_ (.A(_08395_),
    .B(_00074_),
    .Z(_08396_));
 NOR3_X4 _33933_ (.A1(_08371_),
    .A2(_08354_),
    .A3(_08396_),
    .ZN(_08397_));
 OAI21_X4 _33934_ (.A(_08038_),
    .B1(_08394_),
    .B2(_08397_),
    .ZN(_08398_));
 OAI211_X2 _33935_ (.A(_07647_),
    .B(_08360_),
    .C1(_08026_),
    .C2(_08035_),
    .ZN(_08399_));
 NAND2_X4 _33936_ (.A1(_08398_),
    .A2(_08399_),
    .ZN(\icache.tag_mem.addr_i [4]));
 NAND3_X1 _33937_ (.A1(_08371_),
    .A2(\bp_fe_pc_gen_1.btb.br_tgt_o [11]),
    .A3(_08341_),
    .ZN(_08400_));
 INV_X1 _33938_ (.A(\bp_fe_pc_gen_1.pc_resume_r [11]),
    .ZN(_08401_));
 INV_X2 _33939_ (.A(fe_cmd_i[45]),
    .ZN(_08402_));
 OAI221_X2 _33940_ (.A(_08400_),
    .B1(_08401_),
    .B2(_08348_),
    .C1(_08402_),
    .C2(_08350_),
    .ZN(_08403_));
 AND2_X1 _33941_ (.A1(_08395_),
    .A2(\bp_fe_pc_gen_1.pc_if1_r [10]),
    .ZN(_08404_));
 XNOR2_X2 _33942_ (.A(_08404_),
    .B(\bp_fe_pc_gen_1.pc_if1_r [11]),
    .ZN(_08405_));
 NOR3_X4 _33943_ (.A1(_08371_),
    .A2(_08354_),
    .A3(_08405_),
    .ZN(_08406_));
 OAI21_X4 _33944_ (.A(_08038_),
    .B1(_08403_),
    .B2(_08406_),
    .ZN(_08407_));
 OAI211_X2 _33945_ (.A(_07652_),
    .B(_08360_),
    .C1(_08026_),
    .C2(_08035_),
    .ZN(_08408_));
 NAND2_X4 _33946_ (.A1(_08407_),
    .A2(_08408_),
    .ZN(\icache.tag_mem.addr_i [5]));
 NOR2_X2 _33947_ (.A1(_08321_),
    .A2(_08354_),
    .ZN(_08409_));
 INV_X2 _33948_ (.A(_08409_),
    .ZN(_08410_));
 AND2_X1 _33949_ (.A1(\bp_fe_pc_gen_1.pc_if1_r [3]),
    .A2(\bp_fe_pc_gen_1.pc_if1_r [2]),
    .ZN(_08411_));
 AOI21_X2 _33950_ (.A(\bp_fe_pc_gen_1.pc_if1_r [5]),
    .B1(_08411_),
    .B2(\bp_fe_pc_gen_1.pc_if1_r [4]),
    .ZN(_08412_));
 NOR3_X4 _33951_ (.A1(_08410_),
    .A2(_08356_),
    .A3(_08412_),
    .ZN(_08413_));
 NAND3_X2 _33952_ (.A1(_08321_),
    .A2(net1415),
    .A3(_08341_),
    .ZN(_08414_));
 INV_X1 _33953_ (.A(\bp_fe_pc_gen_1.pc_resume_r [5]),
    .ZN(_08415_));
 INV_X1 _33954_ (.A(fe_cmd_i[39]),
    .ZN(_08416_));
 OAI221_X2 _33955_ (.A(_08414_),
    .B1(_08415_),
    .B2(_08348_),
    .C1(_08416_),
    .C2(_08350_),
    .ZN(_08417_));
 OAI21_X4 _33956_ (.A(_08038_),
    .B1(_08413_),
    .B2(_08417_),
    .ZN(_08418_));
 BUF_X8 _33957_ (.A(_08037_),
    .Z(_08419_));
 AOI21_X4 _33958_ (.A(_07612_),
    .B1(_07614_),
    .B2(_07615_),
    .ZN(_08420_));
 BUF_X8 _33959_ (.A(_08420_),
    .Z(_08421_));
 AND3_X4 _33960_ (.A1(_07604_),
    .A2(_07605_),
    .A3(\icache.lce.N14 ),
    .ZN(_08422_));
 NAND4_X4 _33961_ (.A1(_08421_),
    .A2(_07978_),
    .A3(_07987_),
    .A4(_08422_),
    .ZN(_08423_));
 INV_X16 _33962_ (.A(net1394),
    .ZN(_08424_));
 OR2_X1 _33963_ (.A1(_08424_),
    .A2(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [520]),
    .ZN(_08425_));
 INV_X16 _33964_ (.A(net1397),
    .ZN(_08426_));
 BUF_X32 _33965_ (.A(net1396),
    .Z(_08427_));
 BUF_X16 _33966_ (.A(_08427_),
    .Z(_08428_));
 OAI211_X1 _33967_ (.A(_08425_),
    .B(_08426_),
    .C1(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [2]),
    .C2(_08428_),
    .ZN(_08429_));
 AND2_X2 _33968_ (.A1(_08423_),
    .A2(_08429_),
    .ZN(_08430_));
 BUF_X16 _33969_ (.A(_08430_),
    .Z(_08431_));
 INV_X8 _33970_ (.A(_08431_),
    .ZN(_08432_));
 BUF_X8 _33971_ (.A(_08432_),
    .Z(_08433_));
 BUF_X32 _33972_ (.A(_08433_),
    .Z(_08434_));
 OAI21_X4 _33973_ (.A(_08418_),
    .B1(_08419_),
    .B2(_08434_),
    .ZN(\icache.data_mem_addr_li [38]));
 AOI21_X2 _33974_ (.A(\bp_fe_pc_gen_1.pc_if1_r [4]),
    .B1(\bp_fe_pc_gen_1.pc_if1_r [3]),
    .B2(\bp_fe_pc_gen_1.pc_if1_r [2]),
    .ZN(_08435_));
 NOR3_X4 _33975_ (.A1(_08410_),
    .A2(_08355_),
    .A3(_08435_),
    .ZN(_08436_));
 NAND3_X1 _33976_ (.A1(_08321_),
    .A2(\bp_fe_pc_gen_1.btb.br_tgt_o [4]),
    .A3(_08341_),
    .ZN(_08437_));
 INV_X1 _33977_ (.A(\bp_fe_pc_gen_1.pc_resume_r [4]),
    .ZN(_08438_));
 INV_X1 _33978_ (.A(fe_cmd_i[38]),
    .ZN(_08439_));
 OAI221_X2 _33979_ (.A(_08437_),
    .B1(_08438_),
    .B2(_08348_),
    .C1(_08439_),
    .C2(_08350_),
    .ZN(_08440_));
 OAI21_X4 _33980_ (.A(_08038_),
    .B1(_08436_),
    .B2(_08440_),
    .ZN(_08441_));
 NAND4_X4 _33981_ (.A1(_08421_),
    .A2(_07978_),
    .A3(_07991_),
    .A4(_08422_),
    .ZN(_08442_));
 OR2_X1 _33982_ (.A1(net1395),
    .A2(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1]),
    .ZN(_08443_));
 OAI211_X1 _33983_ (.A(_08443_),
    .B(_08426_),
    .C1(_08424_),
    .C2(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [519]),
    .ZN(_08444_));
 AND2_X4 _33984_ (.A1(_08442_),
    .A2(_08444_),
    .ZN(_08445_));
 BUF_X16 _33985_ (.A(_08445_),
    .Z(_08446_));
 INV_X16 _33986_ (.A(_08446_),
    .ZN(_08447_));
 BUF_X32 _33987_ (.A(_08447_),
    .Z(_08448_));
 OAI21_X4 _33988_ (.A(_08441_),
    .B1(_08419_),
    .B2(_08448_),
    .ZN(\icache.data_mem_addr_li [19]));
 NOR2_X1 _33989_ (.A1(\bp_fe_pc_gen_1.pc_if1_r [3]),
    .A2(\bp_fe_pc_gen_1.pc_if1_r [2]),
    .ZN(_08449_));
 OR3_X1 _33990_ (.A1(_08410_),
    .A2(_08411_),
    .A3(_08449_),
    .ZN(_08450_));
 NAND2_X2 _33991_ (.A1(_08316_),
    .A2(_08317_),
    .ZN(_08451_));
 NOR2_X1 _33992_ (.A1(_08061_),
    .A2(\bp_fe_pc_gen_1.btb.r_tag_r [1]),
    .ZN(_08452_));
 NOR3_X1 _33993_ (.A1(_08039_),
    .A2(_08452_),
    .A3(_08060_),
    .ZN(_08453_));
 INV_X1 _33994_ (.A(\bp_fe_pc_gen_1.btb.r_tag_r [4]),
    .ZN(_08454_));
 AOI22_X1 _33995_ (.A1(_08454_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.data_o [43]),
    .B1(_08040_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.data_o [44]),
    .ZN(_08455_));
 NAND2_X1 _33996_ (.A1(_08061_),
    .A2(\bp_fe_pc_gen_1.btb.r_tag_r [1]),
    .ZN(_08456_));
 AND4_X1 _33997_ (.A1(_08453_),
    .A2(_08455_),
    .A3(_08044_),
    .A4(_08456_),
    .ZN(_08457_));
 INV_X1 _33998_ (.A(net1399),
    .ZN(_08458_));
 NAND2_X1 _33999_ (.A1(_08458_),
    .A2(\bp_fe_pc_gen_1.btb.r_tag_r [6]),
    .ZN(_08459_));
 INV_X1 _34000_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.data_o [47]),
    .ZN(_08460_));
 OAI21_X1 _34001_ (.A(_08459_),
    .B1(\bp_fe_pc_gen_1.btb.r_tag_r [8]),
    .B2(_08460_),
    .ZN(_08461_));
 OAI22_X1 _34002_ (.A1(_08454_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.data_o [43]),
    .B1(_08458_),
    .B2(\bp_fe_pc_gen_1.btb.r_tag_r [6]),
    .ZN(_08462_));
 AND2_X1 _34003_ (.A1(_08460_),
    .A2(\bp_fe_pc_gen_1.btb.r_tag_r [8]),
    .ZN(_08463_));
 NOR4_X1 _34004_ (.A1(_08461_),
    .A2(_08462_),
    .A3(_08463_),
    .A4(_08072_),
    .ZN(_08464_));
 AOI22_X1 _34005_ (.A1(_08046_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.data_o [39]),
    .B1(_08041_),
    .B2(\bp_fe_pc_gen_1.btb.r_tag_r [7]),
    .ZN(_08465_));
 OAI211_X1 _34006_ (.A(_08465_),
    .B(_08063_),
    .C1(\bp_fe_pc_gen_1.btb.r_tag_r [7]),
    .C2(_08041_),
    .ZN(_08466_));
 OAI22_X1 _34007_ (.A1(_08040_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.data_o [44]),
    .B1(_08069_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.data_o [48]),
    .ZN(_08467_));
 NOR3_X1 _34008_ (.A1(_08466_),
    .A2(_08071_),
    .A3(_08467_),
    .ZN(_08468_));
 AND4_X1 _34009_ (.A1(_08059_),
    .A2(_08457_),
    .A3(_08464_),
    .A4(_08468_),
    .ZN(_08469_));
 AND2_X1 _34010_ (.A1(_08451_),
    .A2(_08469_),
    .ZN(_08470_));
 NAND2_X1 _34011_ (.A1(_08470_),
    .A2(_08340_),
    .ZN(_08471_));
 OR2_X1 _34012_ (.A1(_08471_),
    .A2(_00077_),
    .ZN(_08472_));
 NAND3_X1 _34013_ (.A1(_08450_),
    .A2(_08348_),
    .A3(_08472_),
    .ZN(_08473_));
 NAND3_X2 _34014_ (.A1(_08350_),
    .A2(_00076_),
    .A3(_08344_),
    .ZN(_08474_));
 NAND2_X4 _34015_ (.A1(_08473_),
    .A2(_08474_),
    .ZN(_08475_));
 BUF_X8 _34016_ (.A(_08331_),
    .Z(_08476_));
 BUF_X8 _34017_ (.A(_08333_),
    .Z(_08477_));
 OAI21_X4 _34018_ (.A(fe_cmd_i[37]),
    .B1(_08476_),
    .B2(_08477_),
    .ZN(_08478_));
 AND3_X4 _34019_ (.A1(_08475_),
    .A2(_08037_),
    .A3(_08478_),
    .ZN(_08479_));
 INV_X8 _34020_ (.A(_08036_),
    .ZN(_08480_));
 BUF_X8 _34021_ (.A(_08480_),
    .Z(_08481_));
 AND4_X4 _34022_ (.A1(_07978_),
    .A2(_08420_),
    .A3(_07995_),
    .A4(_08422_),
    .ZN(_08482_));
 BUF_X16 _34023_ (.A(_08482_),
    .Z(_08483_));
 NAND2_X1 _34024_ (.A1(_08424_),
    .A2(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [0]),
    .ZN(_08484_));
 NAND2_X1 _34025_ (.A1(net1395),
    .A2(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [518]),
    .ZN(_08485_));
 AOI21_X4 _34026_ (.A(net1397),
    .B1(_08484_),
    .B2(_08485_),
    .ZN(_08486_));
 BUF_X16 _34027_ (.A(_08486_),
    .Z(_08487_));
 NOR2_X2 _34028_ (.A1(_08483_),
    .A2(_08487_),
    .ZN(_08488_));
 BUF_X16 _34029_ (.A(_08488_),
    .Z(_08489_));
 BUF_X16 _34030_ (.A(_08489_),
    .Z(_08490_));
 BUF_X16 _34031_ (.A(_08490_),
    .Z(_08491_));
 INV_X4 _34032_ (.A(_08491_),
    .ZN(_08492_));
 AOI21_X4 _34033_ (.A(_08479_),
    .B1(_08481_),
    .B2(_08492_),
    .ZN(\icache.data_mem_addr_li [27]));
 AOI21_X4 _34034_ (.A(_08479_),
    .B1(_08481_),
    .B2(_08491_),
    .ZN(\icache.data_mem_addr_li [0]));
 BUF_X16 _34035_ (.A(_08446_),
    .Z(_08493_));
 BUF_X16 _34036_ (.A(_08493_),
    .Z(_08494_));
 OAI21_X4 _34037_ (.A(_08441_),
    .B1(_08419_),
    .B2(_08494_),
    .ZN(\icache.data_mem_addr_li [10]));
 BUF_X16 _34038_ (.A(_08431_),
    .Z(_08495_));
 BUF_X16 _34039_ (.A(_08495_),
    .Z(_08496_));
 OAI21_X4 _34040_ (.A(_08418_),
    .B1(_08419_),
    .B2(_08496_),
    .ZN(\icache.data_mem_addr_li [11]));
 AND2_X1 _34041_ (.A1(_08420_),
    .A2(_07978_),
    .ZN(_08497_));
 AND2_X1 _34042_ (.A1(_08497_),
    .A2(_08422_),
    .ZN(_08498_));
 BUF_X8 _34043_ (.A(_08498_),
    .Z(_08499_));
 BUF_X16 _34044_ (.A(_08426_),
    .Z(_08500_));
 BUF_X16 _34045_ (.A(_08500_),
    .Z(_08501_));
 AOI22_X2 _34046_ (.A1(_08499_),
    .A2(_07626_),
    .B1(_08501_),
    .B2(lce_req_o[13]),
    .ZN(_08502_));
 OAI21_X4 _34047_ (.A(_08359_),
    .B1(_08419_),
    .B2(_08502_),
    .ZN(\icache.data_mem_addr_li [12]));
 AOI22_X2 _34048_ (.A1(_08499_),
    .A2(_07632_),
    .B1(_08501_),
    .B2(lce_req_o[14]),
    .ZN(_08503_));
 OAI21_X4 _34049_ (.A(_08369_),
    .B1(_08419_),
    .B2(_08503_),
    .ZN(\icache.data_mem_addr_li [13]));
 AOI22_X2 _34050_ (.A1(_08499_),
    .A2(_07637_),
    .B1(_08501_),
    .B2(lce_req_o[15]),
    .ZN(_08504_));
 OAI21_X4 _34051_ (.A(_08379_),
    .B1(_08419_),
    .B2(_08504_),
    .ZN(\icache.data_mem_addr_li [14]));
 AOI22_X2 _34052_ (.A1(_08499_),
    .A2(_07642_),
    .B1(_08501_),
    .B2(lce_req_o[16]),
    .ZN(_08505_));
 OAI21_X4 _34053_ (.A(_08389_),
    .B1(_08419_),
    .B2(_08505_),
    .ZN(\icache.data_mem_addr_li [15]));
 AOI22_X2 _34054_ (.A1(_08499_),
    .A2(_07647_),
    .B1(_08501_),
    .B2(lce_req_o[17]),
    .ZN(_08506_));
 OAI21_X4 _34055_ (.A(_08398_),
    .B1(_08419_),
    .B2(_08506_),
    .ZN(\icache.data_mem_addr_li [16]));
 AOI22_X2 _34056_ (.A1(_08499_),
    .A2(_07652_),
    .B1(_08501_),
    .B2(lce_req_o[18]),
    .ZN(_08507_));
 OAI21_X4 _34057_ (.A(_08407_),
    .B1(_08419_),
    .B2(_08507_),
    .ZN(\icache.data_mem_addr_li [17]));
 OR2_X2 _34058_ (.A1(_08017_),
    .A2(_08024_),
    .ZN(_08508_));
 INV_X1 _34059_ (.A(_08028_),
    .ZN(_08509_));
 NOR2_X4 _34060_ (.A1(_08509_),
    .A2(fe_cmd_i[73]),
    .ZN(_08510_));
 NOR2_X4 _34061_ (.A1(_08510_),
    .A2(_08322_),
    .ZN(_08511_));
 INV_X4 _34062_ (.A(_08511_),
    .ZN(_08512_));
 AND2_X4 _34063_ (.A1(_08508_),
    .A2(_08512_),
    .ZN(_08513_));
 INV_X1 _34064_ (.A(\bp_fe_pc_gen_1.itlb_miss_i ),
    .ZN(_08514_));
 NAND4_X4 _34065_ (.A1(_08513_),
    .A2(\icache.itlb_icache_data_resp_ready_o ),
    .A3(\icache.itlb_icache_data_resp_v_i ),
    .A4(_08514_),
    .ZN(_08515_));
 BUF_X32 _34066_ (.A(reset_i),
    .Z(_08516_));
 NOR2_X4 _34067_ (.A1(_08515_),
    .A2(_08516_),
    .ZN(_08517_));
 BUF_X16 _34068_ (.A(_08517_),
    .Z(_08518_));
 BUF_X8 _34069_ (.A(_08518_),
    .Z(\icache.N29 ));
 INV_X8 _34070_ (.A(_08516_),
    .ZN(_08519_));
 AND2_X1 _34071_ (.A1(_08037_),
    .A2(_08519_),
    .ZN(_08520_));
 BUF_X8 _34072_ (.A(_08520_),
    .Z(_08521_));
 BUF_X16 _34073_ (.A(_08521_),
    .Z(\icache.N25 ));
 NOR2_X4 _34074_ (.A1(_08511_),
    .A2(_08344_),
    .ZN(_08522_));
 BUF_X4 _34075_ (.A(_08522_),
    .Z(_08523_));
 BUF_X8 _34076_ (.A(fe_cmd_i[34]),
    .Z(_08524_));
 BUF_X4 _34077_ (.A(_08511_),
    .Z(_08525_));
 AOI22_X1 _34078_ (.A1(_08523_),
    .A2(\bp_fe_pc_gen_1.pc_if2_r [0]),
    .B1(_08524_),
    .B2(_08525_),
    .ZN(_08526_));
 BUF_X4 _34079_ (.A(_08512_),
    .Z(_08527_));
 NAND3_X1 _34080_ (.A1(_08527_),
    .A2(\bp_fe_pc_gen_1.pc_resume_r [0]),
    .A3(_08344_),
    .ZN(_08528_));
 NAND2_X1 _34081_ (.A1(_08526_),
    .A2(_08528_),
    .ZN(_00688_));
 BUF_X8 _34082_ (.A(fe_cmd_i[35]),
    .Z(_08529_));
 AOI22_X1 _34083_ (.A1(_08523_),
    .A2(\bp_fe_pc_gen_1.pc_if2_r [1]),
    .B1(_08529_),
    .B2(_08525_),
    .ZN(_08530_));
 NAND3_X1 _34084_ (.A1(_08527_),
    .A2(\bp_fe_pc_gen_1.pc_resume_r [1]),
    .A3(_08344_),
    .ZN(_08531_));
 NAND2_X1 _34085_ (.A1(_08530_),
    .A2(_08531_),
    .ZN(_00699_));
 BUF_X4 _34086_ (.A(_08512_),
    .Z(_08532_));
 BUF_X4 _34087_ (.A(_08337_),
    .Z(_08533_));
 NAND3_X1 _34088_ (.A1(_08532_),
    .A2(\bp_fe_pc_gen_1.pc_if2_r [2]),
    .A3(_08533_),
    .ZN(_08534_));
 NAND3_X1 _34089_ (.A1(_08532_),
    .A2(\bp_fe_pc_gen_1.pc_resume_r [2]),
    .A3(_08344_),
    .ZN(_08535_));
 INV_X1 _34090_ (.A(fe_cmd_i[36]),
    .ZN(_08536_));
 OAI211_X1 _34091_ (.A(_08534_),
    .B(_08535_),
    .C1(_08536_),
    .C2(_08527_),
    .ZN(_00710_));
 BUF_X8 _34092_ (.A(fe_cmd_i[37]),
    .Z(_08537_));
 AOI22_X1 _34093_ (.A1(_08523_),
    .A2(\bp_fe_pc_gen_1.pc_if2_r [3]),
    .B1(_08537_),
    .B2(_08525_),
    .ZN(_08538_));
 NAND3_X1 _34094_ (.A1(_08527_),
    .A2(\bp_fe_pc_gen_1.pc_resume_r [3]),
    .A3(_08344_),
    .ZN(_08539_));
 NAND2_X1 _34095_ (.A1(_08538_),
    .A2(_08539_),
    .ZN(_00720_));
 NAND3_X1 _34096_ (.A1(_08532_),
    .A2(\bp_fe_pc_gen_1.pc_if2_r [4]),
    .A3(_08533_),
    .ZN(_08540_));
 OR2_X1 _34097_ (.A1(_08511_),
    .A2(_08337_),
    .ZN(_08541_));
 BUF_X8 _34098_ (.A(_08541_),
    .Z(_08542_));
 BUF_X8 _34099_ (.A(_08542_),
    .Z(_08543_));
 OAI221_X1 _34100_ (.A(_08540_),
    .B1(_08439_),
    .B2(_08527_),
    .C1(_08543_),
    .C2(_08438_),
    .ZN(_00721_));
 NAND3_X1 _34101_ (.A1(_08532_),
    .A2(\bp_fe_pc_gen_1.pc_if2_r [5]),
    .A3(_08533_),
    .ZN(_08544_));
 OAI221_X1 _34102_ (.A(_08544_),
    .B1(_08416_),
    .B2(_08527_),
    .C1(_08543_),
    .C2(_08415_),
    .ZN(_00722_));
 NAND3_X1 _34103_ (.A1(_08532_),
    .A2(\bp_fe_pc_gen_1.pc_if2_r [6]),
    .A3(_08533_),
    .ZN(_08545_));
 OAI221_X1 _34104_ (.A(_08545_),
    .B1(_08349_),
    .B2(_08527_),
    .C1(_08543_),
    .C2(_08343_),
    .ZN(_00723_));
 NAND3_X1 _34105_ (.A1(_08532_),
    .A2(\bp_fe_pc_gen_1.pc_if2_r [7]),
    .A3(_08533_),
    .ZN(_08546_));
 OAI221_X1 _34106_ (.A(_08546_),
    .B1(_08364_),
    .B2(_08527_),
    .C1(_08542_),
    .C2(_08363_),
    .ZN(_00724_));
 NAND3_X1 _34107_ (.A1(_08532_),
    .A2(\bp_fe_pc_gen_1.pc_if2_r [8]),
    .A3(_08533_),
    .ZN(_08547_));
 OAI221_X1 _34108_ (.A(_08547_),
    .B1(_08374_),
    .B2(_08527_),
    .C1(_08542_),
    .C2(_08373_),
    .ZN(_00725_));
 NAND3_X1 _34109_ (.A1(_08532_),
    .A2(\bp_fe_pc_gen_1.pc_if2_r [9]),
    .A3(_08533_),
    .ZN(_08548_));
 OAI221_X1 _34110_ (.A(_08548_),
    .B1(_08383_),
    .B2(_08527_),
    .C1(_08542_),
    .C2(_08382_),
    .ZN(_00726_));
 NAND3_X1 _34111_ (.A1(_08512_),
    .A2(\bp_fe_pc_gen_1.pc_if2_r [10]),
    .A3(_08533_),
    .ZN(_08549_));
 OAI221_X1 _34112_ (.A(_08549_),
    .B1(_08393_),
    .B2(_08532_),
    .C1(_08542_),
    .C2(_08392_),
    .ZN(_00689_));
 NAND3_X1 _34113_ (.A1(_08512_),
    .A2(\bp_fe_pc_gen_1.pc_if2_r [11]),
    .A3(_08533_),
    .ZN(_08550_));
 OAI221_X1 _34114_ (.A(_08550_),
    .B1(_08402_),
    .B2(_08532_),
    .C1(_08542_),
    .C2(_08401_),
    .ZN(_00690_));
 BUF_X32 _34115_ (.A(fe_cmd_i[46]),
    .Z(_08551_));
 AOI22_X1 _34116_ (.A1(_08523_),
    .A2(\bp_fe_pc_gen_1.pc_if2_r [12]),
    .B1(_08551_),
    .B2(_08525_),
    .ZN(_08552_));
 INV_X2 _34117_ (.A(\bp_fe_pc_gen_1.pc_resume_r [12]),
    .ZN(_08553_));
 BUF_X8 _34118_ (.A(_08542_),
    .Z(_08554_));
 OAI21_X1 _34119_ (.A(_08552_),
    .B1(_08553_),
    .B2(_08554_),
    .ZN(_00691_));
 BUF_X32 _34120_ (.A(fe_cmd_i[47]),
    .Z(_08555_));
 AOI22_X1 _34121_ (.A1(_08523_),
    .A2(\bp_fe_pc_gen_1.pc_if2_r [13]),
    .B1(_08555_),
    .B2(_08525_),
    .ZN(_08556_));
 INV_X1 _34122_ (.A(\bp_fe_pc_gen_1.pc_resume_r [13]),
    .ZN(_08557_));
 OAI21_X1 _34123_ (.A(_08556_),
    .B1(_08557_),
    .B2(_08554_),
    .ZN(_00692_));
 BUF_X32 _34124_ (.A(fe_cmd_i[48]),
    .Z(_08558_));
 AOI22_X1 _34125_ (.A1(_08523_),
    .A2(\bp_fe_pc_gen_1.pc_if2_r [14]),
    .B1(_08558_),
    .B2(_08525_),
    .ZN(_08559_));
 INV_X1 _34126_ (.A(\bp_fe_pc_gen_1.pc_resume_r [14]),
    .ZN(_08560_));
 OAI21_X1 _34127_ (.A(_08559_),
    .B1(_08560_),
    .B2(_08554_),
    .ZN(_00693_));
 BUF_X32 _34128_ (.A(fe_cmd_i[49]),
    .Z(_08561_));
 AOI22_X2 _34129_ (.A1(_08523_),
    .A2(\bp_fe_pc_gen_1.pc_if2_r [15]),
    .B1(_08561_),
    .B2(_08525_),
    .ZN(_08562_));
 INV_X1 _34130_ (.A(\bp_fe_pc_gen_1.pc_resume_r [15]),
    .ZN(_08563_));
 OAI21_X1 _34131_ (.A(_08562_),
    .B1(_08563_),
    .B2(_08554_),
    .ZN(_00694_));
 BUF_X32 _34132_ (.A(fe_cmd_i[50]),
    .Z(_08564_));
 AOI22_X1 _34133_ (.A1(_08523_),
    .A2(\bp_fe_pc_gen_1.pc_if2_r [16]),
    .B1(_08564_),
    .B2(_08525_),
    .ZN(_08565_));
 INV_X2 _34134_ (.A(\bp_fe_pc_gen_1.pc_resume_r [16]),
    .ZN(_08566_));
 OAI21_X1 _34135_ (.A(_08565_),
    .B1(_08566_),
    .B2(_08554_),
    .ZN(_00695_));
 BUF_X32 _34136_ (.A(fe_cmd_i[51]),
    .Z(_08567_));
 AOI22_X1 _34137_ (.A1(_08523_),
    .A2(\bp_fe_pc_gen_1.pc_if2_r [17]),
    .B1(_08567_),
    .B2(_08525_),
    .ZN(_08568_));
 INV_X1 _34138_ (.A(\bp_fe_pc_gen_1.pc_resume_r [17]),
    .ZN(_08569_));
 OAI21_X1 _34139_ (.A(_08568_),
    .B1(_08569_),
    .B2(_08554_),
    .ZN(_00696_));
 BUF_X4 _34140_ (.A(_08522_),
    .Z(_08570_));
 BUF_X32 _34141_ (.A(fe_cmd_i[52]),
    .Z(_08571_));
 BUF_X4 _34142_ (.A(_08511_),
    .Z(_08572_));
 AOI22_X1 _34143_ (.A1(_08570_),
    .A2(\bp_fe_pc_gen_1.pc_if2_r [18]),
    .B1(_08571_),
    .B2(_08572_),
    .ZN(_08573_));
 INV_X1 _34144_ (.A(\bp_fe_pc_gen_1.pc_resume_r [18]),
    .ZN(_08574_));
 OAI21_X1 _34145_ (.A(_08573_),
    .B1(_08574_),
    .B2(_08554_),
    .ZN(_00697_));
 BUF_X16 _34146_ (.A(fe_cmd_i[53]),
    .Z(_08575_));
 AOI22_X1 _34147_ (.A1(_08570_),
    .A2(\bp_fe_pc_gen_1.pc_if2_r [19]),
    .B1(_08575_),
    .B2(_08572_),
    .ZN(_08576_));
 INV_X1 _34148_ (.A(\bp_fe_pc_gen_1.pc_resume_r [19]),
    .ZN(_08577_));
 OAI21_X1 _34149_ (.A(_08576_),
    .B1(_08577_),
    .B2(_08554_),
    .ZN(_00698_));
 BUF_X32 _34150_ (.A(fe_cmd_i[54]),
    .Z(_08578_));
 AOI22_X1 _34151_ (.A1(_08570_),
    .A2(\bp_fe_pc_gen_1.pc_if2_r [20]),
    .B1(_08578_),
    .B2(_08572_),
    .ZN(_08579_));
 INV_X1 _34152_ (.A(\bp_fe_pc_gen_1.pc_resume_r [20]),
    .ZN(_08580_));
 OAI21_X1 _34153_ (.A(_08579_),
    .B1(_08580_),
    .B2(_08554_),
    .ZN(_00700_));
 BUF_X32 _34154_ (.A(fe_cmd_i[55]),
    .Z(_08581_));
 AOI22_X1 _34155_ (.A1(_08570_),
    .A2(\bp_fe_pc_gen_1.pc_if2_r [21]),
    .B1(_08581_),
    .B2(_08572_),
    .ZN(_08582_));
 INV_X1 _34156_ (.A(\bp_fe_pc_gen_1.pc_resume_r [21]),
    .ZN(_08583_));
 OAI21_X1 _34157_ (.A(_08582_),
    .B1(_08583_),
    .B2(_08554_),
    .ZN(_00701_));
 BUF_X32 _34158_ (.A(fe_cmd_i[56]),
    .Z(_08584_));
 AOI22_X1 _34159_ (.A1(_08570_),
    .A2(\bp_fe_pc_gen_1.pc_if2_r [22]),
    .B1(_08584_),
    .B2(_08572_),
    .ZN(_08585_));
 INV_X1 _34160_ (.A(\bp_fe_pc_gen_1.pc_resume_r [22]),
    .ZN(_08586_));
 BUF_X4 _34161_ (.A(_08542_),
    .Z(_08587_));
 OAI21_X1 _34162_ (.A(_08585_),
    .B1(_08586_),
    .B2(_08587_),
    .ZN(_00702_));
 BUF_X32 _34163_ (.A(fe_cmd_i[57]),
    .Z(_08588_));
 AOI22_X1 _34164_ (.A1(_08570_),
    .A2(\bp_fe_pc_gen_1.pc_if2_r [23]),
    .B1(_08588_),
    .B2(_08572_),
    .ZN(_08589_));
 INV_X1 _34165_ (.A(\bp_fe_pc_gen_1.pc_resume_r [23]),
    .ZN(_08590_));
 OAI21_X1 _34166_ (.A(_08589_),
    .B1(_08590_),
    .B2(_08587_),
    .ZN(_00703_));
 BUF_X32 _34167_ (.A(fe_cmd_i[58]),
    .Z(_08591_));
 AOI22_X1 _34168_ (.A1(_08570_),
    .A2(\bp_fe_pc_gen_1.pc_if2_r [24]),
    .B1(_08591_),
    .B2(_08572_),
    .ZN(_08592_));
 INV_X1 _34169_ (.A(\bp_fe_pc_gen_1.pc_resume_r [24]),
    .ZN(_08593_));
 OAI21_X1 _34170_ (.A(_08592_),
    .B1(_08593_),
    .B2(_08587_),
    .ZN(_00704_));
 BUF_X32 _34171_ (.A(fe_cmd_i[59]),
    .Z(_08594_));
 AOI22_X1 _34172_ (.A1(_08570_),
    .A2(\bp_fe_pc_gen_1.pc_if2_r [25]),
    .B1(_08594_),
    .B2(_08572_),
    .ZN(_08595_));
 INV_X1 _34173_ (.A(\bp_fe_pc_gen_1.pc_resume_r [25]),
    .ZN(_08596_));
 OAI21_X1 _34174_ (.A(_08595_),
    .B1(_08596_),
    .B2(_08587_),
    .ZN(_00705_));
 BUF_X32 _34175_ (.A(fe_cmd_i[60]),
    .Z(_08597_));
 AOI22_X1 _34176_ (.A1(_08570_),
    .A2(\bp_fe_pc_gen_1.pc_if2_r [26]),
    .B1(_08597_),
    .B2(_08572_),
    .ZN(_08598_));
 INV_X1 _34177_ (.A(\bp_fe_pc_gen_1.pc_resume_r [26]),
    .ZN(_08599_));
 OAI21_X1 _34178_ (.A(_08598_),
    .B1(_08599_),
    .B2(_08587_),
    .ZN(_00706_));
 BUF_X32 _34179_ (.A(fe_cmd_i[61]),
    .Z(_08600_));
 AOI22_X1 _34180_ (.A1(_08570_),
    .A2(\bp_fe_pc_gen_1.pc_if2_r [27]),
    .B1(_08600_),
    .B2(_08572_),
    .ZN(_08601_));
 INV_X1 _34181_ (.A(\bp_fe_pc_gen_1.pc_resume_r [27]),
    .ZN(_08602_));
 OAI21_X1 _34182_ (.A(_08601_),
    .B1(_08602_),
    .B2(_08587_),
    .ZN(_00707_));
 BUF_X4 _34183_ (.A(_08522_),
    .Z(_08603_));
 BUF_X32 _34184_ (.A(fe_cmd_i[62]),
    .Z(_08604_));
 BUF_X4 _34185_ (.A(_08511_),
    .Z(_08605_));
 AOI22_X1 _34186_ (.A1(_08603_),
    .A2(\bp_fe_pc_gen_1.pc_if2_r [28]),
    .B1(_08604_),
    .B2(_08605_),
    .ZN(_08606_));
 INV_X1 _34187_ (.A(\bp_fe_pc_gen_1.pc_resume_r [28]),
    .ZN(_08607_));
 OAI21_X1 _34188_ (.A(_08606_),
    .B1(_08607_),
    .B2(_08587_),
    .ZN(_00708_));
 BUF_X32 _34189_ (.A(fe_cmd_i[63]),
    .Z(_08608_));
 AOI22_X1 _34190_ (.A1(_08603_),
    .A2(\bp_fe_pc_gen_1.pc_if2_r [29]),
    .B1(_08608_),
    .B2(_08605_),
    .ZN(_08609_));
 INV_X1 _34191_ (.A(\bp_fe_pc_gen_1.pc_resume_r [29]),
    .ZN(_08610_));
 OAI21_X1 _34192_ (.A(_08609_),
    .B1(_08610_),
    .B2(_08587_),
    .ZN(_00709_));
 BUF_X32 _34193_ (.A(fe_cmd_i[64]),
    .Z(_08611_));
 AOI22_X1 _34194_ (.A1(_08603_),
    .A2(\bp_fe_pc_gen_1.pc_if2_r [30]),
    .B1(_08611_),
    .B2(_08605_),
    .ZN(_08612_));
 INV_X1 _34195_ (.A(\bp_fe_pc_gen_1.pc_resume_r [30]),
    .ZN(_08613_));
 OAI21_X1 _34196_ (.A(_08612_),
    .B1(_08613_),
    .B2(_08587_),
    .ZN(_00711_));
 BUF_X32 _34197_ (.A(fe_cmd_i[65]),
    .Z(_08614_));
 AOI22_X1 _34198_ (.A1(_08603_),
    .A2(\bp_fe_pc_gen_1.pc_if2_r [31]),
    .B1(_08614_),
    .B2(_08605_),
    .ZN(_08615_));
 INV_X1 _34199_ (.A(\bp_fe_pc_gen_1.pc_resume_r [31]),
    .ZN(_08616_));
 OAI21_X1 _34200_ (.A(_08615_),
    .B1(_08616_),
    .B2(_08587_),
    .ZN(_00712_));
 BUF_X32 _34201_ (.A(fe_cmd_i[66]),
    .Z(_08617_));
 AOI22_X1 _34202_ (.A1(_08603_),
    .A2(\bp_fe_pc_gen_1.pc_if2_r [32]),
    .B1(_08617_),
    .B2(_08605_),
    .ZN(_08618_));
 INV_X1 _34203_ (.A(\bp_fe_pc_gen_1.pc_resume_r [32]),
    .ZN(_08619_));
 OAI21_X1 _34204_ (.A(_08618_),
    .B1(_08619_),
    .B2(_08543_),
    .ZN(_00713_));
 BUF_X32 _34205_ (.A(fe_cmd_i[67]),
    .Z(_08620_));
 AOI22_X1 _34206_ (.A1(_08603_),
    .A2(\bp_fe_pc_gen_1.pc_if2_r [33]),
    .B1(_08620_),
    .B2(_08605_),
    .ZN(_08621_));
 INV_X1 _34207_ (.A(\bp_fe_pc_gen_1.pc_resume_r [33]),
    .ZN(_08622_));
 OAI21_X1 _34208_ (.A(_08621_),
    .B1(_08622_),
    .B2(_08543_),
    .ZN(_00714_));
 BUF_X32 _34209_ (.A(fe_cmd_i[68]),
    .Z(_08623_));
 AOI22_X1 _34210_ (.A1(_08603_),
    .A2(\bp_fe_pc_gen_1.pc_if2_r [34]),
    .B1(_08623_),
    .B2(_08605_),
    .ZN(_08624_));
 INV_X1 _34211_ (.A(\bp_fe_pc_gen_1.pc_resume_r [34]),
    .ZN(_08625_));
 OAI21_X1 _34212_ (.A(_08624_),
    .B1(_08625_),
    .B2(_08543_),
    .ZN(_00715_));
 BUF_X32 _34213_ (.A(fe_cmd_i[69]),
    .Z(_08626_));
 AOI22_X1 _34214_ (.A1(_08603_),
    .A2(\bp_fe_pc_gen_1.pc_if2_r [35]),
    .B1(_08626_),
    .B2(_08605_),
    .ZN(_08627_));
 INV_X1 _34215_ (.A(\bp_fe_pc_gen_1.pc_resume_r [35]),
    .ZN(_08628_));
 OAI21_X1 _34216_ (.A(_08627_),
    .B1(_08628_),
    .B2(_08543_),
    .ZN(_00716_));
 BUF_X32 _34217_ (.A(fe_cmd_i[70]),
    .Z(_08629_));
 AOI22_X1 _34218_ (.A1(_08603_),
    .A2(\bp_fe_pc_gen_1.pc_if2_r [36]),
    .B1(_08629_),
    .B2(_08605_),
    .ZN(_08630_));
 INV_X1 _34219_ (.A(\bp_fe_pc_gen_1.pc_resume_r [36]),
    .ZN(_08631_));
 OAI21_X1 _34220_ (.A(_08630_),
    .B1(_08631_),
    .B2(_08543_),
    .ZN(_00717_));
 BUF_X32 _34221_ (.A(fe_cmd_i[71]),
    .Z(_08632_));
 AOI22_X1 _34222_ (.A1(_08603_),
    .A2(\bp_fe_pc_gen_1.pc_if2_r [37]),
    .B1(_08632_),
    .B2(_08605_),
    .ZN(_08633_));
 INV_X1 _34223_ (.A(\bp_fe_pc_gen_1.pc_resume_r [37]),
    .ZN(_08634_));
 OAI21_X1 _34224_ (.A(_08633_),
    .B1(_08634_),
    .B2(_08543_),
    .ZN(_00718_));
 BUF_X32 _34225_ (.A(fe_cmd_i[72]),
    .Z(_08635_));
 AOI22_X1 _34226_ (.A1(_08522_),
    .A2(\bp_fe_pc_gen_1.pc_if2_r [38]),
    .B1(_08635_),
    .B2(_08511_),
    .ZN(_08636_));
 INV_X1 _34227_ (.A(\bp_fe_pc_gen_1.pc_resume_r [38]),
    .ZN(_08637_));
 OAI21_X1 _34228_ (.A(_08636_),
    .B1(_08637_),
    .B2(_08543_),
    .ZN(_00719_));
 AOI21_X4 _34229_ (.A(_00080_),
    .B1(_00079_),
    .B2(_00078_),
    .ZN(_08638_));
 AND2_X1 _34230_ (.A1(\bp_fe_pc_gen_1.pc_v_if2_r ),
    .A2(\bp_fe_pc_gen_1.itlb_miss_if2_r ),
    .ZN(_08639_));
 NOR2_X4 _34231_ (.A1(_08638_),
    .A2(_08639_),
    .ZN(_08640_));
 OAI21_X4 _34232_ (.A(_08640_),
    .B1(\icache.N8 ),
    .B2(\icache.N7 ),
    .ZN(_08641_));
 AND2_X2 _34233_ (.A1(_08641_),
    .A2(\bp_fe_pc_gen_1.pc_v_if2_r ),
    .ZN(_08642_));
 BUF_X16 _34234_ (.A(_08642_),
    .Z(_08643_));
 BUF_X16 _34235_ (.A(_08643_),
    .Z(_08644_));
 BUF_X32 _34236_ (.A(_08644_),
    .Z(fe_queue_o[99]));
 INV_X1 _34237_ (.A(_08513_),
    .ZN(_08645_));
 OR3_X2 _34238_ (.A1(_08645_),
    .A2(_00080_),
    .A3(\bp_fe_pc_gen_1.itlb_miss_if2_r ),
    .ZN(_08646_));
 INV_X8 _34239_ (.A(_08643_),
    .ZN(_08647_));
 NAND2_X4 _34240_ (.A1(_08646_),
    .A2(_08647_),
    .ZN(_08648_));
 BUF_X4 _34241_ (.A(fe_queue_ready_i),
    .Z(_08649_));
 AND2_X4 _34242_ (.A1(_08648_),
    .A2(_08649_),
    .ZN(fe_queue_v_o));
 BUF_X16 _34243_ (.A(_08516_),
    .Z(_08650_));
 BUF_X8 _34244_ (.A(_08650_),
    .Z(_08651_));
 AOI21_X4 _34245_ (.A(_00080_),
    .B1(_08648_),
    .B2(fe_queue_ready_i),
    .ZN(_08652_));
 OAI21_X4 _34246_ (.A(_08512_),
    .B1(_08652_),
    .B2(_08643_),
    .ZN(_08653_));
 AND2_X1 _34247_ (.A1(_08653_),
    .A2(_08337_),
    .ZN(_08654_));
 NOR4_X4 _34248_ (.A1(_08026_),
    .A2(\bp_fe_pc_gen_1.state_r [0]),
    .A3(_08335_),
    .A4(_08035_),
    .ZN(_08655_));
 NOR2_X2 _34249_ (.A1(_08654_),
    .A2(_08655_),
    .ZN(_08656_));
 BUF_X8 _34250_ (.A(_08656_),
    .Z(_08657_));
 BUF_X8 _34251_ (.A(_08657_),
    .Z(_08658_));
 NOR2_X1 _34252_ (.A1(_08658_),
    .A2(\bp_fe_pc_gen_1.N79 ),
    .ZN(_08659_));
 INV_X2 _34253_ (.A(\bp_fe_pc_gen_1.pc_if2_r [0]),
    .ZN(_08660_));
 BUF_X8 _34254_ (.A(_08658_),
    .Z(_08661_));
 AOI211_X1 _34255_ (.A(_08651_),
    .B(_08659_),
    .C1(_08660_),
    .C2(_08661_),
    .ZN(_00649_));
 BUF_X8 _34256_ (.A(_08519_),
    .Z(_08662_));
 INV_X1 _34257_ (.A(_08656_),
    .ZN(_08663_));
 BUF_X8 _34258_ (.A(_08663_),
    .Z(_08664_));
 BUF_X8 _34259_ (.A(_08664_),
    .Z(_08665_));
 OAI21_X1 _34260_ (.A(_08662_),
    .B1(_08665_),
    .B2(\bp_fe_pc_gen_1.pc_if2_r [1]),
    .ZN(_08666_));
 INV_X1 _34261_ (.A(\bp_fe_pc_gen_1.N80 ),
    .ZN(_08667_));
 BUF_X8 _34262_ (.A(_08664_),
    .Z(_08668_));
 AOI21_X1 _34263_ (.A(_08666_),
    .B1(_08667_),
    .B2(_08668_),
    .ZN(_00660_));
 BUF_X4 _34264_ (.A(_08663_),
    .Z(_08669_));
 OAI21_X1 _34265_ (.A(_08662_),
    .B1(_08669_),
    .B2(\bp_fe_pc_gen_1.pc_if2_r [2]),
    .ZN(_08670_));
 INV_X1 _34266_ (.A(\bp_fe_pc_gen_1.pc_if1_r [2]),
    .ZN(_08671_));
 AOI21_X1 _34267_ (.A(_08670_),
    .B1(_08671_),
    .B2(_08668_),
    .ZN(_00671_));
 BUF_X8 _34268_ (.A(_08657_),
    .Z(_08672_));
 MUX2_X1 _34269_ (.A(\bp_fe_pc_gen_1.pc_if1_r [3]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [3]),
    .S(_08672_),
    .Z(_08673_));
 BUF_X16 _34270_ (.A(_08519_),
    .Z(_08674_));
 BUF_X8 _34271_ (.A(_08674_),
    .Z(_08675_));
 AND2_X1 _34272_ (.A1(_08673_),
    .A2(_08675_),
    .ZN(_00681_));
 MUX2_X1 _34273_ (.A(\bp_fe_pc_gen_1.pc_if1_r [4]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [4]),
    .S(_08672_),
    .Z(_08676_));
 AND2_X1 _34274_ (.A1(_08676_),
    .A2(_08675_),
    .ZN(_00682_));
 MUX2_X1 _34275_ (.A(\bp_fe_pc_gen_1.pc_if1_r [5]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [5]),
    .S(_08672_),
    .Z(_08677_));
 AND2_X1 _34276_ (.A1(_08677_),
    .A2(_08675_),
    .ZN(_00683_));
 MUX2_X1 _34277_ (.A(\bp_fe_pc_gen_1.pc_if1_r [6]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [6]),
    .S(_08672_),
    .Z(_08678_));
 AND2_X1 _34278_ (.A1(_08678_),
    .A2(_08675_),
    .ZN(_00684_));
 MUX2_X1 _34279_ (.A(\bp_fe_pc_gen_1.pc_if1_r [7]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [7]),
    .S(_08672_),
    .Z(_08679_));
 AND2_X1 _34280_ (.A1(_08679_),
    .A2(_08675_),
    .ZN(_00685_));
 BUF_X8 _34281_ (.A(_08656_),
    .Z(_08680_));
 MUX2_X1 _34282_ (.A(\bp_fe_pc_gen_1.pc_if1_r [8]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [8]),
    .S(_08680_),
    .Z(_08681_));
 AND2_X1 _34283_ (.A1(_08681_),
    .A2(_08675_),
    .ZN(_00686_));
 OAI21_X1 _34284_ (.A(_08662_),
    .B1(_08669_),
    .B2(\bp_fe_pc_gen_1.pc_if2_r [9]),
    .ZN(_08682_));
 AOI21_X1 _34285_ (.A(_08682_),
    .B1(_08386_),
    .B2(_08668_),
    .ZN(_00687_));
 MUX2_X1 _34286_ (.A(\bp_fe_pc_gen_1.pc_if1_r [10]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [10]),
    .S(_08680_),
    .Z(_08683_));
 AND2_X1 _34287_ (.A1(_08683_),
    .A2(_08675_),
    .ZN(_00650_));
 MUX2_X1 _34288_ (.A(\bp_fe_pc_gen_1.pc_if1_r [11]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [11]),
    .S(_08680_),
    .Z(_08684_));
 AND2_X1 _34289_ (.A1(_08684_),
    .A2(_08675_),
    .ZN(_00651_));
 MUX2_X1 _34290_ (.A(\bp_fe_pc_gen_1.pc_if1_r [12]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [12]),
    .S(_08680_),
    .Z(_08685_));
 AND2_X1 _34291_ (.A1(_08685_),
    .A2(_08675_),
    .ZN(_00652_));
 OAI21_X1 _34292_ (.A(_08662_),
    .B1(_08669_),
    .B2(\bp_fe_pc_gen_1.pc_if2_r [13]),
    .ZN(_08686_));
 INV_X1 _34293_ (.A(\bp_fe_pc_gen_1.pc_if1_r [13]),
    .ZN(_08687_));
 AOI21_X1 _34294_ (.A(_08686_),
    .B1(_08687_),
    .B2(_08668_),
    .ZN(_00653_));
 MUX2_X1 _34295_ (.A(\bp_fe_pc_gen_1.pc_if1_r [14]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [14]),
    .S(_08680_),
    .Z(_08688_));
 BUF_X8 _34296_ (.A(_08674_),
    .Z(_08689_));
 AND2_X1 _34297_ (.A1(_08688_),
    .A2(_08689_),
    .ZN(_00654_));
 OAI21_X1 _34298_ (.A(_08662_),
    .B1(_08669_),
    .B2(\bp_fe_pc_gen_1.pc_if2_r [15]),
    .ZN(_08690_));
 INV_X1 _34299_ (.A(\bp_fe_pc_gen_1.pc_if1_r [15]),
    .ZN(_08691_));
 AOI21_X1 _34300_ (.A(_08690_),
    .B1(_08691_),
    .B2(_08668_),
    .ZN(_00655_));
 MUX2_X1 _34301_ (.A(\bp_fe_pc_gen_1.pc_if1_r [16]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [16]),
    .S(_08680_),
    .Z(_08692_));
 AND2_X1 _34302_ (.A1(_08692_),
    .A2(_08689_),
    .ZN(_00656_));
 BUF_X4 _34303_ (.A(_08519_),
    .Z(_08693_));
 OAI21_X1 _34304_ (.A(_08693_),
    .B1(_08669_),
    .B2(\bp_fe_pc_gen_1.pc_if2_r [17]),
    .ZN(_08694_));
 INV_X1 _34305_ (.A(\bp_fe_pc_gen_1.pc_if1_r [17]),
    .ZN(_08695_));
 AOI21_X1 _34306_ (.A(_08694_),
    .B1(_08695_),
    .B2(_08668_),
    .ZN(_00657_));
 MUX2_X1 _34307_ (.A(\bp_fe_pc_gen_1.pc_if1_r [18]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [18]),
    .S(_08680_),
    .Z(_08696_));
 AND2_X1 _34308_ (.A1(_08696_),
    .A2(_08689_),
    .ZN(_00658_));
 OAI21_X1 _34309_ (.A(_08693_),
    .B1(_08669_),
    .B2(\bp_fe_pc_gen_1.pc_if2_r [19]),
    .ZN(_08697_));
 INV_X1 _34310_ (.A(\bp_fe_pc_gen_1.pc_if1_r [19]),
    .ZN(_08698_));
 AOI21_X1 _34311_ (.A(_08697_),
    .B1(_08698_),
    .B2(_08668_),
    .ZN(_00659_));
 MUX2_X1 _34312_ (.A(\bp_fe_pc_gen_1.pc_if1_r [20]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [20]),
    .S(_08680_),
    .Z(_08699_));
 AND2_X1 _34313_ (.A1(_08699_),
    .A2(_08689_),
    .ZN(_00661_));
 OAI21_X1 _34314_ (.A(_08693_),
    .B1(_08669_),
    .B2(\bp_fe_pc_gen_1.pc_if2_r [21]),
    .ZN(_08700_));
 INV_X1 _34315_ (.A(\bp_fe_pc_gen_1.pc_if1_r [21]),
    .ZN(_08701_));
 AOI21_X1 _34316_ (.A(_08700_),
    .B1(_08701_),
    .B2(_08668_),
    .ZN(_00662_));
 MUX2_X1 _34317_ (.A(\bp_fe_pc_gen_1.pc_if1_r [22]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [22]),
    .S(_08680_),
    .Z(_08702_));
 AND2_X1 _34318_ (.A1(_08702_),
    .A2(_08689_),
    .ZN(_00663_));
 OAI21_X1 _34319_ (.A(_08693_),
    .B1(_08669_),
    .B2(\bp_fe_pc_gen_1.pc_if2_r [23]),
    .ZN(_08703_));
 INV_X1 _34320_ (.A(\bp_fe_pc_gen_1.pc_if1_r [23]),
    .ZN(_08704_));
 AOI21_X1 _34321_ (.A(_08703_),
    .B1(_08704_),
    .B2(_08668_),
    .ZN(_00664_));
 MUX2_X1 _34322_ (.A(\bp_fe_pc_gen_1.pc_if1_r [24]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [24]),
    .S(_08680_),
    .Z(_08705_));
 AND2_X1 _34323_ (.A1(_08705_),
    .A2(_08689_),
    .ZN(_00665_));
 OAI21_X1 _34324_ (.A(_08693_),
    .B1(_08669_),
    .B2(\bp_fe_pc_gen_1.pc_if2_r [25]),
    .ZN(_08706_));
 INV_X1 _34325_ (.A(\bp_fe_pc_gen_1.pc_if1_r [25]),
    .ZN(_08707_));
 AOI21_X1 _34326_ (.A(_08706_),
    .B1(_08707_),
    .B2(_08668_),
    .ZN(_00666_));
 MUX2_X1 _34327_ (.A(\bp_fe_pc_gen_1.pc_if1_r [26]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [26]),
    .S(_08657_),
    .Z(_08708_));
 AND2_X1 _34328_ (.A1(_08708_),
    .A2(_08689_),
    .ZN(_00667_));
 OAI21_X1 _34329_ (.A(_08693_),
    .B1(_08669_),
    .B2(\bp_fe_pc_gen_1.pc_if2_r [27]),
    .ZN(_08709_));
 INV_X1 _34330_ (.A(\bp_fe_pc_gen_1.pc_if1_r [27]),
    .ZN(_08710_));
 BUF_X4 _34331_ (.A(_08664_),
    .Z(_08711_));
 AOI21_X1 _34332_ (.A(_08709_),
    .B1(_08710_),
    .B2(_08711_),
    .ZN(_00668_));
 MUX2_X1 _34333_ (.A(\bp_fe_pc_gen_1.pc_if1_r [28]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [28]),
    .S(_08657_),
    .Z(_08712_));
 AND2_X1 _34334_ (.A1(_08712_),
    .A2(_08689_),
    .ZN(_00669_));
 OAI21_X1 _34335_ (.A(_08693_),
    .B1(_08664_),
    .B2(\bp_fe_pc_gen_1.pc_if2_r [29]),
    .ZN(_08713_));
 INV_X1 _34336_ (.A(\bp_fe_pc_gen_1.pc_if1_r [29]),
    .ZN(_08714_));
 AOI21_X1 _34337_ (.A(_08713_),
    .B1(_08714_),
    .B2(_08711_),
    .ZN(_00670_));
 MUX2_X1 _34338_ (.A(\bp_fe_pc_gen_1.pc_if1_r [30]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [30]),
    .S(_08657_),
    .Z(_08715_));
 AND2_X1 _34339_ (.A1(_08715_),
    .A2(_08689_),
    .ZN(_00672_));
 OAI21_X1 _34340_ (.A(_08693_),
    .B1(_08664_),
    .B2(\bp_fe_pc_gen_1.pc_if2_r [31]),
    .ZN(_08716_));
 INV_X1 _34341_ (.A(\bp_fe_pc_gen_1.pc_if1_r [31]),
    .ZN(_08717_));
 AOI21_X1 _34342_ (.A(_08716_),
    .B1(_08717_),
    .B2(_08711_),
    .ZN(_00673_));
 MUX2_X1 _34343_ (.A(\bp_fe_pc_gen_1.pc_if1_r [32]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [32]),
    .S(_08657_),
    .Z(_08718_));
 AND2_X1 _34344_ (.A1(_08718_),
    .A2(_08689_),
    .ZN(_00674_));
 OAI21_X1 _34345_ (.A(_08693_),
    .B1(_08664_),
    .B2(\bp_fe_pc_gen_1.pc_if2_r [33]),
    .ZN(_08719_));
 INV_X1 _34346_ (.A(\bp_fe_pc_gen_1.pc_if1_r [33]),
    .ZN(_08720_));
 AOI21_X1 _34347_ (.A(_08719_),
    .B1(_08720_),
    .B2(_08711_),
    .ZN(_00675_));
 MUX2_X1 _34348_ (.A(\bp_fe_pc_gen_1.pc_if1_r [34]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [34]),
    .S(_08657_),
    .Z(_08721_));
 BUF_X8 _34349_ (.A(_08519_),
    .Z(_08722_));
 BUF_X8 _34350_ (.A(_08722_),
    .Z(_08723_));
 AND2_X1 _34351_ (.A1(_08721_),
    .A2(_08723_),
    .ZN(_00676_));
 OAI21_X1 _34352_ (.A(_08693_),
    .B1(_08664_),
    .B2(\bp_fe_pc_gen_1.pc_if2_r [35]),
    .ZN(_08724_));
 INV_X1 _34353_ (.A(\bp_fe_pc_gen_1.pc_if1_r [35]),
    .ZN(_08725_));
 AOI21_X1 _34354_ (.A(_08724_),
    .B1(_08725_),
    .B2(_08711_),
    .ZN(_00677_));
 MUX2_X1 _34355_ (.A(\bp_fe_pc_gen_1.pc_if1_r [36]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [36]),
    .S(_08657_),
    .Z(_08726_));
 AND2_X1 _34356_ (.A1(_08726_),
    .A2(_08723_),
    .ZN(_00678_));
 BUF_X8 _34357_ (.A(_08519_),
    .Z(_08727_));
 OAI21_X1 _34358_ (.A(_08727_),
    .B1(_08664_),
    .B2(\bp_fe_pc_gen_1.pc_if2_r [37]),
    .ZN(_08728_));
 INV_X2 _34359_ (.A(\bp_fe_pc_gen_1.pc_if1_r [37]),
    .ZN(_08729_));
 AOI21_X1 _34360_ (.A(_08728_),
    .B1(_08729_),
    .B2(_08711_),
    .ZN(_00679_));
 MUX2_X1 _34361_ (.A(\bp_fe_pc_gen_1.pc_if1_r [38]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [38]),
    .S(_08657_),
    .Z(_08730_));
 AND2_X1 _34362_ (.A1(_08730_),
    .A2(_08723_),
    .ZN(_00680_));
 BUF_X4 _34363_ (.A(_08655_),
    .Z(_08731_));
 BUF_X4 _34364_ (.A(_08653_),
    .Z(_08732_));
 AOI211_X1 _34365_ (.A(\bp_fe_pc_gen_1.N79 ),
    .B(_08731_),
    .C1(_08732_),
    .C2(_08533_),
    .ZN(_08733_));
 AND2_X1 _34366_ (.A1(_08371_),
    .A2(_08341_),
    .ZN(_08734_));
 INV_X4 _34367_ (.A(_08334_),
    .ZN(_08735_));
 AOI22_X2 _34368_ (.A1(_08734_),
    .A2(net1417),
    .B1(fe_cmd_i[34]),
    .B2(_08735_),
    .ZN(_08736_));
 AOI22_X1 _34369_ (.A1(_08409_),
    .A2(\bp_fe_pc_gen_1.N79 ),
    .B1(\bp_fe_pc_gen_1.pc_resume_r [0]),
    .B2(_08345_),
    .ZN(_08737_));
 AND2_X1 _34370_ (.A1(_08736_),
    .A2(_08737_),
    .ZN(_08738_));
 AOI211_X1 _34371_ (.A(_08651_),
    .B(_08733_),
    .C1(_08738_),
    .C2(_08711_),
    .ZN(_00610_));
 NOR3_X1 _34372_ (.A1(_08371_),
    .A2(_08667_),
    .A3(_08354_),
    .ZN(_08739_));
 AOI221_X4 _34373_ (.A(_08739_),
    .B1(fe_cmd_i[35]),
    .B2(_08735_),
    .C1(\bp_fe_pc_gen_1.pc_resume_r [1]),
    .C2(_08345_),
    .ZN(_08740_));
 NAND4_X4 _34374_ (.A1(_08451_),
    .A2(net1416),
    .A3(_08341_),
    .A4(_08469_),
    .ZN(_08741_));
 AND3_X1 _34375_ (.A1(_08740_),
    .A2(_08664_),
    .A3(_08741_),
    .ZN(_08742_));
 AOI211_X1 _34376_ (.A(_08651_),
    .B(_08742_),
    .C1(_08667_),
    .C2(_08661_),
    .ZN(_00621_));
 NOR2_X2 _34377_ (.A1(_08350_),
    .A2(_08536_),
    .ZN(_08743_));
 NAND2_X1 _34378_ (.A1(_08321_),
    .A2(_08340_),
    .ZN(_08744_));
 OR2_X1 _34379_ (.A1(_08744_),
    .A2(_00082_),
    .ZN(_08745_));
 OR3_X1 _34380_ (.A1(_08321_),
    .A2(\bp_fe_pc_gen_1.pc_if1_r [2]),
    .A3(_08354_),
    .ZN(_08746_));
 NAND3_X1 _34381_ (.A1(_08745_),
    .A2(_08348_),
    .A3(_08746_),
    .ZN(_08747_));
 NAND3_X1 _34382_ (.A1(_08334_),
    .A2(_00081_),
    .A3(_08344_),
    .ZN(_08748_));
 AOI211_X1 _34383_ (.A(_08672_),
    .B(_08743_),
    .C1(_08747_),
    .C2(_08748_),
    .ZN(_08749_));
 AOI211_X1 _34384_ (.A(_08651_),
    .B(_08749_),
    .C1(_08671_),
    .C2(_08661_),
    .ZN(_00632_));
 BUF_X4 _34385_ (.A(_08337_),
    .Z(_08750_));
 AOI211_X1 _34386_ (.A(\bp_fe_pc_gen_1.pc_if1_r [3]),
    .B(_08731_),
    .C1(_08732_),
    .C2(_08750_),
    .ZN(_08751_));
 AND2_X1 _34387_ (.A1(_08475_),
    .A2(_08478_),
    .ZN(_08752_));
 AOI211_X1 _34388_ (.A(_08651_),
    .B(_08751_),
    .C1(_08752_),
    .C2(_08711_),
    .ZN(_00642_));
 BUF_X4 _34389_ (.A(_08650_),
    .Z(_08753_));
 AOI211_X1 _34390_ (.A(\bp_fe_pc_gen_1.pc_if1_r [4]),
    .B(_08731_),
    .C1(_08732_),
    .C2(_08750_),
    .ZN(_08754_));
 NOR2_X4 _34391_ (.A1(_08436_),
    .A2(_08440_),
    .ZN(_08755_));
 AOI211_X1 _34392_ (.A(_08753_),
    .B(_08754_),
    .C1(_08755_),
    .C2(_08711_),
    .ZN(_00643_));
 AOI211_X1 _34393_ (.A(\bp_fe_pc_gen_1.pc_if1_r [5]),
    .B(_08731_),
    .C1(_08732_),
    .C2(_08750_),
    .ZN(_08756_));
 NOR2_X4 _34394_ (.A1(_08413_),
    .A2(_08417_),
    .ZN(_08757_));
 AOI211_X1 _34395_ (.A(_08753_),
    .B(_08756_),
    .C1(_08757_),
    .C2(_08711_),
    .ZN(_00644_));
 AOI211_X1 _34396_ (.A(\bp_fe_pc_gen_1.pc_if1_r [6]),
    .B(_08731_),
    .C1(_08732_),
    .C2(_08750_),
    .ZN(_08758_));
 NOR2_X4 _34397_ (.A1(_08351_),
    .A2(_08358_),
    .ZN(_08759_));
 BUF_X8 _34398_ (.A(_08664_),
    .Z(_08760_));
 AOI211_X1 _34399_ (.A(_08753_),
    .B(_08758_),
    .C1(_08759_),
    .C2(_08760_),
    .ZN(_00645_));
 AOI211_X1 _34400_ (.A(\bp_fe_pc_gen_1.pc_if1_r [7]),
    .B(_08731_),
    .C1(_08732_),
    .C2(_08750_),
    .ZN(_08761_));
 NOR2_X4 _34401_ (.A1(_08365_),
    .A2(_08368_),
    .ZN(_08762_));
 AOI211_X1 _34402_ (.A(_08753_),
    .B(_08761_),
    .C1(_08762_),
    .C2(_08760_),
    .ZN(_00646_));
 AOI211_X1 _34403_ (.A(\bp_fe_pc_gen_1.pc_if1_r [8]),
    .B(_08731_),
    .C1(_08732_),
    .C2(_08750_),
    .ZN(_08763_));
 NOR2_X2 _34404_ (.A1(_08375_),
    .A2(_08378_),
    .ZN(_08764_));
 AOI211_X1 _34405_ (.A(_08753_),
    .B(_08763_),
    .C1(_08764_),
    .C2(_08760_),
    .ZN(_00647_));
 NOR3_X1 _34406_ (.A1(_08384_),
    .A2(_08388_),
    .A3(_08672_),
    .ZN(_08765_));
 AOI211_X1 _34407_ (.A(_08753_),
    .B(_08765_),
    .C1(_08386_),
    .C2(_08661_),
    .ZN(_00648_));
 AOI211_X1 _34408_ (.A(\bp_fe_pc_gen_1.pc_if1_r [10]),
    .B(_08731_),
    .C1(_08732_),
    .C2(_08750_),
    .ZN(_08766_));
 NOR2_X2 _34409_ (.A1(_08394_),
    .A2(_08397_),
    .ZN(_08767_));
 AOI211_X1 _34410_ (.A(_08753_),
    .B(_08766_),
    .C1(_08767_),
    .C2(_08760_),
    .ZN(_00611_));
 AOI211_X1 _34411_ (.A(\bp_fe_pc_gen_1.pc_if1_r [11]),
    .B(_08731_),
    .C1(_08732_),
    .C2(_08750_),
    .ZN(_08768_));
 NOR2_X2 _34412_ (.A1(_08403_),
    .A2(_08406_),
    .ZN(_08769_));
 AOI211_X1 _34413_ (.A(_08753_),
    .B(_08768_),
    .C1(_08769_),
    .C2(_08760_),
    .ZN(_00612_));
 AOI211_X1 _34414_ (.A(\bp_fe_pc_gen_1.pc_if1_r [12]),
    .B(_08731_),
    .C1(_08732_),
    .C2(_08750_),
    .ZN(_08770_));
 BUF_X8 _34415_ (.A(_08339_),
    .Z(_08771_));
 NAND3_X2 _34416_ (.A1(_08319_),
    .A2(\bp_fe_pc_gen_1.btb.br_tgt_o [12]),
    .A3(_08771_),
    .ZN(_08772_));
 BUF_X4 _34417_ (.A(_08331_),
    .Z(_08773_));
 BUF_X8 _34418_ (.A(_08333_),
    .Z(_08774_));
 OAI21_X2 _34419_ (.A(fe_cmd_i[46]),
    .B1(_08773_),
    .B2(_08774_),
    .ZN(_08775_));
 BUF_X8 _34420_ (.A(_08346_),
    .Z(_08776_));
 OAI211_X4 _34421_ (.A(_08772_),
    .B(_08775_),
    .C1(_08553_),
    .C2(_08776_),
    .ZN(_08777_));
 BUF_X8 _34422_ (.A(_08318_),
    .Z(_08778_));
 BUF_X8 _34423_ (.A(_08352_),
    .Z(_08779_));
 NAND2_X1 _34424_ (.A1(_08404_),
    .A2(\bp_fe_pc_gen_1.pc_if1_r [11]),
    .ZN(_08780_));
 XNOR2_X2 _34425_ (.A(_08780_),
    .B(_00083_),
    .ZN(_08781_));
 NOR3_X2 _34426_ (.A1(_08778_),
    .A2(_08779_),
    .A3(_08781_),
    .ZN(_08782_));
 NOR2_X4 _34427_ (.A1(_08777_),
    .A2(_08782_),
    .ZN(_08783_));
 BUF_X16 _34428_ (.A(_08783_),
    .Z(_08784_));
 AOI211_X1 _34429_ (.A(_08753_),
    .B(_08770_),
    .C1(_08784_),
    .C2(_08760_),
    .ZN(_00613_));
 BUF_X8 _34430_ (.A(_08318_),
    .Z(_08785_));
 BUF_X8 _34431_ (.A(_08785_),
    .Z(_08786_));
 NAND3_X2 _34432_ (.A1(_08786_),
    .A2(\bp_fe_pc_gen_1.btb.br_tgt_o [13]),
    .A3(_08340_),
    .ZN(_08787_));
 OAI21_X2 _34433_ (.A(fe_cmd_i[47]),
    .B1(_08476_),
    .B2(_08477_),
    .ZN(_08788_));
 OAI211_X4 _34434_ (.A(_08787_),
    .B(_08788_),
    .C1(_08557_),
    .C2(_08347_),
    .ZN(_08789_));
 BUF_X4 _34435_ (.A(_08657_),
    .Z(_08790_));
 AND3_X1 _34436_ (.A1(_08404_),
    .A2(\bp_fe_pc_gen_1.pc_if1_r [11]),
    .A3(\bp_fe_pc_gen_1.pc_if1_r [12]),
    .ZN(_08791_));
 XNOR2_X1 _34437_ (.A(_08791_),
    .B(\bp_fe_pc_gen_1.pc_if1_r [13]),
    .ZN(_08792_));
 NOR3_X2 _34438_ (.A1(_08320_),
    .A2(_08353_),
    .A3(_08792_),
    .ZN(_08793_));
 NOR3_X1 _34439_ (.A1(_08789_),
    .A2(_08790_),
    .A3(_08793_),
    .ZN(_08794_));
 AOI211_X1 _34440_ (.A(_08753_),
    .B(_08794_),
    .C1(_08687_),
    .C2(_08661_),
    .ZN(_00614_));
 BUF_X4 _34441_ (.A(_08650_),
    .Z(_08795_));
 BUF_X4 _34442_ (.A(_08655_),
    .Z(_08796_));
 BUF_X4 _34443_ (.A(_08653_),
    .Z(_08797_));
 AOI211_X1 _34444_ (.A(\bp_fe_pc_gen_1.pc_if1_r [14]),
    .B(_08796_),
    .C1(_08797_),
    .C2(_08750_),
    .ZN(_08798_));
 AND3_X1 _34445_ (.A1(_08318_),
    .A2(net1412),
    .A3(_08338_),
    .ZN(_08799_));
 AOI221_X2 _34446_ (.A(_08799_),
    .B1(fe_cmd_i[48]),
    .B2(_08735_),
    .C1(\bp_fe_pc_gen_1.pc_resume_r [14]),
    .C2(_08345_),
    .ZN(_08800_));
 NAND2_X1 _34447_ (.A1(_08791_),
    .A2(\bp_fe_pc_gen_1.pc_if1_r [13]),
    .ZN(_08801_));
 XNOR2_X2 _34448_ (.A(_08801_),
    .B(_00084_),
    .ZN(_08802_));
 OR3_X4 _34449_ (.A1(_08778_),
    .A2(_08779_),
    .A3(_08802_),
    .ZN(_08803_));
 AND2_X4 _34450_ (.A1(net212),
    .A2(_08803_),
    .ZN(_08804_));
 BUF_X16 _34451_ (.A(_08804_),
    .Z(_08805_));
 AOI211_X1 _34452_ (.A(_08795_),
    .B(_08798_),
    .C1(_08805_),
    .C2(_08760_),
    .ZN(_00615_));
 NAND3_X2 _34453_ (.A1(_08319_),
    .A2(net1411),
    .A3(_08771_),
    .ZN(_08806_));
 OAI21_X2 _34454_ (.A(fe_cmd_i[49]),
    .B1(_08773_),
    .B2(_08774_),
    .ZN(_08807_));
 OAI211_X4 _34455_ (.A(_08806_),
    .B(_08807_),
    .C1(_08563_),
    .C2(_08776_),
    .ZN(_08808_));
 AND3_X1 _34456_ (.A1(_08791_),
    .A2(\bp_fe_pc_gen_1.pc_if1_r [13]),
    .A3(\bp_fe_pc_gen_1.pc_if1_r [14]),
    .ZN(_08809_));
 XNOR2_X2 _34457_ (.A(_08809_),
    .B(\bp_fe_pc_gen_1.pc_if1_r [15]),
    .ZN(_08810_));
 NOR3_X4 _34458_ (.A1(_08786_),
    .A2(_08779_),
    .A3(_08810_),
    .ZN(_08811_));
 NOR3_X1 _34459_ (.A1(_08808_),
    .A2(_08790_),
    .A3(_08811_),
    .ZN(_08812_));
 AOI211_X1 _34460_ (.A(_08795_),
    .B(_08812_),
    .C1(_08691_),
    .C2(_08661_),
    .ZN(_00616_));
 BUF_X4 _34461_ (.A(_08337_),
    .Z(_08813_));
 AOI211_X1 _34462_ (.A(\bp_fe_pc_gen_1.pc_if1_r [16]),
    .B(_08796_),
    .C1(_08797_),
    .C2(_08813_),
    .ZN(_08814_));
 NAND3_X2 _34463_ (.A1(_08319_),
    .A2(net1410),
    .A3(_08771_),
    .ZN(_08815_));
 OAI21_X2 _34464_ (.A(fe_cmd_i[50]),
    .B1(_08773_),
    .B2(_08774_),
    .ZN(_08816_));
 OAI211_X4 _34465_ (.A(_08815_),
    .B(_08816_),
    .C1(_08566_),
    .C2(_08776_),
    .ZN(_08817_));
 NAND2_X1 _34466_ (.A1(_08809_),
    .A2(\bp_fe_pc_gen_1.pc_if1_r [15]),
    .ZN(_08818_));
 XNOR2_X2 _34467_ (.A(_08818_),
    .B(_00085_),
    .ZN(_08819_));
 NOR3_X2 _34468_ (.A1(_08786_),
    .A2(_08779_),
    .A3(_08819_),
    .ZN(_08820_));
 NOR2_X4 _34469_ (.A1(_08817_),
    .A2(_08820_),
    .ZN(_08821_));
 BUF_X16 _34470_ (.A(_08821_),
    .Z(_08822_));
 AOI211_X1 _34471_ (.A(_08795_),
    .B(_08814_),
    .C1(_08822_),
    .C2(_08760_),
    .ZN(_00617_));
 NAND3_X4 _34472_ (.A1(_08785_),
    .A2(\bp_fe_pc_gen_1.btb.br_tgt_o [17]),
    .A3(_08771_),
    .ZN(_08823_));
 OAI21_X2 _34473_ (.A(fe_cmd_i[51]),
    .B1(_08773_),
    .B2(_08774_),
    .ZN(_08824_));
 OAI211_X4 _34474_ (.A(_08823_),
    .B(_08824_),
    .C1(_08569_),
    .C2(_08776_),
    .ZN(_08825_));
 AND3_X2 _34475_ (.A1(_08809_),
    .A2(\bp_fe_pc_gen_1.pc_if1_r [15]),
    .A3(\bp_fe_pc_gen_1.pc_if1_r [16]),
    .ZN(_08826_));
 XNOR2_X1 _34476_ (.A(_08826_),
    .B(\bp_fe_pc_gen_1.pc_if1_r [17]),
    .ZN(_08827_));
 NOR3_X2 _34477_ (.A1(_08778_),
    .A2(_08779_),
    .A3(_08827_),
    .ZN(_08828_));
 NOR3_X1 _34478_ (.A1(_08825_),
    .A2(_08790_),
    .A3(_08828_),
    .ZN(_08829_));
 AOI211_X1 _34479_ (.A(_08795_),
    .B(_08829_),
    .C1(_08695_),
    .C2(_08661_),
    .ZN(_00618_));
 AOI211_X1 _34480_ (.A(\bp_fe_pc_gen_1.pc_if1_r [18]),
    .B(_08796_),
    .C1(_08797_),
    .C2(_08813_),
    .ZN(_08830_));
 NAND3_X2 _34481_ (.A1(_08320_),
    .A2(net1409),
    .A3(_08340_),
    .ZN(_08831_));
 OAI21_X2 _34482_ (.A(fe_cmd_i[52]),
    .B1(_08476_),
    .B2(_08477_),
    .ZN(_08832_));
 OAI211_X4 _34483_ (.A(_08831_),
    .B(_08832_),
    .C1(_08574_),
    .C2(_08347_),
    .ZN(_08833_));
 NAND2_X1 _34484_ (.A1(_08826_),
    .A2(\bp_fe_pc_gen_1.pc_if1_r [17]),
    .ZN(_08834_));
 XNOR2_X2 _34485_ (.A(_08834_),
    .B(_00086_),
    .ZN(_08835_));
 NOR3_X2 _34486_ (.A1(_08320_),
    .A2(_08353_),
    .A3(_08835_),
    .ZN(_08836_));
 NOR2_X4 _34487_ (.A1(_08833_),
    .A2(_08836_),
    .ZN(_08837_));
 BUF_X8 _34488_ (.A(_08837_),
    .Z(_08838_));
 AOI211_X1 _34489_ (.A(_08795_),
    .B(_08830_),
    .C1(_08838_),
    .C2(_08760_),
    .ZN(_00619_));
 NAND3_X2 _34490_ (.A1(_08778_),
    .A2(net1408),
    .A3(_08340_),
    .ZN(_08839_));
 OAI21_X2 _34491_ (.A(fe_cmd_i[53]),
    .B1(_08476_),
    .B2(_08477_),
    .ZN(_08840_));
 OAI211_X4 _34492_ (.A(_08839_),
    .B(_08840_),
    .C1(_08577_),
    .C2(_08347_),
    .ZN(_08841_));
 AND3_X1 _34493_ (.A1(_08826_),
    .A2(\bp_fe_pc_gen_1.pc_if1_r [17]),
    .A3(\bp_fe_pc_gen_1.pc_if1_r [18]),
    .ZN(_08842_));
 XNOR2_X2 _34494_ (.A(_08842_),
    .B(\bp_fe_pc_gen_1.pc_if1_r [19]),
    .ZN(_08843_));
 NOR3_X4 _34495_ (.A1(_08786_),
    .A2(_08353_),
    .A3(_08843_),
    .ZN(_08844_));
 NOR3_X1 _34496_ (.A1(_08841_),
    .A2(_08790_),
    .A3(_08844_),
    .ZN(_08845_));
 AOI211_X1 _34497_ (.A(_08795_),
    .B(_08845_),
    .C1(_08698_),
    .C2(_08661_),
    .ZN(_00620_));
 AOI211_X1 _34498_ (.A(\bp_fe_pc_gen_1.pc_if1_r [20]),
    .B(_08796_),
    .C1(_08797_),
    .C2(_08813_),
    .ZN(_08846_));
 AND3_X1 _34499_ (.A1(_08318_),
    .A2(\bp_fe_pc_gen_1.btb.br_tgt_o [20]),
    .A3(_08339_),
    .ZN(_08847_));
 AOI221_X2 _34500_ (.A(_08847_),
    .B1(fe_cmd_i[54]),
    .B2(_08735_),
    .C1(\bp_fe_pc_gen_1.pc_resume_r [20]),
    .C2(_08345_),
    .ZN(_08848_));
 NAND2_X1 _34501_ (.A1(_08842_),
    .A2(\bp_fe_pc_gen_1.pc_if1_r [19]),
    .ZN(_08849_));
 XNOR2_X1 _34502_ (.A(_08849_),
    .B(_00087_),
    .ZN(_08850_));
 OR3_X4 _34503_ (.A1(_08320_),
    .A2(_08353_),
    .A3(_08850_),
    .ZN(_08851_));
 AND2_X4 _34504_ (.A1(net210),
    .A2(_08851_),
    .ZN(_08852_));
 BUF_X8 _34505_ (.A(_08852_),
    .Z(_08853_));
 AOI211_X1 _34506_ (.A(_08795_),
    .B(_08846_),
    .C1(_08853_),
    .C2(_08760_),
    .ZN(_00622_));
 NAND3_X2 _34507_ (.A1(_08778_),
    .A2(net1407),
    .A3(_08340_),
    .ZN(_08854_));
 OAI21_X2 _34508_ (.A(fe_cmd_i[55]),
    .B1(_08476_),
    .B2(_08477_),
    .ZN(_08855_));
 OAI211_X4 _34509_ (.A(_08854_),
    .B(_08855_),
    .C1(_08583_),
    .C2(_08347_),
    .ZN(_08856_));
 AND3_X1 _34510_ (.A1(_08842_),
    .A2(\bp_fe_pc_gen_1.pc_if1_r [19]),
    .A3(\bp_fe_pc_gen_1.pc_if1_r [20]),
    .ZN(_08857_));
 XNOR2_X2 _34511_ (.A(_08857_),
    .B(\bp_fe_pc_gen_1.pc_if1_r [21]),
    .ZN(_08858_));
 NOR3_X2 _34512_ (.A1(_08320_),
    .A2(_08353_),
    .A3(_08858_),
    .ZN(_08859_));
 NOR3_X1 _34513_ (.A1(_08856_),
    .A2(_08790_),
    .A3(_08859_),
    .ZN(_08860_));
 AOI211_X1 _34514_ (.A(_08795_),
    .B(_08860_),
    .C1(_08701_),
    .C2(_08661_),
    .ZN(_00623_));
 AOI211_X1 _34515_ (.A(\bp_fe_pc_gen_1.pc_if1_r [22]),
    .B(_08796_),
    .C1(_08797_),
    .C2(_08813_),
    .ZN(_08861_));
 NAND3_X2 _34516_ (.A1(_08318_),
    .A2(net1406),
    .A3(_08339_),
    .ZN(_08862_));
 OAI21_X2 _34517_ (.A(fe_cmd_i[56]),
    .B1(_08331_),
    .B2(_08333_),
    .ZN(_08863_));
 OAI211_X4 _34518_ (.A(_08862_),
    .B(_08863_),
    .C1(_08586_),
    .C2(_08346_),
    .ZN(_08864_));
 NAND2_X1 _34519_ (.A1(_08857_),
    .A2(\bp_fe_pc_gen_1.pc_if1_r [21]),
    .ZN(_08865_));
 XNOR2_X1 _34520_ (.A(_08865_),
    .B(_00088_),
    .ZN(_08866_));
 NOR3_X2 _34521_ (.A1(_08785_),
    .A2(_08352_),
    .A3(_08866_),
    .ZN(_08867_));
 NOR2_X4 _34522_ (.A1(_08864_),
    .A2(_08867_),
    .ZN(_08868_));
 AOI211_X1 _34523_ (.A(_08795_),
    .B(_08861_),
    .C1(_08868_),
    .C2(_08665_),
    .ZN(_00624_));
 NAND3_X2 _34524_ (.A1(_08778_),
    .A2(\bp_fe_pc_gen_1.btb.br_tgt_o [23]),
    .A3(_08771_),
    .ZN(_08869_));
 OAI21_X2 _34525_ (.A(fe_cmd_i[57]),
    .B1(_08476_),
    .B2(_08477_),
    .ZN(_08870_));
 OAI211_X4 _34526_ (.A(_08869_),
    .B(_08870_),
    .C1(_08590_),
    .C2(_08347_),
    .ZN(_08871_));
 AND3_X1 _34527_ (.A1(_08857_),
    .A2(\bp_fe_pc_gen_1.pc_if1_r [21]),
    .A3(\bp_fe_pc_gen_1.pc_if1_r [22]),
    .ZN(_08872_));
 XNOR2_X2 _34528_ (.A(_08872_),
    .B(\bp_fe_pc_gen_1.pc_if1_r [23]),
    .ZN(_08873_));
 NOR3_X4 _34529_ (.A1(_08786_),
    .A2(_08353_),
    .A3(_08873_),
    .ZN(_08874_));
 NOR3_X1 _34530_ (.A1(_08871_),
    .A2(_08790_),
    .A3(_08874_),
    .ZN(_08875_));
 AOI211_X1 _34531_ (.A(_08795_),
    .B(_08875_),
    .C1(_08704_),
    .C2(_08658_),
    .ZN(_00625_));
 BUF_X4 _34532_ (.A(_08650_),
    .Z(_08876_));
 AOI211_X1 _34533_ (.A(\bp_fe_pc_gen_1.pc_if1_r [24]),
    .B(_08796_),
    .C1(_08797_),
    .C2(_08813_),
    .ZN(_08877_));
 NAND3_X2 _34534_ (.A1(_08778_),
    .A2(\bp_fe_pc_gen_1.btb.br_tgt_o [24]),
    .A3(_08340_),
    .ZN(_08878_));
 OAI21_X2 _34535_ (.A(fe_cmd_i[58]),
    .B1(_08476_),
    .B2(_08477_),
    .ZN(_08879_));
 OAI211_X4 _34536_ (.A(_08878_),
    .B(_08879_),
    .C1(_08593_),
    .C2(_08347_),
    .ZN(_08880_));
 NAND2_X1 _34537_ (.A1(_08872_),
    .A2(\bp_fe_pc_gen_1.pc_if1_r [23]),
    .ZN(_08881_));
 XNOR2_X2 _34538_ (.A(_08881_),
    .B(_00089_),
    .ZN(_08882_));
 NOR3_X2 _34539_ (.A1(_08320_),
    .A2(_08353_),
    .A3(_08882_),
    .ZN(_08883_));
 NOR2_X4 _34540_ (.A1(_08880_),
    .A2(_08883_),
    .ZN(_08884_));
 BUF_X8 _34541_ (.A(_08884_),
    .Z(_08885_));
 AOI211_X1 _34542_ (.A(_08876_),
    .B(_08877_),
    .C1(_08885_),
    .C2(_08665_),
    .ZN(_00626_));
 NAND3_X2 _34543_ (.A1(_08318_),
    .A2(\bp_fe_pc_gen_1.btb.br_tgt_o [25]),
    .A3(_08339_),
    .ZN(_08886_));
 OAI21_X2 _34544_ (.A(fe_cmd_i[59]),
    .B1(_08331_),
    .B2(_08333_),
    .ZN(_08887_));
 OAI211_X4 _34545_ (.A(_08886_),
    .B(_08887_),
    .C1(_08596_),
    .C2(_08346_),
    .ZN(_08888_));
 AND3_X1 _34546_ (.A1(_08872_),
    .A2(\bp_fe_pc_gen_1.pc_if1_r [23]),
    .A3(\bp_fe_pc_gen_1.pc_if1_r [24]),
    .ZN(_08889_));
 XNOR2_X1 _34547_ (.A(_08889_),
    .B(\bp_fe_pc_gen_1.pc_if1_r [25]),
    .ZN(_08890_));
 NOR3_X2 _34548_ (.A1(_08785_),
    .A2(_08352_),
    .A3(_08890_),
    .ZN(_08891_));
 NOR3_X1 _34549_ (.A1(_08888_),
    .A2(_08790_),
    .A3(_08891_),
    .ZN(_08892_));
 AOI211_X1 _34550_ (.A(_08876_),
    .B(_08892_),
    .C1(_08707_),
    .C2(_08658_),
    .ZN(_00627_));
 AOI211_X1 _34551_ (.A(\bp_fe_pc_gen_1.pc_if1_r [26]),
    .B(_08796_),
    .C1(_08797_),
    .C2(_08813_),
    .ZN(_08893_));
 NAND3_X2 _34552_ (.A1(_08320_),
    .A2(\bp_fe_pc_gen_1.btb.br_tgt_o [26]),
    .A3(_08340_),
    .ZN(_08894_));
 OAI21_X2 _34553_ (.A(fe_cmd_i[60]),
    .B1(_08476_),
    .B2(_08477_),
    .ZN(_08895_));
 OAI211_X4 _34554_ (.A(_08894_),
    .B(_08895_),
    .C1(_08599_),
    .C2(_08347_),
    .ZN(_08896_));
 NAND2_X1 _34555_ (.A1(_08889_),
    .A2(\bp_fe_pc_gen_1.pc_if1_r [25]),
    .ZN(_08897_));
 XNOR2_X2 _34556_ (.A(_08897_),
    .B(_00090_),
    .ZN(_08898_));
 NOR3_X4 _34557_ (.A1(_08320_),
    .A2(_08354_),
    .A3(_08898_),
    .ZN(_08899_));
 NOR2_X4 _34558_ (.A1(_08896_),
    .A2(_08899_),
    .ZN(_08900_));
 BUF_X8 _34559_ (.A(_08900_),
    .Z(_08901_));
 AOI211_X1 _34560_ (.A(_08876_),
    .B(_08893_),
    .C1(_08901_),
    .C2(_08665_),
    .ZN(_00628_));
 NAND3_X2 _34561_ (.A1(_08319_),
    .A2(\bp_fe_pc_gen_1.btb.br_tgt_o [27]),
    .A3(_08771_),
    .ZN(_08902_));
 OAI21_X2 _34562_ (.A(fe_cmd_i[61]),
    .B1(_08773_),
    .B2(_08774_),
    .ZN(_08903_));
 OAI211_X4 _34563_ (.A(_08902_),
    .B(_08903_),
    .C1(_08602_),
    .C2(_08776_),
    .ZN(_08904_));
 AND3_X1 _34564_ (.A1(_08889_),
    .A2(\bp_fe_pc_gen_1.pc_if1_r [25]),
    .A3(\bp_fe_pc_gen_1.pc_if1_r [26]),
    .ZN(_08905_));
 XNOR2_X1 _34565_ (.A(_08905_),
    .B(\bp_fe_pc_gen_1.pc_if1_r [27]),
    .ZN(_08906_));
 NOR3_X2 _34566_ (.A1(_08786_),
    .A2(_08779_),
    .A3(_08906_),
    .ZN(_08907_));
 NOR3_X1 _34567_ (.A1(_08904_),
    .A2(_08790_),
    .A3(_08907_),
    .ZN(_08908_));
 AOI211_X1 _34568_ (.A(_08876_),
    .B(_08908_),
    .C1(_08710_),
    .C2(_08658_),
    .ZN(_00629_));
 AOI211_X1 _34569_ (.A(\bp_fe_pc_gen_1.pc_if1_r [28]),
    .B(_08796_),
    .C1(_08797_),
    .C2(_08813_),
    .ZN(_08909_));
 NAND3_X2 _34570_ (.A1(_08785_),
    .A2(\bp_fe_pc_gen_1.btb.br_tgt_o [28]),
    .A3(_08339_),
    .ZN(_08910_));
 OAI21_X2 _34571_ (.A(fe_cmd_i[62]),
    .B1(_08773_),
    .B2(_08774_),
    .ZN(_08911_));
 OAI211_X4 _34572_ (.A(_08910_),
    .B(_08911_),
    .C1(_08607_),
    .C2(_08776_),
    .ZN(_08912_));
 NAND2_X1 _34573_ (.A1(_08905_),
    .A2(\bp_fe_pc_gen_1.pc_if1_r [27]),
    .ZN(_08913_));
 XNOR2_X1 _34574_ (.A(_08913_),
    .B(_00091_),
    .ZN(_08914_));
 NOR3_X2 _34575_ (.A1(_08319_),
    .A2(_08352_),
    .A3(_08914_),
    .ZN(_08915_));
 NOR2_X4 _34576_ (.A1(_08912_),
    .A2(_08915_),
    .ZN(_08916_));
 BUF_X8 _34577_ (.A(_08916_),
    .Z(_08917_));
 AOI211_X1 _34578_ (.A(_08876_),
    .B(_08909_),
    .C1(_08917_),
    .C2(_08665_),
    .ZN(_00630_));
 NAND3_X2 _34579_ (.A1(_08318_),
    .A2(\bp_fe_pc_gen_1.btb.br_tgt_o [29]),
    .A3(_08338_),
    .ZN(_08918_));
 OAI21_X2 _34580_ (.A(fe_cmd_i[63]),
    .B1(_08331_),
    .B2(_08333_),
    .ZN(_08919_));
 OAI211_X4 _34581_ (.A(_08918_),
    .B(_08919_),
    .C1(_08610_),
    .C2(_08346_),
    .ZN(_08920_));
 AND3_X1 _34582_ (.A1(_08905_),
    .A2(\bp_fe_pc_gen_1.pc_if1_r [27]),
    .A3(\bp_fe_pc_gen_1.pc_if1_r [28]),
    .ZN(_08921_));
 XNOR2_X2 _34583_ (.A(_08921_),
    .B(\bp_fe_pc_gen_1.pc_if1_r [29]),
    .ZN(_08922_));
 NOR3_X2 _34584_ (.A1(_08318_),
    .A2(_08352_),
    .A3(_08922_),
    .ZN(_08923_));
 NOR3_X1 _34585_ (.A1(_08920_),
    .A2(_08790_),
    .A3(_08923_),
    .ZN(_08924_));
 AOI211_X1 _34586_ (.A(_08876_),
    .B(_08924_),
    .C1(_08714_),
    .C2(_08658_),
    .ZN(_00631_));
 AOI211_X1 _34587_ (.A(\bp_fe_pc_gen_1.pc_if1_r [30]),
    .B(_08796_),
    .C1(_08797_),
    .C2(_08813_),
    .ZN(_08925_));
 NAND3_X2 _34588_ (.A1(_08785_),
    .A2(\bp_fe_pc_gen_1.btb.br_tgt_o [30]),
    .A3(_08771_),
    .ZN(_08926_));
 OAI21_X2 _34589_ (.A(fe_cmd_i[64]),
    .B1(_08773_),
    .B2(_08774_),
    .ZN(_08927_));
 OAI211_X4 _34590_ (.A(_08926_),
    .B(_08927_),
    .C1(_08613_),
    .C2(_08776_),
    .ZN(_08928_));
 NAND2_X1 _34591_ (.A1(_08921_),
    .A2(\bp_fe_pc_gen_1.pc_if1_r [29]),
    .ZN(_08929_));
 XNOR2_X2 _34592_ (.A(_08929_),
    .B(_00092_),
    .ZN(_08930_));
 NOR3_X4 _34593_ (.A1(_08778_),
    .A2(_08779_),
    .A3(_08930_),
    .ZN(_08931_));
 NOR2_X4 _34594_ (.A1(_08928_),
    .A2(_08931_),
    .ZN(_08932_));
 BUF_X8 _34595_ (.A(_08932_),
    .Z(_08933_));
 AOI211_X1 _34596_ (.A(_08876_),
    .B(_08925_),
    .C1(_08933_),
    .C2(_08665_),
    .ZN(_00633_));
 NAND3_X2 _34597_ (.A1(_08778_),
    .A2(net1405),
    .A3(_08771_),
    .ZN(_08934_));
 OAI21_X2 _34598_ (.A(fe_cmd_i[65]),
    .B1(_08476_),
    .B2(_08477_),
    .ZN(_08935_));
 OAI211_X4 _34599_ (.A(_08934_),
    .B(_08935_),
    .C1(_08616_),
    .C2(_08347_),
    .ZN(_08936_));
 AND3_X1 _34600_ (.A1(_08921_),
    .A2(\bp_fe_pc_gen_1.pc_if1_r [29]),
    .A3(\bp_fe_pc_gen_1.pc_if1_r [30]),
    .ZN(_08937_));
 XNOR2_X1 _34601_ (.A(_08937_),
    .B(\bp_fe_pc_gen_1.pc_if1_r [31]),
    .ZN(_08938_));
 NOR3_X2 _34602_ (.A1(_08786_),
    .A2(_08353_),
    .A3(_08938_),
    .ZN(_08939_));
 NOR3_X1 _34603_ (.A1(_08936_),
    .A2(_08790_),
    .A3(_08939_),
    .ZN(_08940_));
 AOI211_X1 _34604_ (.A(_08876_),
    .B(_08940_),
    .C1(_08717_),
    .C2(_08658_),
    .ZN(_00634_));
 AOI211_X1 _34605_ (.A(\bp_fe_pc_gen_1.pc_if1_r [32]),
    .B(_08796_),
    .C1(_08797_),
    .C2(_08813_),
    .ZN(_08941_));
 NAND3_X2 _34606_ (.A1(_08318_),
    .A2(net1404),
    .A3(_08339_),
    .ZN(_08942_));
 OAI21_X2 _34607_ (.A(fe_cmd_i[66]),
    .B1(_08331_),
    .B2(_08333_),
    .ZN(_08943_));
 OAI211_X4 _34608_ (.A(_08942_),
    .B(_08943_),
    .C1(_08619_),
    .C2(_08346_),
    .ZN(_08944_));
 NAND2_X1 _34609_ (.A1(_08937_),
    .A2(\bp_fe_pc_gen_1.pc_if1_r [31]),
    .ZN(_08945_));
 XNOR2_X2 _34610_ (.A(_08945_),
    .B(_00093_),
    .ZN(_08946_));
 NOR3_X2 _34611_ (.A1(_08785_),
    .A2(_08352_),
    .A3(_08946_),
    .ZN(_08947_));
 NOR2_X4 _34612_ (.A1(_08944_),
    .A2(_08947_),
    .ZN(_08948_));
 BUF_X8 _34613_ (.A(_08948_),
    .Z(_08949_));
 AOI211_X1 _34614_ (.A(_08876_),
    .B(_08941_),
    .C1(_08949_),
    .C2(_08665_),
    .ZN(_00635_));
 NAND3_X2 _34615_ (.A1(_08785_),
    .A2(net1403),
    .A3(_08339_),
    .ZN(_08950_));
 OAI21_X2 _34616_ (.A(fe_cmd_i[67]),
    .B1(_08331_),
    .B2(_08333_),
    .ZN(_08951_));
 OAI211_X4 _34617_ (.A(_08950_),
    .B(_08951_),
    .C1(_08622_),
    .C2(_08346_),
    .ZN(_08952_));
 AND3_X2 _34618_ (.A1(_08937_),
    .A2(\bp_fe_pc_gen_1.pc_if1_r [31]),
    .A3(\bp_fe_pc_gen_1.pc_if1_r [32]),
    .ZN(_08953_));
 XNOR2_X1 _34619_ (.A(_08953_),
    .B(\bp_fe_pc_gen_1.pc_if1_r [33]),
    .ZN(_08954_));
 NOR3_X2 _34620_ (.A1(_08319_),
    .A2(_08352_),
    .A3(_08954_),
    .ZN(_08955_));
 NOR3_X1 _34621_ (.A1(_08952_),
    .A2(_08672_),
    .A3(_08955_),
    .ZN(_08956_));
 AOI211_X1 _34622_ (.A(_08876_),
    .B(_08956_),
    .C1(_08720_),
    .C2(_08658_),
    .ZN(_00636_));
 BUF_X8 _34623_ (.A(_08650_),
    .Z(_08957_));
 AOI211_X2 _34624_ (.A(\bp_fe_pc_gen_1.pc_if1_r [34]),
    .B(_08655_),
    .C1(_08653_),
    .C2(_08813_),
    .ZN(_08958_));
 NAND3_X4 _34625_ (.A1(_08785_),
    .A2(\bp_fe_pc_gen_1.btb.br_tgt_o [34]),
    .A3(_08339_),
    .ZN(_08959_));
 OAI21_X2 _34626_ (.A(fe_cmd_i[68]),
    .B1(_08773_),
    .B2(_08774_),
    .ZN(_08960_));
 OAI211_X4 _34627_ (.A(_08959_),
    .B(_08960_),
    .C1(_08625_),
    .C2(_08776_),
    .ZN(_08961_));
 NAND2_X1 _34628_ (.A1(_08953_),
    .A2(\bp_fe_pc_gen_1.pc_if1_r [33]),
    .ZN(_08962_));
 XNOR2_X2 _34629_ (.A(_08962_),
    .B(_00094_),
    .ZN(_08963_));
 NOR3_X2 _34630_ (.A1(_08778_),
    .A2(_08779_),
    .A3(_08963_),
    .ZN(_08964_));
 NOR2_X4 _34631_ (.A1(_08961_),
    .A2(_08964_),
    .ZN(_08965_));
 BUF_X8 _34632_ (.A(_08965_),
    .Z(_08966_));
 AOI211_X1 _34633_ (.A(_08957_),
    .B(_08958_),
    .C1(_08966_),
    .C2(_08665_),
    .ZN(_00637_));
 NAND3_X2 _34634_ (.A1(_08786_),
    .A2(\bp_fe_pc_gen_1.btb.br_tgt_o [35]),
    .A3(_08340_),
    .ZN(_08967_));
 OAI21_X2 _34635_ (.A(fe_cmd_i[69]),
    .B1(_08476_),
    .B2(_08477_),
    .ZN(_08968_));
 OAI211_X4 _34636_ (.A(_08967_),
    .B(_08968_),
    .C1(_08628_),
    .C2(_08347_),
    .ZN(_08969_));
 AND3_X2 _34637_ (.A1(_08953_),
    .A2(\bp_fe_pc_gen_1.pc_if1_r [33]),
    .A3(\bp_fe_pc_gen_1.pc_if1_r [34]),
    .ZN(_08970_));
 XNOR2_X2 _34638_ (.A(_08970_),
    .B(\bp_fe_pc_gen_1.pc_if1_r [35]),
    .ZN(_08971_));
 NOR3_X2 _34639_ (.A1(_08320_),
    .A2(_08353_),
    .A3(_08971_),
    .ZN(_08972_));
 NOR3_X1 _34640_ (.A1(_08969_),
    .A2(_08672_),
    .A3(_08972_),
    .ZN(_08973_));
 AOI211_X1 _34641_ (.A(_08957_),
    .B(_08973_),
    .C1(_08725_),
    .C2(_08658_),
    .ZN(_00638_));
 AOI211_X1 _34642_ (.A(\bp_fe_pc_gen_1.pc_if1_r [36]),
    .B(_08655_),
    .C1(_08653_),
    .C2(_08337_),
    .ZN(_08974_));
 NAND3_X2 _34643_ (.A1(_08319_),
    .A2(\bp_fe_pc_gen_1.btb.br_tgt_o [36]),
    .A3(_08771_),
    .ZN(_08975_));
 OAI21_X2 _34644_ (.A(fe_cmd_i[70]),
    .B1(_08773_),
    .B2(_08774_),
    .ZN(_08976_));
 OAI211_X4 _34645_ (.A(_08975_),
    .B(_08976_),
    .C1(_08631_),
    .C2(_08776_),
    .ZN(_08977_));
 NAND2_X1 _34646_ (.A1(_08970_),
    .A2(\bp_fe_pc_gen_1.pc_if1_r [35]),
    .ZN(_08978_));
 XNOR2_X2 _34647_ (.A(_08978_),
    .B(_00095_),
    .ZN(_08979_));
 NOR3_X2 _34648_ (.A1(_08786_),
    .A2(_08779_),
    .A3(_08979_),
    .ZN(_08980_));
 NOR2_X4 _34649_ (.A1(_08977_),
    .A2(_08980_),
    .ZN(_08981_));
 BUF_X8 _34650_ (.A(_08981_),
    .Z(_08982_));
 AOI211_X1 _34651_ (.A(_08957_),
    .B(_08974_),
    .C1(_08982_),
    .C2(_08665_),
    .ZN(_00639_));
 NAND3_X2 _34652_ (.A1(_08785_),
    .A2(\bp_fe_pc_gen_1.btb.br_tgt_o [37]),
    .A3(_08339_),
    .ZN(_08983_));
 OAI21_X2 _34653_ (.A(fe_cmd_i[71]),
    .B1(_08331_),
    .B2(_08333_),
    .ZN(_08984_));
 OAI211_X4 _34654_ (.A(_08983_),
    .B(_08984_),
    .C1(_08634_),
    .C2(_08346_),
    .ZN(_08985_));
 NAND3_X2 _34655_ (.A1(_08970_),
    .A2(\bp_fe_pc_gen_1.pc_if1_r [35]),
    .A3(\bp_fe_pc_gen_1.pc_if1_r [36]),
    .ZN(_08986_));
 XNOR2_X2 _34656_ (.A(_08986_),
    .B(_08729_),
    .ZN(_08987_));
 NOR3_X2 _34657_ (.A1(_08319_),
    .A2(_08352_),
    .A3(_08987_),
    .ZN(_08988_));
 NOR3_X1 _34658_ (.A1(_08985_),
    .A2(_08672_),
    .A3(_08988_),
    .ZN(_08989_));
 AOI211_X1 _34659_ (.A(_08957_),
    .B(_08989_),
    .C1(_08729_),
    .C2(_08658_),
    .ZN(_00640_));
 AOI211_X1 _34660_ (.A(\bp_fe_pc_gen_1.pc_if1_r [38]),
    .B(_08655_),
    .C1(_08653_),
    .C2(_08337_),
    .ZN(_08990_));
 NAND3_X2 _34661_ (.A1(_08319_),
    .A2(net1402),
    .A3(_08771_),
    .ZN(_08991_));
 OAI21_X2 _34662_ (.A(fe_cmd_i[72]),
    .B1(_08773_),
    .B2(_08774_),
    .ZN(_08992_));
 OAI211_X4 _34663_ (.A(_08991_),
    .B(_08992_),
    .C1(_08637_),
    .C2(_08776_),
    .ZN(_08993_));
 NOR2_X1 _34664_ (.A1(_08986_),
    .A2(_08729_),
    .ZN(_08994_));
 XNOR2_X2 _34665_ (.A(_08994_),
    .B(\bp_fe_pc_gen_1.pc_if1_r [38]),
    .ZN(_08995_));
 NOR3_X2 _34666_ (.A1(_08786_),
    .A2(_08779_),
    .A3(_08995_),
    .ZN(_08996_));
 NOR2_X4 _34667_ (.A1(_08993_),
    .A2(_08996_),
    .ZN(_08997_));
 AOI211_X1 _34668_ (.A(_08957_),
    .B(_08990_),
    .C1(_08997_),
    .C2(_08665_),
    .ZN(_00641_));
 BUF_X8 _34669_ (.A(_08516_),
    .Z(_08998_));
 BUF_X8 _34670_ (.A(_08998_),
    .Z(_08999_));
 NOR2_X1 _34671_ (.A1(_08661_),
    .A2(_08999_),
    .ZN(_00729_));
 BUF_X8 _34672_ (.A(_08998_),
    .Z(_09000_));
 NAND2_X2 _34673_ (.A1(_08652_),
    .A2(_08523_),
    .ZN(_09001_));
 NOR3_X1 _34674_ (.A1(_08037_),
    .A2(\bp_fe_pc_gen_1.state_r [0]),
    .A3(_08335_),
    .ZN(_09002_));
 AOI21_X1 _34675_ (.A(_09002_),
    .B1(_08033_),
    .B2(_08525_),
    .ZN(_09003_));
 AOI21_X1 _34676_ (.A(_09000_),
    .B1(_09001_),
    .B2(_09003_),
    .ZN(_00730_));
 NOR2_X1 _34677_ (.A1(_08514_),
    .A2(_08999_),
    .ZN(_00609_));
 AND2_X1 _34678_ (.A1(_08038_),
    .A2(_08723_),
    .ZN(_00727_));
 OAI211_X1 _34679_ (.A(_08674_),
    .B(\bp_fe_pc_gen_1.pc_v_if1_r ),
    .C1(_08649_),
    .C2(_00080_),
    .ZN(_09004_));
 NOR3_X1 _34680_ (.A1(_08645_),
    .A2(\bp_fe_pc_gen_1.itlb_miss_if2_r ),
    .A3(_09004_),
    .ZN(_00728_));
 INV_X1 _34681_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [0]),
    .ZN(_09005_));
 BUF_X8 _34682_ (.A(_08641_),
    .Z(_09006_));
 BUF_X8 _34683_ (.A(_09006_),
    .Z(_09007_));
 BUF_X8 _34684_ (.A(\bp_fe_pc_gen_1.pc_v_if2_r ),
    .Z(_09008_));
 BUF_X8 _34685_ (.A(_09008_),
    .Z(_09009_));
 AOI21_X4 _34686_ (.A(_09005_),
    .B1(_09007_),
    .B2(_09009_),
    .ZN(fe_queue_o[1]));
 INV_X1 _34687_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [1]),
    .ZN(_09010_));
 AOI21_X4 _34688_ (.A(_09010_),
    .B1(_09007_),
    .B2(_09009_),
    .ZN(fe_queue_o[2]));
 INV_X1 _34689_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [2]),
    .ZN(_09011_));
 AOI21_X4 _34690_ (.A(_09011_),
    .B1(_09007_),
    .B2(_09009_),
    .ZN(fe_queue_o[3]));
 INV_X1 _34691_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [3]),
    .ZN(_09012_));
 AOI21_X4 _34692_ (.A(_09012_),
    .B1(_09007_),
    .B2(_09009_),
    .ZN(fe_queue_o[4]));
 INV_X1 _34693_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [4]),
    .ZN(_09013_));
 AOI21_X4 _34694_ (.A(_09013_),
    .B1(_09007_),
    .B2(_09009_),
    .ZN(fe_queue_o[5]));
 INV_X1 _34695_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [5]),
    .ZN(_09014_));
 AOI21_X4 _34696_ (.A(_09014_),
    .B1(_09007_),
    .B2(_09009_),
    .ZN(fe_queue_o[6]));
 INV_X1 _34697_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [6]),
    .ZN(_09015_));
 AOI21_X4 _34698_ (.A(_09015_),
    .B1(_09007_),
    .B2(_09009_),
    .ZN(fe_queue_o[7]));
 INV_X1 _34699_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [7]),
    .ZN(_09016_));
 AOI21_X4 _34700_ (.A(_09016_),
    .B1(_09007_),
    .B2(_09009_),
    .ZN(fe_queue_o[8]));
 INV_X1 _34701_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [8]),
    .ZN(_09017_));
 AOI21_X4 _34702_ (.A(_09017_),
    .B1(_09007_),
    .B2(_09009_),
    .ZN(fe_queue_o[9]));
 INV_X1 _34703_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [9]),
    .ZN(_09018_));
 AOI21_X4 _34704_ (.A(_09018_),
    .B1(_09007_),
    .B2(_09009_),
    .ZN(fe_queue_o[10]));
 INV_X2 _34705_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [10]),
    .ZN(_09019_));
 BUF_X8 _34706_ (.A(_09006_),
    .Z(_09020_));
 BUF_X8 _34707_ (.A(_09008_),
    .Z(_09021_));
 AOI21_X4 _34708_ (.A(_09019_),
    .B1(_09020_),
    .B2(_09021_),
    .ZN(fe_queue_o[11]));
 INV_X1 _34709_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [11]),
    .ZN(_09022_));
 AOI21_X4 _34710_ (.A(_09022_),
    .B1(_09020_),
    .B2(_09021_),
    .ZN(fe_queue_o[12]));
 INV_X1 _34711_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [12]),
    .ZN(_09023_));
 AOI21_X4 _34712_ (.A(_09023_),
    .B1(_09020_),
    .B2(_09021_),
    .ZN(fe_queue_o[13]));
 INV_X1 _34713_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [13]),
    .ZN(_09024_));
 AOI21_X4 _34714_ (.A(_09024_),
    .B1(_09020_),
    .B2(_09021_),
    .ZN(fe_queue_o[14]));
 INV_X1 _34715_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [14]),
    .ZN(_09025_));
 AOI21_X4 _34716_ (.A(_09025_),
    .B1(_09020_),
    .B2(_09021_),
    .ZN(fe_queue_o[15]));
 INV_X1 _34717_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [15]),
    .ZN(_09026_));
 AOI21_X4 _34718_ (.A(_09026_),
    .B1(_09020_),
    .B2(_09021_),
    .ZN(fe_queue_o[16]));
 INV_X1 _34719_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [16]),
    .ZN(_09027_));
 AOI21_X4 _34720_ (.A(_09027_),
    .B1(_09020_),
    .B2(_09021_),
    .ZN(fe_queue_o[17]));
 INV_X1 _34721_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [17]),
    .ZN(_09028_));
 AOI21_X4 _34722_ (.A(_09028_),
    .B1(_09020_),
    .B2(_09021_),
    .ZN(fe_queue_o[18]));
 INV_X1 _34723_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [18]),
    .ZN(_09029_));
 AOI21_X4 _34724_ (.A(_09029_),
    .B1(_09020_),
    .B2(_09021_),
    .ZN(fe_queue_o[19]));
 INV_X1 _34725_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [19]),
    .ZN(_09030_));
 AOI21_X4 _34726_ (.A(_09030_),
    .B1(_09020_),
    .B2(_09021_),
    .ZN(fe_queue_o[20]));
 INV_X1 _34727_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [20]),
    .ZN(_09031_));
 AOI21_X4 _34728_ (.A(_09031_),
    .B1(_09006_),
    .B2(_09008_),
    .ZN(fe_queue_o[21]));
 INV_X1 _34729_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [21]),
    .ZN(_09032_));
 AOI21_X4 _34730_ (.A(_09032_),
    .B1(_09006_),
    .B2(_09008_),
    .ZN(fe_queue_o[22]));
 INV_X1 _34731_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [22]),
    .ZN(_09033_));
 AOI21_X4 _34732_ (.A(_09033_),
    .B1(_09006_),
    .B2(_09008_),
    .ZN(fe_queue_o[23]));
 INV_X1 _34733_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [23]),
    .ZN(_09034_));
 AOI21_X4 _34734_ (.A(_09034_),
    .B1(_09006_),
    .B2(_09008_),
    .ZN(fe_queue_o[24]));
 INV_X1 _34735_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [24]),
    .ZN(_09035_));
 AOI21_X4 _34736_ (.A(_09035_),
    .B1(_09006_),
    .B2(_09008_),
    .ZN(fe_queue_o[25]));
 INV_X1 _34737_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [25]),
    .ZN(_09036_));
 AOI21_X4 _34738_ (.A(_09036_),
    .B1(_09006_),
    .B2(_09008_),
    .ZN(fe_queue_o[26]));
 INV_X1 _34739_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [26]),
    .ZN(_09037_));
 AOI21_X4 _34740_ (.A(_09037_),
    .B1(_09006_),
    .B2(_09008_),
    .ZN(fe_queue_o[27]));
 INV_X2 _34741_ (.A(net1389),
    .ZN(_09038_));
 BUF_X8 _34742_ (.A(_09038_),
    .Z(_09039_));
 INV_X4 _34743_ (.A(net1264),
    .ZN(_09040_));
 BUF_X8 _34744_ (.A(_09040_),
    .Z(_09041_));
 BUF_X8 _34745_ (.A(_09041_),
    .Z(_09042_));
 XNOR2_X2 _34746_ (.A(_07583_),
    .B(\icache.addr_tv_r [4]),
    .ZN(_09043_));
 INV_X2 _34747_ (.A(_09043_),
    .ZN(_09044_));
 BUF_X8 _34748_ (.A(_09044_),
    .Z(_09045_));
 NOR2_X4 _34749_ (.A1(_07592_),
    .A2(_07600_),
    .ZN(_09046_));
 XNOR2_X2 _34750_ (.A(_09046_),
    .B(\icache.addr_tv_r [3]),
    .ZN(_09047_));
 BUF_X8 _34751_ (.A(_09047_),
    .Z(_09048_));
 NOR2_X4 _34752_ (.A1(_09045_),
    .A2(_09048_),
    .ZN(_09049_));
 AND2_X4 _34753_ (.A1(_07573_),
    .A2(_07578_),
    .ZN(_09050_));
 INV_X1 _34754_ (.A(\icache.addr_tv_r [5]),
    .ZN(_09051_));
 XNOR2_X2 _34755_ (.A(_09050_),
    .B(_09051_),
    .ZN(_09052_));
 BUF_X4 _34756_ (.A(_09052_),
    .Z(_09053_));
 BUF_X8 _34757_ (.A(_09053_),
    .Z(_09054_));
 AND2_X1 _34758_ (.A1(_09049_),
    .A2(_09054_),
    .ZN(_09055_));
 BUF_X8 _34759_ (.A(_09055_),
    .Z(_09056_));
 INV_X4 _34760_ (.A(_09056_),
    .ZN(_09057_));
 BUF_X4 _34761_ (.A(_09057_),
    .Z(_09058_));
 AND2_X4 _34762_ (.A1(_09047_),
    .A2(_09043_),
    .ZN(_09059_));
 AND2_X4 _34763_ (.A1(_09059_),
    .A2(_09053_),
    .ZN(_09060_));
 INV_X8 _34764_ (.A(_09060_),
    .ZN(_09061_));
 BUF_X8 _34765_ (.A(_09061_),
    .Z(_09062_));
 AND2_X2 _34766_ (.A1(_09044_),
    .A2(_09047_),
    .ZN(_09063_));
 BUF_X8 _34767_ (.A(_09063_),
    .Z(_09064_));
 BUF_X8 _34768_ (.A(_09064_),
    .Z(_09065_));
 BUF_X8 _34769_ (.A(_09065_),
    .Z(_09066_));
 INV_X2 _34770_ (.A(_09052_),
    .ZN(_09067_));
 BUF_X4 _34771_ (.A(_09067_),
    .Z(_09068_));
 BUF_X8 _34772_ (.A(_09068_),
    .Z(_09069_));
 BUF_X8 _34773_ (.A(_09069_),
    .Z(_09070_));
 NAND3_X2 _34774_ (.A1(_09066_),
    .A2(\icache.data_set_select_mux.data_i [480]),
    .A3(_09070_),
    .ZN(_09071_));
 NOR2_X4 _34775_ (.A1(_09047_),
    .A2(_09043_),
    .ZN(_09072_));
 AND2_X2 _34776_ (.A1(_09072_),
    .A2(_09067_),
    .ZN(_09073_));
 INV_X2 _34777_ (.A(_09073_),
    .ZN(_09074_));
 BUF_X8 _34778_ (.A(_09074_),
    .Z(_09075_));
 BUF_X8 _34779_ (.A(_09075_),
    .Z(_09076_));
 BUF_X16 _34780_ (.A(_09076_),
    .Z(_09077_));
 OAI21_X4 _34781_ (.A(_09071_),
    .B1(_09077_),
    .B2(_00111_),
    .ZN(_09078_));
 BUF_X8 _34782_ (.A(_09045_),
    .Z(_09079_));
 BUF_X8 _34783_ (.A(_09079_),
    .Z(_09080_));
 BUF_X8 _34784_ (.A(_09080_),
    .Z(_09081_));
 INV_X1 _34785_ (.A(_09047_),
    .ZN(_09082_));
 BUF_X4 _34786_ (.A(_09082_),
    .Z(_09083_));
 BUF_X8 _34787_ (.A(_09083_),
    .Z(_09084_));
 BUF_X8 _34788_ (.A(_09084_),
    .Z(_09085_));
 BUF_X8 _34789_ (.A(_09085_),
    .Z(_09086_));
 BUF_X8 _34790_ (.A(_09054_),
    .Z(_09087_));
 BUF_X8 _34791_ (.A(_09087_),
    .Z(_09088_));
 NOR4_X4 _34792_ (.A1(_09081_),
    .A2(_09086_),
    .A3(_09088_),
    .A4(_00110_),
    .ZN(_09089_));
 BUF_X4 _34793_ (.A(_09054_),
    .Z(_09090_));
 BUF_X8 _34794_ (.A(_09090_),
    .Z(_09091_));
 BUF_X4 _34795_ (.A(_09048_),
    .Z(_09092_));
 BUF_X8 _34796_ (.A(_09092_),
    .Z(_09093_));
 NOR4_X1 _34797_ (.A1(_09081_),
    .A2(_09091_),
    .A3(_09093_),
    .A4(_00109_),
    .ZN(_09094_));
 NOR3_X2 _34798_ (.A1(_09078_),
    .A2(_09089_),
    .A3(_09094_),
    .ZN(_09095_));
 BUF_X4 _34799_ (.A(_09069_),
    .Z(_09096_));
 BUF_X8 _34800_ (.A(_09084_),
    .Z(_09097_));
 BUF_X8 _34801_ (.A(_09097_),
    .Z(_09098_));
 BUF_X4 _34802_ (.A(_09043_),
    .Z(_09099_));
 BUF_X4 _34803_ (.A(_09099_),
    .Z(_09100_));
 BUF_X4 _34804_ (.A(_09100_),
    .Z(_09101_));
 OR4_X1 _34805_ (.A1(_00108_),
    .A2(_09096_),
    .A3(_09098_),
    .A4(_09101_),
    .ZN(_09102_));
 AND2_X4 _34806_ (.A1(_09072_),
    .A2(_09052_),
    .ZN(_09103_));
 INV_X2 _34807_ (.A(_09103_),
    .ZN(_09104_));
 BUF_X8 _34808_ (.A(_09104_),
    .Z(_09105_));
 BUF_X4 _34809_ (.A(_09105_),
    .Z(_09106_));
 OR2_X1 _34810_ (.A1(_09106_),
    .A2(_00107_),
    .ZN(_09107_));
 AND4_X4 _34811_ (.A1(_09062_),
    .A2(_09095_),
    .A3(_09102_),
    .A4(_09107_),
    .ZN(_09108_));
 BUF_X8 _34812_ (.A(_09054_),
    .Z(_09109_));
 BUF_X8 _34813_ (.A(_09109_),
    .Z(_09110_));
 BUF_X4 _34814_ (.A(_09110_),
    .Z(_09111_));
 BUF_X8 _34815_ (.A(_09048_),
    .Z(_09112_));
 BUF_X4 _34816_ (.A(_09112_),
    .Z(_09113_));
 BUF_X4 _34817_ (.A(_09113_),
    .Z(_09114_));
 BUF_X4 _34818_ (.A(_09101_),
    .Z(_09115_));
 AND4_X1 _34819_ (.A1(_00106_),
    .A2(_09111_),
    .A3(_09114_),
    .A4(_09115_),
    .ZN(_09116_));
 OAI221_X2 _34820_ (.A(_09042_),
    .B1(_00105_),
    .B2(_09058_),
    .C1(_09108_),
    .C2(_09116_),
    .ZN(_09117_));
 BUF_X8 _34821_ (.A(net1263),
    .Z(_09118_));
 NAND2_X1 _34822_ (.A1(_09118_),
    .A2(_00104_),
    .ZN(_09119_));
 AOI21_X2 _34823_ (.A(_09039_),
    .B1(_09117_),
    .B2(_09119_),
    .ZN(_09120_));
 BUF_X4 _34824_ (.A(net1390),
    .Z(_09121_));
 BUF_X8 _34825_ (.A(_09070_),
    .Z(_09122_));
 BUF_X8 _34826_ (.A(_09079_),
    .Z(_09123_));
 BUF_X8 _34827_ (.A(_09123_),
    .Z(_09124_));
 BUF_X4 _34828_ (.A(_09124_),
    .Z(_09125_));
 BUF_X4 _34829_ (.A(_09093_),
    .Z(_09126_));
 OR4_X2 _34830_ (.A1(_00097_),
    .A2(_09122_),
    .A3(_09125_),
    .A4(_09126_),
    .ZN(_09127_));
 BUF_X4 _34831_ (.A(_09064_),
    .Z(_09128_));
 BUF_X8 _34832_ (.A(_09128_),
    .Z(_09129_));
 BUF_X8 _34833_ (.A(_09068_),
    .Z(_09130_));
 BUF_X8 _34834_ (.A(_09130_),
    .Z(_09131_));
 NAND3_X1 _34835_ (.A1(_09129_),
    .A2(\icache.data_set_select_mux.data_i [448]),
    .A3(_09131_),
    .ZN(_09132_));
 BUF_X8 _34836_ (.A(_09076_),
    .Z(_09133_));
 OAI21_X1 _34837_ (.A(_09132_),
    .B1(_09133_),
    .B2(_00103_),
    .ZN(_09134_));
 BUF_X8 _34838_ (.A(_09085_),
    .Z(_09135_));
 BUF_X8 _34839_ (.A(_09079_),
    .Z(_09136_));
 BUF_X8 _34840_ (.A(_09136_),
    .Z(_09137_));
 BUF_X8 _34841_ (.A(_09090_),
    .Z(_09138_));
 NOR4_X1 _34842_ (.A1(_09135_),
    .A2(_09137_),
    .A3(_09138_),
    .A4(_00102_),
    .ZN(_09139_));
 BUF_X8 _34843_ (.A(_09087_),
    .Z(_09140_));
 BUF_X8 _34844_ (.A(_09112_),
    .Z(_09141_));
 NOR4_X2 _34845_ (.A1(_09137_),
    .A2(_09140_),
    .A3(_09141_),
    .A4(_00101_),
    .ZN(_09142_));
 OR3_X4 _34846_ (.A1(_09134_),
    .A2(_09139_),
    .A3(_09142_),
    .ZN(_09143_));
 BUF_X4 _34847_ (.A(_09068_),
    .Z(_09144_));
 BUF_X8 _34848_ (.A(_09144_),
    .Z(_09145_));
 BUF_X8 _34849_ (.A(_09145_),
    .Z(_09146_));
 BUF_X8 _34850_ (.A(_09146_),
    .Z(_09147_));
 BUF_X8 _34851_ (.A(_09135_),
    .Z(_09148_));
 BUF_X4 _34852_ (.A(_09100_),
    .Z(_09149_));
 BUF_X4 _34853_ (.A(_09149_),
    .Z(_09150_));
 NOR4_X2 _34854_ (.A1(_09147_),
    .A2(_09148_),
    .A3(_00100_),
    .A4(_09150_),
    .ZN(_09151_));
 BUF_X8 _34855_ (.A(_09105_),
    .Z(_09152_));
 BUF_X8 _34856_ (.A(_09152_),
    .Z(_09153_));
 OAI21_X2 _34857_ (.A(_09062_),
    .B1(_09153_),
    .B2(_00099_),
    .ZN(_09154_));
 NOR3_X4 _34858_ (.A1(_09143_),
    .A2(_09151_),
    .A3(_09154_),
    .ZN(_09155_));
 BUF_X4 _34859_ (.A(_09059_),
    .Z(_09156_));
 AND3_X1 _34860_ (.A1(_09156_),
    .A2(_00098_),
    .A3(_09111_),
    .ZN(_09157_));
 OAI211_X4 _34861_ (.A(_09042_),
    .B(_09127_),
    .C1(_09155_),
    .C2(_09157_),
    .ZN(_09158_));
 NAND2_X1 _34862_ (.A1(_09118_),
    .A2(_00096_),
    .ZN(_09159_));
 AOI21_X2 _34863_ (.A(_09121_),
    .B1(_09158_),
    .B2(_09159_),
    .ZN(_09160_));
 NOR3_X4 _34864_ (.A1(_09120_),
    .A2(_09160_),
    .A3(fe_queue_o[99]),
    .ZN(fe_queue_o[28]));
 AND2_X4 _34865_ (.A1(_09049_),
    .A2(_09069_),
    .ZN(_09161_));
 INV_X1 _34866_ (.A(_09161_),
    .ZN(_09162_));
 NOR2_X1 _34867_ (.A1(_09162_),
    .A2(_00125_),
    .ZN(_09163_));
 NAND3_X1 _34868_ (.A1(_09129_),
    .A2(\icache.data_set_select_mux.data_i [481]),
    .A3(_09131_),
    .ZN(_09164_));
 OAI21_X4 _34869_ (.A(_09164_),
    .B1(_09133_),
    .B2(_00127_),
    .ZN(_09165_));
 BUF_X4 _34870_ (.A(_09087_),
    .Z(_09166_));
 NOR4_X2 _34871_ (.A1(_09081_),
    .A2(_09086_),
    .A3(_09166_),
    .A4(_00126_),
    .ZN(_09167_));
 NOR3_X4 _34872_ (.A1(_09163_),
    .A2(_09165_),
    .A3(_09167_),
    .ZN(_09168_));
 OR4_X1 _34873_ (.A1(_00124_),
    .A2(_09096_),
    .A3(_09098_),
    .A4(_09101_),
    .ZN(_09169_));
 OR4_X1 _34874_ (.A1(_00123_),
    .A2(_09096_),
    .A3(_09101_),
    .A4(_09093_),
    .ZN(_09170_));
 AND4_X4 _34875_ (.A1(_09062_),
    .A2(_09168_),
    .A3(_09169_),
    .A4(_09170_),
    .ZN(_09171_));
 BUF_X8 _34876_ (.A(_09110_),
    .Z(_09172_));
 AND4_X1 _34877_ (.A1(_00122_),
    .A2(_09172_),
    .A3(_09114_),
    .A4(_09115_),
    .ZN(_09173_));
 OAI221_X2 _34878_ (.A(_09042_),
    .B1(_00121_),
    .B2(_09058_),
    .C1(_09171_),
    .C2(_09173_),
    .ZN(_09174_));
 NAND2_X1 _34879_ (.A1(_09118_),
    .A2(_00120_),
    .ZN(_09175_));
 AOI21_X2 _34880_ (.A(_09039_),
    .B1(_09174_),
    .B2(_09175_),
    .ZN(_09176_));
 BUF_X8 _34881_ (.A(_09040_),
    .Z(_09177_));
 BUF_X8 _34882_ (.A(_09177_),
    .Z(_09178_));
 NAND3_X2 _34883_ (.A1(_09066_),
    .A2(\icache.data_set_select_mux.data_i [449]),
    .A3(_09070_),
    .ZN(_09179_));
 OAI21_X2 _34884_ (.A(_09179_),
    .B1(_09077_),
    .B2(_00119_),
    .ZN(_09180_));
 NOR4_X2 _34885_ (.A1(_09135_),
    .A2(_09137_),
    .A3(_09091_),
    .A4(_00118_),
    .ZN(_09181_));
 NOR4_X2 _34886_ (.A1(_09081_),
    .A2(_09091_),
    .A3(_09093_),
    .A4(_00117_),
    .ZN(_09182_));
 NOR3_X4 _34887_ (.A1(_09180_),
    .A2(_09181_),
    .A3(_09182_),
    .ZN(_09183_));
 OR4_X1 _34888_ (.A1(_00116_),
    .A2(_09096_),
    .A3(_09098_),
    .A4(_09101_),
    .ZN(_09184_));
 BUF_X4 _34889_ (.A(_09144_),
    .Z(_09185_));
 BUF_X4 _34890_ (.A(_09099_),
    .Z(_09186_));
 OR4_X1 _34891_ (.A1(_00115_),
    .A2(_09185_),
    .A3(_09186_),
    .A4(_09112_),
    .ZN(_09187_));
 AND2_X1 _34892_ (.A1(_09187_),
    .A2(_09062_),
    .ZN(_09188_));
 AND3_X2 _34893_ (.A1(_09183_),
    .A2(_09184_),
    .A3(_09188_),
    .ZN(_09189_));
 AND3_X1 _34894_ (.A1(_09156_),
    .A2(_00114_),
    .A3(_09172_),
    .ZN(_09190_));
 OAI221_X2 _34895_ (.A(_09178_),
    .B1(_00113_),
    .B2(_09058_),
    .C1(_09189_),
    .C2(_09190_),
    .ZN(_09191_));
 NAND2_X2 _34896_ (.A1(_09118_),
    .A2(_00112_),
    .ZN(_09192_));
 AOI21_X2 _34897_ (.A(_09121_),
    .B1(_09191_),
    .B2(_09192_),
    .ZN(_09193_));
 NOR3_X4 _34898_ (.A1(_09176_),
    .A2(fe_queue_o[99]),
    .A3(_09193_),
    .ZN(fe_queue_o[29]));
 BUF_X8 _34899_ (.A(_09177_),
    .Z(_09194_));
 BUF_X8 _34900_ (.A(_09075_),
    .Z(_09195_));
 NOR2_X2 _34901_ (.A1(_09195_),
    .A2(_00135_),
    .ZN(_09196_));
 BUF_X4 _34902_ (.A(_09064_),
    .Z(_09197_));
 BUF_X8 _34903_ (.A(_09144_),
    .Z(_09198_));
 AND3_X1 _34904_ (.A1(_09197_),
    .A2(\icache.data_set_select_mux.data_i [450]),
    .A3(_09198_),
    .ZN(_09199_));
 BUF_X4 _34905_ (.A(_09083_),
    .Z(_09200_));
 BUF_X8 _34906_ (.A(_09200_),
    .Z(_09201_));
 BUF_X4 _34907_ (.A(_09053_),
    .Z(_09202_));
 BUF_X4 _34908_ (.A(_09202_),
    .Z(_09203_));
 NOR4_X4 _34909_ (.A1(_09124_),
    .A2(_09201_),
    .A3(_09203_),
    .A4(_00134_),
    .ZN(_09204_));
 NOR3_X4 _34910_ (.A1(_09196_),
    .A2(_09199_),
    .A3(_09204_),
    .ZN(_09205_));
 BUF_X4 _34911_ (.A(_09045_),
    .Z(_09206_));
 BUF_X8 _34912_ (.A(_09206_),
    .Z(_09207_));
 BUF_X4 _34913_ (.A(_09048_),
    .Z(_09208_));
 OR4_X4 _34914_ (.A1(_00133_),
    .A2(_09207_),
    .A3(_09203_),
    .A4(_09208_),
    .ZN(_09209_));
 BUF_X4 _34915_ (.A(_09084_),
    .Z(_09210_));
 BUF_X4 _34916_ (.A(_09099_),
    .Z(_09211_));
 OR4_X1 _34917_ (.A1(_00132_),
    .A2(_09198_),
    .A3(_09210_),
    .A4(_09211_),
    .ZN(_09212_));
 NOR2_X1 _34918_ (.A1(_09152_),
    .A2(_00131_),
    .ZN(_09213_));
 BUF_X8 _34919_ (.A(_09060_),
    .Z(_09214_));
 NOR2_X4 _34920_ (.A1(_09213_),
    .A2(_09214_),
    .ZN(_09215_));
 AND4_X2 _34921_ (.A1(_09205_),
    .A2(_09209_),
    .A3(_09212_),
    .A4(_09215_),
    .ZN(_09216_));
 BUF_X8 _34922_ (.A(_09110_),
    .Z(_09217_));
 AND4_X1 _34923_ (.A1(_00130_),
    .A2(_09217_),
    .A3(_09114_),
    .A4(_09115_),
    .ZN(_09218_));
 OAI221_X2 _34924_ (.A(_09194_),
    .B1(_00129_),
    .B2(_09058_),
    .C1(_09216_),
    .C2(_09218_),
    .ZN(_09219_));
 BUF_X4 _34925_ (.A(net1264),
    .Z(_09220_));
 NAND2_X1 _34926_ (.A1(_09220_),
    .A2(_00128_),
    .ZN(_09221_));
 AOI21_X1 _34927_ (.A(_09121_),
    .B1(_09219_),
    .B2(_09221_),
    .ZN(_09222_));
 BUF_X4 _34928_ (.A(_09121_),
    .Z(_09223_));
 NAND3_X1 _34929_ (.A1(_09066_),
    .A2(\icache.data_set_select_mux.data_i [482]),
    .A3(_09096_),
    .ZN(_09224_));
 OAI21_X1 _34930_ (.A(_09224_),
    .B1(_09077_),
    .B2(_00143_),
    .ZN(_09225_));
 NOR4_X4 _34931_ (.A1(_09081_),
    .A2(_09086_),
    .A3(_09166_),
    .A4(_00142_),
    .ZN(_09226_));
 BUF_X8 _34932_ (.A(_09080_),
    .Z(_09227_));
 NOR4_X4 _34933_ (.A1(_09227_),
    .A2(_09091_),
    .A3(_09093_),
    .A4(_00141_),
    .ZN(_09228_));
 NOR3_X2 _34934_ (.A1(_09225_),
    .A2(_09226_),
    .A3(_09228_),
    .ZN(_09229_));
 BUF_X8 _34935_ (.A(_09069_),
    .Z(_09230_));
 BUF_X8 _34936_ (.A(_09083_),
    .Z(_09231_));
 BUF_X4 _34937_ (.A(_09231_),
    .Z(_09232_));
 OR4_X2 _34938_ (.A1(_00140_),
    .A2(_09230_),
    .A3(_09232_),
    .A4(_09101_),
    .ZN(_09233_));
 OR2_X4 _34939_ (.A1(_09106_),
    .A2(_00139_),
    .ZN(_09234_));
 NAND3_X4 _34940_ (.A1(_09229_),
    .A2(_09233_),
    .A3(_09234_),
    .ZN(_09235_));
 NOR4_X2 _34941_ (.A1(_09147_),
    .A2(_09148_),
    .A3(_00138_),
    .A4(_09125_),
    .ZN(_09236_));
 BUF_X4 _34942_ (.A(_09146_),
    .Z(_09237_));
 BUF_X8 _34943_ (.A(_09079_),
    .Z(_09238_));
 BUF_X8 _34944_ (.A(_09238_),
    .Z(_09239_));
 BUF_X4 _34945_ (.A(_09239_),
    .Z(_09240_));
 BUF_X4 _34946_ (.A(_09113_),
    .Z(_09241_));
 NOR4_X2 _34947_ (.A1(_09237_),
    .A2(_09240_),
    .A3(_09241_),
    .A4(_00137_),
    .ZN(_09242_));
 NOR3_X4 _34948_ (.A1(_09235_),
    .A2(_09236_),
    .A3(_09242_),
    .ZN(_09243_));
 MUX2_X1 _34949_ (.A(_00136_),
    .B(_09243_),
    .S(_09178_),
    .Z(_09244_));
 AOI211_X2 _34950_ (.A(fe_queue_o[99]),
    .B(_09222_),
    .C1(_09223_),
    .C2(_09244_),
    .ZN(fe_queue_o[30]));
 BUF_X8 _34951_ (.A(_09040_),
    .Z(_09245_));
 NOR2_X1 _34952_ (.A1(_09195_),
    .A2(_00151_),
    .ZN(_09246_));
 AND3_X1 _34953_ (.A1(_09065_),
    .A2(\icache.data_set_select_mux.data_i [451]),
    .A3(_09069_),
    .ZN(_09247_));
 NOR4_X1 _34954_ (.A1(_09080_),
    .A2(_09085_),
    .A3(_09090_),
    .A4(_00150_),
    .ZN(_09248_));
 NOR3_X1 _34955_ (.A1(_09246_),
    .A2(_09247_),
    .A3(_09248_),
    .ZN(_09249_));
 OR4_X1 _34956_ (.A1(_00149_),
    .A2(_09136_),
    .A3(_09087_),
    .A4(_09092_),
    .ZN(_09250_));
 OR4_X2 _34957_ (.A1(_00148_),
    .A2(_09185_),
    .A3(_09097_),
    .A4(_09186_),
    .ZN(_09251_));
 AND3_X2 _34958_ (.A1(_09249_),
    .A2(_09250_),
    .A3(_09251_),
    .ZN(_09252_));
 OR2_X1 _34959_ (.A1(_09153_),
    .A2(_00147_),
    .ZN(_09253_));
 BUF_X4 _34960_ (.A(_09045_),
    .Z(_09254_));
 BUF_X4 _34961_ (.A(_09254_),
    .Z(_09255_));
 OR4_X1 _34962_ (.A1(_00146_),
    .A2(_09096_),
    .A3(_09232_),
    .A4(_09255_),
    .ZN(_09256_));
 NAND3_X1 _34963_ (.A1(_09252_),
    .A2(_09253_),
    .A3(_09256_),
    .ZN(_09257_));
 BUF_X8 _34964_ (.A(_09080_),
    .Z(_09258_));
 BUF_X8 _34965_ (.A(_09258_),
    .Z(_09259_));
 NOR4_X1 _34966_ (.A1(_09147_),
    .A2(_09259_),
    .A3(_09126_),
    .A4(_00145_),
    .ZN(_09260_));
 OAI21_X1 _34967_ (.A(_09245_),
    .B1(_09257_),
    .B2(_09260_),
    .ZN(_09261_));
 BUF_X4 _34968_ (.A(_09038_),
    .Z(_09262_));
 OR2_X1 _34969_ (.A1(_09041_),
    .A2(_00144_),
    .ZN(_09263_));
 AND3_X1 _34970_ (.A1(_09261_),
    .A2(_09262_),
    .A3(_09263_),
    .ZN(_09264_));
 NAND3_X2 _34971_ (.A1(_09066_),
    .A2(\icache.data_set_select_mux.data_i [483]),
    .A3(_09230_),
    .ZN(_09265_));
 OAI21_X4 _34972_ (.A(_09265_),
    .B1(_09077_),
    .B2(_00159_),
    .ZN(_09266_));
 BUF_X8 _34973_ (.A(_09085_),
    .Z(_09267_));
 NOR4_X2 _34974_ (.A1(_09239_),
    .A2(_09267_),
    .A3(_09166_),
    .A4(_00158_),
    .ZN(_09268_));
 NOR4_X2 _34975_ (.A1(_09227_),
    .A2(_09088_),
    .A3(_09093_),
    .A4(_00157_),
    .ZN(_09269_));
 NOR3_X4 _34976_ (.A1(_09266_),
    .A2(_09268_),
    .A3(_09269_),
    .ZN(_09270_));
 BUF_X4 _34977_ (.A(_09069_),
    .Z(_09271_));
 BUF_X4 _34978_ (.A(_09186_),
    .Z(_09272_));
 OR4_X2 _34979_ (.A1(_00156_),
    .A2(_09271_),
    .A3(_09232_),
    .A4(_09272_),
    .ZN(_09273_));
 OR2_X2 _34980_ (.A1(_09106_),
    .A2(_00155_),
    .ZN(_09274_));
 NAND3_X4 _34981_ (.A1(_09270_),
    .A2(_09273_),
    .A3(_09274_),
    .ZN(_09275_));
 BUF_X4 _34982_ (.A(_09146_),
    .Z(_09276_));
 NOR4_X2 _34983_ (.A1(_09276_),
    .A2(_09148_),
    .A3(_00154_),
    .A4(_09125_),
    .ZN(_09277_));
 NOR4_X2 _34984_ (.A1(_09237_),
    .A2(_09240_),
    .A3(_09241_),
    .A4(_00153_),
    .ZN(_09278_));
 NOR3_X4 _34985_ (.A1(_09275_),
    .A2(_09277_),
    .A3(_09278_),
    .ZN(_09279_));
 BUF_X4 _34986_ (.A(_09177_),
    .Z(_09280_));
 MUX2_X1 _34987_ (.A(_00152_),
    .B(_09279_),
    .S(_09280_),
    .Z(_09281_));
 AOI211_X2 _34988_ (.A(fe_queue_o[99]),
    .B(_09264_),
    .C1(_09223_),
    .C2(_09281_),
    .ZN(fe_queue_o[31]));
 NOR2_X1 _34989_ (.A1(_09195_),
    .A2(_00167_),
    .ZN(_09282_));
 AND3_X1 _34990_ (.A1(_09065_),
    .A2(\icache.data_set_select_mux.data_i [452]),
    .A3(_09069_),
    .ZN(_09283_));
 NOR4_X1 _34991_ (.A1(_09080_),
    .A2(_09085_),
    .A3(_09090_),
    .A4(_00166_),
    .ZN(_09284_));
 NOR3_X1 _34992_ (.A1(_09282_),
    .A2(_09283_),
    .A3(_09284_),
    .ZN(_09285_));
 OR4_X1 _34993_ (.A1(_00165_),
    .A2(_09136_),
    .A3(_09087_),
    .A4(_09092_),
    .ZN(_09286_));
 OR4_X2 _34994_ (.A1(_00164_),
    .A2(_09185_),
    .A3(_09097_),
    .A4(_09186_),
    .ZN(_09287_));
 AND3_X2 _34995_ (.A1(_09285_),
    .A2(_09286_),
    .A3(_09287_),
    .ZN(_09288_));
 OR2_X1 _34996_ (.A1(_09153_),
    .A2(_00163_),
    .ZN(_09289_));
 OR4_X1 _34997_ (.A1(_00162_),
    .A2(_09096_),
    .A3(_09232_),
    .A4(_09255_),
    .ZN(_09290_));
 NAND3_X1 _34998_ (.A1(_09288_),
    .A2(_09289_),
    .A3(_09290_),
    .ZN(_09291_));
 NOR4_X1 _34999_ (.A1(_09147_),
    .A2(_09259_),
    .A3(_09126_),
    .A4(_00161_),
    .ZN(_09292_));
 OAI21_X2 _35000_ (.A(_09245_),
    .B1(_09291_),
    .B2(_09292_),
    .ZN(_09293_));
 OR2_X1 _35001_ (.A1(_09041_),
    .A2(_00160_),
    .ZN(_09294_));
 AND3_X1 _35002_ (.A1(_09293_),
    .A2(_09262_),
    .A3(_09294_),
    .ZN(_09295_));
 NOR2_X1 _35003_ (.A1(_09074_),
    .A2(_00175_),
    .ZN(_09296_));
 AND3_X1 _35004_ (.A1(_09064_),
    .A2(\icache.data_set_select_mux.data_i [484]),
    .A3(_09067_),
    .ZN(_09297_));
 NOR4_X1 _35005_ (.A1(_09045_),
    .A2(_09083_),
    .A3(_09053_),
    .A4(_00174_),
    .ZN(_09298_));
 NOR3_X1 _35006_ (.A1(_09296_),
    .A2(_09297_),
    .A3(_09298_),
    .ZN(_09299_));
 OR4_X2 _35007_ (.A1(_00173_),
    .A2(_09045_),
    .A3(_09053_),
    .A4(_09047_),
    .ZN(_09300_));
 OR4_X1 _35008_ (.A1(_00172_),
    .A2(_09068_),
    .A3(_09083_),
    .A4(_09043_),
    .ZN(_09301_));
 AND3_X1 _35009_ (.A1(_09299_),
    .A2(_09300_),
    .A3(_09301_),
    .ZN(_09302_));
 MUX2_X2 _35010_ (.A(_00171_),
    .B(_09302_),
    .S(_09105_),
    .Z(_09303_));
 MUX2_X2 _35011_ (.A(_00170_),
    .B(_09303_),
    .S(_09061_),
    .Z(_09304_));
 OR4_X1 _35012_ (.A1(_00169_),
    .A2(_09146_),
    .A3(_09081_),
    .A4(_09113_),
    .ZN(_09305_));
 AND2_X2 _35013_ (.A1(_09304_),
    .A2(_09305_),
    .ZN(_09306_));
 MUX2_X1 _35014_ (.A(_00168_),
    .B(_09306_),
    .S(_09178_),
    .Z(_09307_));
 BUF_X8 _35015_ (.A(net1389),
    .Z(_09308_));
 AOI211_X2 _35016_ (.A(fe_queue_o[99]),
    .B(_09295_),
    .C1(_09307_),
    .C2(_09308_),
    .ZN(fe_queue_o[32]));
 NAND3_X1 _35017_ (.A1(_09129_),
    .A2(\icache.data_set_select_mux.data_i [453]),
    .A3(_09131_),
    .ZN(_09309_));
 OAI21_X2 _35018_ (.A(_09309_),
    .B1(_09133_),
    .B2(_00183_),
    .ZN(_09310_));
 AND2_X4 _35019_ (.A1(_09064_),
    .A2(_09202_),
    .ZN(_09311_));
 BUF_X4 _35020_ (.A(_09054_),
    .Z(_09312_));
 BUF_X4 _35021_ (.A(_09312_),
    .Z(_09313_));
 NOR4_X2 _35022_ (.A1(_09124_),
    .A2(_09201_),
    .A3(_09313_),
    .A4(_00182_),
    .ZN(_09314_));
 BUF_X4 _35023_ (.A(_09048_),
    .Z(_09315_));
 BUF_X8 _35024_ (.A(_09315_),
    .Z(_09316_));
 NOR4_X2 _35025_ (.A1(_09255_),
    .A2(_09313_),
    .A3(_09316_),
    .A4(_00181_),
    .ZN(_09317_));
 NOR4_X4 _35026_ (.A1(_09310_),
    .A2(_09311_),
    .A3(_09314_),
    .A4(_09317_),
    .ZN(_09318_));
 AND4_X1 _35027_ (.A1(_00180_),
    .A2(_09258_),
    .A3(_09113_),
    .A4(_09110_),
    .ZN(_09319_));
 OAI221_X2 _35028_ (.A(_09062_),
    .B1(_00179_),
    .B2(_09153_),
    .C1(_09318_),
    .C2(_09319_),
    .ZN(_09320_));
 NAND4_X4 _35029_ (.A1(_09111_),
    .A2(_09114_),
    .A3(_00178_),
    .A4(_09115_),
    .ZN(_09321_));
 AOI21_X4 _35030_ (.A(_09056_),
    .B1(_09320_),
    .B2(_09321_),
    .ZN(_09322_));
 BUF_X8 _35031_ (.A(_09049_),
    .Z(_09323_));
 AND3_X1 _35032_ (.A1(_09323_),
    .A2(_00177_),
    .A3(_09111_),
    .ZN(_09324_));
 OAI21_X1 _35033_ (.A(_09042_),
    .B1(_09322_),
    .B2(_09324_),
    .ZN(_09325_));
 NAND2_X2 _35034_ (.A1(_09118_),
    .A2(_00176_),
    .ZN(_09326_));
 AOI21_X2 _35035_ (.A(_09308_),
    .B1(_09325_),
    .B2(_09326_),
    .ZN(_09327_));
 NAND4_X2 _35036_ (.A1(_09148_),
    .A2(_00187_),
    .A3(_09259_),
    .A4(_09172_),
    .ZN(_09328_));
 BUF_X8 _35037_ (.A(_09065_),
    .Z(_09329_));
 NAND3_X2 _35038_ (.A1(_09329_),
    .A2(\icache.data_set_select_mux.data_i [485]),
    .A3(_09131_),
    .ZN(_09330_));
 OAI21_X4 _35039_ (.A(_09330_),
    .B1(_09133_),
    .B2(_00191_),
    .ZN(_09331_));
 BUF_X8 _35040_ (.A(_09123_),
    .Z(_09332_));
 NOR4_X2 _35041_ (.A1(_09086_),
    .A2(_09332_),
    .A3(_09138_),
    .A4(_00190_),
    .ZN(_09333_));
 BUF_X8 _35042_ (.A(_09092_),
    .Z(_09334_));
 NOR4_X2 _35043_ (.A1(_09137_),
    .A2(_09140_),
    .A3(_09334_),
    .A4(_00189_),
    .ZN(_09335_));
 NOR3_X4 _35044_ (.A1(_09331_),
    .A2(_09333_),
    .A3(_09335_),
    .ZN(_09336_));
 INV_X4 _35045_ (.A(_09311_),
    .ZN(_09337_));
 OAI21_X2 _35046_ (.A(_09336_),
    .B1(_00188_),
    .B2(_09337_),
    .ZN(_09338_));
 OAI21_X4 _35047_ (.A(_09328_),
    .B1(_09338_),
    .B2(_09103_),
    .ZN(_09339_));
 BUF_X8 _35048_ (.A(_09198_),
    .Z(_09340_));
 BUF_X4 _35049_ (.A(_09207_),
    .Z(_09341_));
 OR4_X2 _35050_ (.A1(_00186_),
    .A2(_09340_),
    .A3(_09135_),
    .A4(_09341_),
    .ZN(_09342_));
 BUF_X8 _35051_ (.A(_09316_),
    .Z(_09343_));
 OR4_X1 _35052_ (.A1(_00185_),
    .A2(_09340_),
    .A3(_09341_),
    .A4(_09343_),
    .ZN(_09344_));
 NAND4_X4 _35053_ (.A1(_09339_),
    .A2(_09042_),
    .A3(_09342_),
    .A4(_09344_),
    .ZN(_09345_));
 NAND2_X1 _35054_ (.A1(_09118_),
    .A2(_00184_),
    .ZN(_09346_));
 AOI21_X2 _35055_ (.A(_09039_),
    .B1(_09345_),
    .B2(_09346_),
    .ZN(_09347_));
 NOR3_X4 _35056_ (.A1(_09327_),
    .A2(fe_queue_o[99]),
    .A3(_09347_),
    .ZN(fe_queue_o[33]));
 BUF_X4 _35057_ (.A(_08644_),
    .Z(_09348_));
 AND3_X1 _35058_ (.A1(_09065_),
    .A2(\icache.data_set_select_mux.data_i [454]),
    .A3(_09069_),
    .ZN(_09349_));
 NOR4_X2 _35059_ (.A1(_09085_),
    .A2(_09254_),
    .A3(_09090_),
    .A4(_00198_),
    .ZN(_09350_));
 NOR4_X1 _35060_ (.A1(_09109_),
    .A2(_09112_),
    .A3(_00199_),
    .A4(_09100_),
    .ZN(_09351_));
 OR3_X1 _35061_ (.A1(_09349_),
    .A2(_09350_),
    .A3(_09351_),
    .ZN(_09352_));
 NOR4_X1 _35062_ (.A1(_09258_),
    .A2(_09091_),
    .A3(_09093_),
    .A4(_00197_),
    .ZN(_09353_));
 BUF_X8 _35063_ (.A(_09185_),
    .Z(_09354_));
 NOR4_X1 _35064_ (.A1(_09354_),
    .A2(_09086_),
    .A3(_00196_),
    .A4(_09101_),
    .ZN(_09355_));
 NOR3_X2 _35065_ (.A1(_09352_),
    .A2(_09353_),
    .A3(_09355_),
    .ZN(_09356_));
 OR4_X4 _35066_ (.A1(_00195_),
    .A2(_09070_),
    .A3(_09101_),
    .A4(_09093_),
    .ZN(_09357_));
 BUF_X8 _35067_ (.A(_09091_),
    .Z(_09358_));
 INV_X4 _35068_ (.A(_00194_),
    .ZN(_09359_));
 OAI211_X4 _35069_ (.A(_09115_),
    .B(_09358_),
    .C1(_09148_),
    .C2(_09359_),
    .ZN(_09360_));
 NAND3_X4 _35070_ (.A1(_09356_),
    .A2(_09357_),
    .A3(_09360_),
    .ZN(_09361_));
 NAND3_X1 _35071_ (.A1(_09323_),
    .A2(_00193_),
    .A3(_09111_),
    .ZN(_09362_));
 NAND3_X1 _35072_ (.A1(_09361_),
    .A2(_09245_),
    .A3(_09362_),
    .ZN(_09363_));
 OR2_X1 _35073_ (.A1(_09041_),
    .A2(_00192_),
    .ZN(_09364_));
 AND3_X1 _35074_ (.A1(_09363_),
    .A2(_09262_),
    .A3(_09364_),
    .ZN(_09365_));
 NAND3_X1 _35075_ (.A1(_09064_),
    .A2(\icache.data_set_select_mux.data_i [486]),
    .A3(_09068_),
    .ZN(_09366_));
 OAI21_X2 _35076_ (.A(_09366_),
    .B1(_09074_),
    .B2(_00207_),
    .ZN(_09367_));
 NOR4_X1 _35077_ (.A1(_09084_),
    .A2(_09079_),
    .A3(_09054_),
    .A4(_00206_),
    .ZN(_09368_));
 NOR4_X1 _35078_ (.A1(_09079_),
    .A2(_09054_),
    .A3(_09048_),
    .A4(_00205_),
    .ZN(_09369_));
 NOR3_X1 _35079_ (.A1(_09367_),
    .A2(_09368_),
    .A3(_09369_),
    .ZN(_09370_));
 OR4_X1 _35080_ (.A1(_00204_),
    .A2(_09068_),
    .A3(_09083_),
    .A4(_09099_),
    .ZN(_09371_));
 OR4_X1 _35081_ (.A1(_00203_),
    .A2(_09068_),
    .A3(_09099_),
    .A4(_09048_),
    .ZN(_09372_));
 AND3_X4 _35082_ (.A1(_09370_),
    .A2(_09371_),
    .A3(_09372_),
    .ZN(_09373_));
 MUX2_X2 _35083_ (.A(_00202_),
    .B(_09373_),
    .S(_09061_),
    .Z(_09374_));
 MUX2_X1 _35084_ (.A(_00201_),
    .B(_09374_),
    .S(_09057_),
    .Z(_09375_));
 MUX2_X1 _35085_ (.A(_00200_),
    .B(_09375_),
    .S(_09178_),
    .Z(_09376_));
 AOI211_X2 _35086_ (.A(_09348_),
    .B(_09365_),
    .C1(_09376_),
    .C2(_09308_),
    .ZN(fe_queue_o[34]));
 NOR2_X1 _35087_ (.A1(_09076_),
    .A2(_00215_),
    .ZN(_09377_));
 BUF_X4 _35088_ (.A(_09068_),
    .Z(_09378_));
 AND3_X1 _35089_ (.A1(_09128_),
    .A2(\icache.data_set_select_mux.data_i [455]),
    .A3(_09378_),
    .ZN(_09379_));
 NOR4_X2 _35090_ (.A1(_09123_),
    .A2(_09231_),
    .A3(_09312_),
    .A4(_00214_),
    .ZN(_09380_));
 NOR3_X1 _35091_ (.A1(_09377_),
    .A2(_09379_),
    .A3(_09380_),
    .ZN(_09381_));
 OR4_X2 _35092_ (.A1(_00213_),
    .A2(_09254_),
    .A3(_09312_),
    .A4(_09092_),
    .ZN(_09382_));
 OR4_X1 _35093_ (.A1(_00212_),
    .A2(_09378_),
    .A3(_09231_),
    .A4(_09100_),
    .ZN(_09383_));
 AND3_X1 _35094_ (.A1(_09381_),
    .A2(_09382_),
    .A3(_09383_),
    .ZN(_09384_));
 BUF_X4 _35095_ (.A(_09378_),
    .Z(_09385_));
 OR4_X2 _35096_ (.A1(_00211_),
    .A2(_09385_),
    .A3(_09149_),
    .A4(_09316_),
    .ZN(_09386_));
 AND3_X2 _35097_ (.A1(_09384_),
    .A2(_09062_),
    .A3(_09386_),
    .ZN(_09387_));
 AND3_X1 _35098_ (.A1(_09156_),
    .A2(_00210_),
    .A3(_09172_),
    .ZN(_09388_));
 OAI221_X2 _35099_ (.A(_09194_),
    .B1(_00209_),
    .B2(_09058_),
    .C1(_09387_),
    .C2(_09388_),
    .ZN(_09389_));
 NAND2_X1 _35100_ (.A1(_09220_),
    .A2(_00208_),
    .ZN(_09390_));
 AOI21_X1 _35101_ (.A(_09121_),
    .B1(_09389_),
    .B2(_09390_),
    .ZN(_09391_));
 NOR4_X2 _35102_ (.A1(_09147_),
    .A2(_09259_),
    .A3(_09126_),
    .A4(_00217_),
    .ZN(_09392_));
 NOR2_X1 _35103_ (.A1(_09075_),
    .A2(_00223_),
    .ZN(_09393_));
 AND2_X2 _35104_ (.A1(_09128_),
    .A2(_09130_),
    .ZN(_09394_));
 AOI21_X1 _35105_ (.A(_09393_),
    .B1(\icache.data_set_select_mux.data_i [487]),
    .B2(_09394_),
    .ZN(_09395_));
 OR4_X4 _35106_ (.A1(_00222_),
    .A2(_09231_),
    .A3(_09079_),
    .A4(_09202_),
    .ZN(_09396_));
 OR4_X4 _35107_ (.A1(_00221_),
    .A2(_09206_),
    .A3(_09202_),
    .A4(_09315_),
    .ZN(_09397_));
 AND4_X2 _35108_ (.A1(_09337_),
    .A2(_09395_),
    .A3(_09396_),
    .A4(_09397_),
    .ZN(_09398_));
 AND4_X1 _35109_ (.A1(_00220_),
    .A2(_09081_),
    .A3(_09113_),
    .A4(_09110_),
    .ZN(_09399_));
 OAI221_X2 _35110_ (.A(_09062_),
    .B1(_00219_),
    .B2(_09153_),
    .C1(_09398_),
    .C2(_09399_),
    .ZN(_09400_));
 NAND4_X4 _35111_ (.A1(_09111_),
    .A2(_09114_),
    .A3(_00218_),
    .A4(_09115_),
    .ZN(_09401_));
 AOI21_X4 _35112_ (.A(_09392_),
    .B1(_09400_),
    .B2(_09401_),
    .ZN(_09402_));
 MUX2_X1 _35113_ (.A(_00216_),
    .B(_09402_),
    .S(_09178_),
    .Z(_09403_));
 AOI211_X2 _35114_ (.A(_09348_),
    .B(_09391_),
    .C1(_09403_),
    .C2(_09308_),
    .ZN(fe_queue_o[35]));
 AND3_X1 _35115_ (.A1(_09197_),
    .A2(\icache.data_set_select_mux.data_i [456]),
    .A3(_09185_),
    .ZN(_09404_));
 NOR4_X2 _35116_ (.A1(_09238_),
    .A2(_09085_),
    .A3(_09087_),
    .A4(_00230_),
    .ZN(_09405_));
 NOR4_X1 _35117_ (.A1(_09109_),
    .A2(_09112_),
    .A3(_00231_),
    .A4(_09186_),
    .ZN(_09406_));
 NOR3_X1 _35118_ (.A1(_09404_),
    .A2(_09405_),
    .A3(_09406_),
    .ZN(_09407_));
 OR4_X2 _35119_ (.A1(_00229_),
    .A2(_09136_),
    .A3(_09087_),
    .A4(_09092_),
    .ZN(_09408_));
 OR4_X1 _35120_ (.A1(_00228_),
    .A2(_09185_),
    .A3(_09097_),
    .A4(_09186_),
    .ZN(_09409_));
 AND3_X2 _35121_ (.A1(_09407_),
    .A2(_09408_),
    .A3(_09409_),
    .ZN(_09410_));
 OR2_X4 _35122_ (.A1(_09153_),
    .A2(_00227_),
    .ZN(_09411_));
 OR4_X1 _35123_ (.A1(_00226_),
    .A2(_09096_),
    .A3(_09232_),
    .A4(_09255_),
    .ZN(_09412_));
 NAND3_X1 _35124_ (.A1(_09410_),
    .A2(_09411_),
    .A3(_09412_),
    .ZN(_09413_));
 NOR4_X1 _35125_ (.A1(_09147_),
    .A2(_09259_),
    .A3(_09126_),
    .A4(_00225_),
    .ZN(_09414_));
 OAI21_X2 _35126_ (.A(_09245_),
    .B1(_09413_),
    .B2(_09414_),
    .ZN(_09415_));
 OR2_X1 _35127_ (.A1(_09041_),
    .A2(_00224_),
    .ZN(_09416_));
 AND3_X1 _35128_ (.A1(_09415_),
    .A2(_09262_),
    .A3(_09416_),
    .ZN(_09417_));
 NAND3_X2 _35129_ (.A1(_09329_),
    .A2(\icache.data_set_select_mux.data_i [488]),
    .A3(_09230_),
    .ZN(_09418_));
 OAI21_X4 _35130_ (.A(_09418_),
    .B1(_09077_),
    .B2(_00239_),
    .ZN(_09419_));
 NOR4_X2 _35131_ (.A1(_09239_),
    .A2(_09267_),
    .A3(_09166_),
    .A4(_00238_),
    .ZN(_09420_));
 NOR4_X2 _35132_ (.A1(_09227_),
    .A2(_09088_),
    .A3(_09141_),
    .A4(_00237_),
    .ZN(_09421_));
 NOR3_X4 _35133_ (.A1(_09419_),
    .A2(_09420_),
    .A3(_09421_),
    .ZN(_09422_));
 OR4_X2 _35134_ (.A1(_00236_),
    .A2(_09271_),
    .A3(_09232_),
    .A4(_09272_),
    .ZN(_09423_));
 OR2_X1 _35135_ (.A1(_09106_),
    .A2(_00235_),
    .ZN(_09424_));
 NAND3_X4 _35136_ (.A1(_09422_),
    .A2(_09423_),
    .A3(_09424_),
    .ZN(_09425_));
 BUF_X4 _35137_ (.A(_09086_),
    .Z(_09426_));
 NOR4_X2 _35138_ (.A1(_09276_),
    .A2(_09426_),
    .A3(_00234_),
    .A4(_09125_),
    .ZN(_09427_));
 NOR4_X2 _35139_ (.A1(_09237_),
    .A2(_09240_),
    .A3(_09241_),
    .A4(_00233_),
    .ZN(_09428_));
 NOR3_X4 _35140_ (.A1(_09425_),
    .A2(_09427_),
    .A3(_09428_),
    .ZN(_09429_));
 MUX2_X1 _35141_ (.A(_00232_),
    .B(_09429_),
    .S(_09280_),
    .Z(_09430_));
 AOI211_X2 _35142_ (.A(_09348_),
    .B(_09417_),
    .C1(_09223_),
    .C2(_09430_),
    .ZN(fe_queue_o[36]));
 AND3_X1 _35143_ (.A1(_09129_),
    .A2(\icache.data_set_select_mux.data_i [457]),
    .A3(_09385_),
    .ZN(_09431_));
 BUF_X8 _35144_ (.A(_09231_),
    .Z(_09432_));
 NOR4_X2 _35145_ (.A1(_09332_),
    .A2(_09432_),
    .A3(_09313_),
    .A4(_00246_),
    .ZN(_09433_));
 NOR4_X1 _35146_ (.A1(_09140_),
    .A2(_09334_),
    .A3(_00247_),
    .A4(_09149_),
    .ZN(_09434_));
 NOR3_X2 _35147_ (.A1(_09431_),
    .A2(_09433_),
    .A3(_09434_),
    .ZN(_09435_));
 BUF_X8 _35148_ (.A(_09105_),
    .Z(_09436_));
 NOR2_X4 _35149_ (.A1(_09436_),
    .A2(_00243_),
    .ZN(_09437_));
 NOR2_X4 _35150_ (.A1(_09437_),
    .A2(_09214_),
    .ZN(_09438_));
 OR4_X4 _35151_ (.A1(_00245_),
    .A2(_09238_),
    .A3(_09203_),
    .A4(_09208_),
    .ZN(_09439_));
 OR4_X1 _35152_ (.A1(_00244_),
    .A2(_09145_),
    .A3(_09210_),
    .A4(_09211_),
    .ZN(_09440_));
 AND4_X2 _35153_ (.A1(_09435_),
    .A2(_09438_),
    .A3(_09439_),
    .A4(_09440_),
    .ZN(_09441_));
 AND4_X1 _35154_ (.A1(_00242_),
    .A2(_09217_),
    .A3(_09114_),
    .A4(_09115_),
    .ZN(_09442_));
 OAI221_X2 _35155_ (.A(_09194_),
    .B1(_00241_),
    .B2(_09058_),
    .C1(_09441_),
    .C2(_09442_),
    .ZN(_09443_));
 NAND2_X2 _35156_ (.A1(_09220_),
    .A2(_00240_),
    .ZN(_09444_));
 AOI21_X2 _35157_ (.A(_09121_),
    .B1(_09443_),
    .B2(_09444_),
    .ZN(_09445_));
 NAND3_X2 _35158_ (.A1(_09329_),
    .A2(\icache.data_set_select_mux.data_i [489]),
    .A3(_09230_),
    .ZN(_09446_));
 OAI21_X4 _35159_ (.A(_09446_),
    .B1(_09077_),
    .B2(_00255_),
    .ZN(_09447_));
 NOR4_X2 _35160_ (.A1(_09239_),
    .A2(_09267_),
    .A3(_09166_),
    .A4(_00254_),
    .ZN(_09448_));
 NOR4_X2 _35161_ (.A1(_09227_),
    .A2(_09088_),
    .A3(_09141_),
    .A4(_00253_),
    .ZN(_09449_));
 NOR3_X4 _35162_ (.A1(_09447_),
    .A2(_09448_),
    .A3(_09449_),
    .ZN(_09450_));
 OR4_X2 _35163_ (.A1(_00252_),
    .A2(_09271_),
    .A3(_09232_),
    .A4(_09272_),
    .ZN(_09451_));
 OR2_X2 _35164_ (.A1(_09106_),
    .A2(_00251_),
    .ZN(_09452_));
 NAND3_X4 _35165_ (.A1(_09450_),
    .A2(_09451_),
    .A3(_09452_),
    .ZN(_09453_));
 NOR4_X1 _35166_ (.A1(_09276_),
    .A2(_09426_),
    .A3(_00250_),
    .A4(_09125_),
    .ZN(_09454_));
 NOR4_X1 _35167_ (.A1(_09237_),
    .A2(_09240_),
    .A3(_09241_),
    .A4(_00249_),
    .ZN(_09455_));
 NOR3_X2 _35168_ (.A1(_09453_),
    .A2(_09454_),
    .A3(_09455_),
    .ZN(_09456_));
 MUX2_X1 _35169_ (.A(_00248_),
    .B(_09456_),
    .S(_09280_),
    .Z(_09457_));
 AOI211_X2 _35170_ (.A(_09348_),
    .B(_09445_),
    .C1(_09223_),
    .C2(_09457_),
    .ZN(fe_queue_o[37]));
 NAND3_X1 _35171_ (.A1(_09129_),
    .A2(\icache.data_set_select_mux.data_i [458]),
    .A3(_09385_),
    .ZN(_09458_));
 OAI21_X1 _35172_ (.A(_09458_),
    .B1(_09195_),
    .B2(_00263_),
    .ZN(_09459_));
 NOR4_X1 _35173_ (.A1(_09086_),
    .A2(_09255_),
    .A3(_09138_),
    .A4(_00262_),
    .ZN(_09460_));
 NOR4_X1 _35174_ (.A1(_09137_),
    .A2(_09138_),
    .A3(_09334_),
    .A4(_00261_),
    .ZN(_09461_));
 NOR3_X2 _35175_ (.A1(_09459_),
    .A2(_09460_),
    .A3(_09461_),
    .ZN(_09462_));
 OR4_X1 _35176_ (.A1(_00260_),
    .A2(_09385_),
    .A3(_09201_),
    .A4(_09149_),
    .ZN(_09463_));
 NOR4_X1 _35177_ (.A1(_09354_),
    .A2(_00259_),
    .A3(_09093_),
    .A4(_09149_),
    .ZN(_09464_));
 NOR2_X2 _35178_ (.A1(_09214_),
    .A2(_09464_),
    .ZN(_09465_));
 AND3_X2 _35179_ (.A1(_09462_),
    .A2(_09463_),
    .A3(_09465_),
    .ZN(_09466_));
 AND3_X1 _35180_ (.A1(_09156_),
    .A2(_00258_),
    .A3(_09172_),
    .ZN(_09467_));
 OAI221_X2 _35181_ (.A(_09194_),
    .B1(_00257_),
    .B2(_09058_),
    .C1(_09466_),
    .C2(_09467_),
    .ZN(_09468_));
 NAND2_X1 _35182_ (.A1(_09220_),
    .A2(_00256_),
    .ZN(_09469_));
 AOI21_X2 _35183_ (.A(_09121_),
    .B1(_09468_),
    .B2(_09469_),
    .ZN(_09470_));
 NOR2_X1 _35184_ (.A1(_09074_),
    .A2(_00271_),
    .ZN(_09471_));
 AND3_X1 _35185_ (.A1(_09063_),
    .A2(\icache.data_set_select_mux.data_i [490]),
    .A3(_09067_),
    .ZN(_09472_));
 NOR4_X1 _35186_ (.A1(_09045_),
    .A2(_09083_),
    .A3(_09053_),
    .A4(_00270_),
    .ZN(_09473_));
 NOR3_X1 _35187_ (.A1(_09471_),
    .A2(_09472_),
    .A3(_09473_),
    .ZN(_09474_));
 OR4_X2 _35188_ (.A1(_00269_),
    .A2(_09045_),
    .A3(_09053_),
    .A4(_09047_),
    .ZN(_09475_));
 OR4_X1 _35189_ (.A1(_00268_),
    .A2(_09067_),
    .A3(_09083_),
    .A4(_09043_),
    .ZN(_09476_));
 AND3_X1 _35190_ (.A1(_09474_),
    .A2(_09475_),
    .A3(_09476_),
    .ZN(_09477_));
 MUX2_X2 _35191_ (.A(_00267_),
    .B(_09477_),
    .S(_09105_),
    .Z(_09478_));
 MUX2_X2 _35192_ (.A(_00266_),
    .B(_09478_),
    .S(_09061_),
    .Z(_09479_));
 OR4_X1 _35193_ (.A1(_00265_),
    .A2(_09146_),
    .A3(_09081_),
    .A4(_09113_),
    .ZN(_09480_));
 AND2_X2 _35194_ (.A1(_09479_),
    .A2(_09480_),
    .ZN(_09481_));
 MUX2_X1 _35195_ (.A(_00264_),
    .B(_09481_),
    .S(_09178_),
    .Z(_09482_));
 AOI211_X2 _35196_ (.A(_09348_),
    .B(_09470_),
    .C1(_09482_),
    .C2(_09308_),
    .ZN(fe_queue_o[38]));
 NAND3_X1 _35197_ (.A1(_09197_),
    .A2(\icache.data_set_select_mux.data_i [459]),
    .A3(_09198_),
    .ZN(_09483_));
 OAI21_X2 _35198_ (.A(_09483_),
    .B1(_09195_),
    .B2(_00279_),
    .ZN(_09484_));
 NOR4_X1 _35199_ (.A1(_09098_),
    .A2(_09238_),
    .A3(_09203_),
    .A4(_00278_),
    .ZN(_09485_));
 NOR4_X1 _35200_ (.A1(_09255_),
    .A2(_09313_),
    .A3(_09208_),
    .A4(_00277_),
    .ZN(_09486_));
 OR3_X4 _35201_ (.A1(_09484_),
    .A2(_09485_),
    .A3(_09486_),
    .ZN(_09487_));
 NOR4_X2 _35202_ (.A1(_09340_),
    .A2(_09135_),
    .A3(_00276_),
    .A4(_09150_),
    .ZN(_09488_));
 OAI21_X2 _35203_ (.A(_09062_),
    .B1(_09153_),
    .B2(_00275_),
    .ZN(_09489_));
 NOR3_X4 _35204_ (.A1(_09487_),
    .A2(_09488_),
    .A3(_09489_),
    .ZN(_09490_));
 AND3_X1 _35205_ (.A1(_09156_),
    .A2(_00274_),
    .A3(_09172_),
    .ZN(_09491_));
 OAI221_X2 _35206_ (.A(_09194_),
    .B1(_00273_),
    .B2(_09058_),
    .C1(_09490_),
    .C2(_09491_),
    .ZN(_09492_));
 NAND2_X1 _35207_ (.A1(_09220_),
    .A2(_00272_),
    .ZN(_09493_));
 AOI21_X1 _35208_ (.A(_09121_),
    .B1(_09492_),
    .B2(_09493_),
    .ZN(_09494_));
 NAND3_X1 _35209_ (.A1(_09128_),
    .A2(\icache.data_set_select_mux.data_i [491]),
    .A3(_09378_),
    .ZN(_09495_));
 OAI21_X1 _35210_ (.A(_09495_),
    .B1(_09075_),
    .B2(_00287_),
    .ZN(_09496_));
 BUF_X4 _35211_ (.A(_09053_),
    .Z(_09497_));
 NOR4_X2 _35212_ (.A1(_09206_),
    .A2(_09084_),
    .A3(_09497_),
    .A4(_00286_),
    .ZN(_09498_));
 NOR4_X1 _35213_ (.A1(_09206_),
    .A2(_09497_),
    .A3(_09048_),
    .A4(_00285_),
    .ZN(_09499_));
 NOR4_X2 _35214_ (.A1(_09496_),
    .A2(_09311_),
    .A3(_09498_),
    .A4(_09499_),
    .ZN(_09500_));
 AND4_X1 _35215_ (.A1(_00284_),
    .A2(_09080_),
    .A3(_09112_),
    .A4(_09109_),
    .ZN(_09501_));
 OAI221_X2 _35216_ (.A(_09061_),
    .B1(_00283_),
    .B2(_09152_),
    .C1(_09500_),
    .C2(_09501_),
    .ZN(_09502_));
 NAND4_X1 _35217_ (.A1(_09110_),
    .A2(_09343_),
    .A3(_00282_),
    .A4(_09150_),
    .ZN(_09503_));
 NAND2_X2 _35218_ (.A1(_09502_),
    .A2(_09503_),
    .ZN(_09504_));
 MUX2_X2 _35219_ (.A(_00281_),
    .B(_09504_),
    .S(_09057_),
    .Z(_09505_));
 MUX2_X1 _35220_ (.A(_00280_),
    .B(_09505_),
    .S(_09178_),
    .Z(_09506_));
 AOI211_X2 _35221_ (.A(_09348_),
    .B(_09494_),
    .C1(_09506_),
    .C2(_09308_),
    .ZN(fe_queue_o[39]));
 AND3_X1 _35222_ (.A1(_09065_),
    .A2(\icache.data_set_select_mux.data_i [460]),
    .A3(_09185_),
    .ZN(_09507_));
 NOR4_X2 _35223_ (.A1(_09238_),
    .A2(_09085_),
    .A3(_09087_),
    .A4(_00294_),
    .ZN(_09508_));
 NOR4_X1 _35224_ (.A1(_09109_),
    .A2(_09112_),
    .A3(_00295_),
    .A4(_09186_),
    .ZN(_09509_));
 NOR3_X1 _35225_ (.A1(_09507_),
    .A2(_09508_),
    .A3(_09509_),
    .ZN(_09510_));
 OR4_X2 _35226_ (.A1(_00293_),
    .A2(_09136_),
    .A3(_09090_),
    .A4(_09092_),
    .ZN(_09511_));
 OR4_X1 _35227_ (.A1(_00292_),
    .A2(_09185_),
    .A3(_09097_),
    .A4(_09186_),
    .ZN(_09512_));
 AND3_X2 _35228_ (.A1(_09510_),
    .A2(_09511_),
    .A3(_09512_),
    .ZN(_09513_));
 OR2_X4 _35229_ (.A1(_09106_),
    .A2(_00291_),
    .ZN(_09514_));
 OR4_X1 _35230_ (.A1(_00290_),
    .A2(_09096_),
    .A3(_09232_),
    .A4(_09255_),
    .ZN(_09515_));
 NAND3_X1 _35231_ (.A1(_09513_),
    .A2(_09514_),
    .A3(_09515_),
    .ZN(_09516_));
 NOR4_X1 _35232_ (.A1(_09147_),
    .A2(_09259_),
    .A3(_09126_),
    .A4(_00289_),
    .ZN(_09517_));
 OAI21_X2 _35233_ (.A(_09245_),
    .B1(_09516_),
    .B2(_09517_),
    .ZN(_09518_));
 OR2_X1 _35234_ (.A1(_09177_),
    .A2(_00288_),
    .ZN(_09519_));
 AND3_X1 _35235_ (.A1(_09518_),
    .A2(_09262_),
    .A3(_09519_),
    .ZN(_09520_));
 NAND3_X2 _35236_ (.A1(_09329_),
    .A2(\icache.data_set_select_mux.data_i [492]),
    .A3(_09230_),
    .ZN(_09521_));
 OAI21_X4 _35237_ (.A(_09521_),
    .B1(_09077_),
    .B2(_00303_),
    .ZN(_09522_));
 NOR4_X2 _35238_ (.A1(_09239_),
    .A2(_09267_),
    .A3(_09166_),
    .A4(_00302_),
    .ZN(_09523_));
 NOR4_X2 _35239_ (.A1(_09227_),
    .A2(_09088_),
    .A3(_09141_),
    .A4(_00301_),
    .ZN(_09524_));
 NOR3_X4 _35240_ (.A1(_09522_),
    .A2(_09523_),
    .A3(_09524_),
    .ZN(_09525_));
 OR4_X2 _35241_ (.A1(_00300_),
    .A2(_09271_),
    .A3(_09232_),
    .A4(_09272_),
    .ZN(_09526_));
 OR2_X2 _35242_ (.A1(_09106_),
    .A2(_00299_),
    .ZN(_09527_));
 NAND3_X4 _35243_ (.A1(_09525_),
    .A2(_09526_),
    .A3(_09527_),
    .ZN(_09528_));
 NOR4_X2 _35244_ (.A1(_09276_),
    .A2(_09426_),
    .A3(_00298_),
    .A4(_09125_),
    .ZN(_09529_));
 NOR4_X2 _35245_ (.A1(_09237_),
    .A2(_09240_),
    .A3(_09241_),
    .A4(_00297_),
    .ZN(_09530_));
 NOR3_X4 _35246_ (.A1(_09528_),
    .A2(_09529_),
    .A3(_09530_),
    .ZN(_09531_));
 MUX2_X1 _35247_ (.A(_00296_),
    .B(_09531_),
    .S(_09280_),
    .Z(_09532_));
 AOI211_X2 _35248_ (.A(_09348_),
    .B(_09520_),
    .C1(_09223_),
    .C2(_09532_),
    .ZN(fe_queue_o[40]));
 OAI21_X1 _35249_ (.A(_09039_),
    .B1(_09042_),
    .B2(_00304_),
    .ZN(_09533_));
 NOR4_X1 _35250_ (.A1(_09122_),
    .A2(_09426_),
    .A3(_00306_),
    .A4(_09258_),
    .ZN(_09534_));
 NAND3_X1 _35251_ (.A1(_09329_),
    .A2(\icache.data_set_select_mux.data_i [461]),
    .A3(_09131_),
    .ZN(_09535_));
 OAI21_X2 _35252_ (.A(_09535_),
    .B1(_09133_),
    .B2(_00311_),
    .ZN(_09536_));
 NOR4_X2 _35253_ (.A1(_09086_),
    .A2(_09332_),
    .A3(_09138_),
    .A4(_00310_),
    .ZN(_09537_));
 NOR4_X2 _35254_ (.A1(_09137_),
    .A2(_09140_),
    .A3(_09334_),
    .A4(_00309_),
    .ZN(_09538_));
 NOR3_X4 _35255_ (.A1(_09536_),
    .A2(_09537_),
    .A3(_09538_),
    .ZN(_09539_));
 OR4_X1 _35256_ (.A1(_00308_),
    .A2(_09131_),
    .A3(_09432_),
    .A4(_09149_),
    .ZN(_09540_));
 NAND3_X2 _35257_ (.A1(_09539_),
    .A2(_09153_),
    .A3(_09540_),
    .ZN(_09541_));
 NAND3_X4 _35258_ (.A1(_09072_),
    .A2(_00307_),
    .A3(_09172_),
    .ZN(_09542_));
 AOI211_X2 _35259_ (.A(_09056_),
    .B(_09534_),
    .C1(_09541_),
    .C2(_09542_),
    .ZN(_09543_));
 AOI21_X2 _35260_ (.A(_09543_),
    .B1(_00305_),
    .B2(_09056_),
    .ZN(_09544_));
 AOI21_X2 _35261_ (.A(_09533_),
    .B1(_09544_),
    .B2(_09042_),
    .ZN(_09545_));
 NAND4_X2 _35262_ (.A1(_09148_),
    .A2(_00315_),
    .A3(_09259_),
    .A4(_09172_),
    .ZN(_09546_));
 NAND3_X2 _35263_ (.A1(_09129_),
    .A2(\icache.data_set_select_mux.data_i [493]),
    .A3(_09131_),
    .ZN(_09547_));
 OAI21_X4 _35264_ (.A(_09547_),
    .B1(_09133_),
    .B2(_00319_),
    .ZN(_09548_));
 NOR4_X2 _35265_ (.A1(_09086_),
    .A2(_09332_),
    .A3(_09138_),
    .A4(_00318_),
    .ZN(_09549_));
 NOR4_X2 _35266_ (.A1(_09137_),
    .A2(_09140_),
    .A3(_09334_),
    .A4(_00317_),
    .ZN(_09550_));
 NOR3_X4 _35267_ (.A1(_09548_),
    .A2(_09549_),
    .A3(_09550_),
    .ZN(_09551_));
 OAI21_X2 _35268_ (.A(_09551_),
    .B1(_00316_),
    .B2(_09337_),
    .ZN(_09552_));
 OAI21_X4 _35269_ (.A(_09546_),
    .B1(_09552_),
    .B2(_09103_),
    .ZN(_09553_));
 OR4_X2 _35270_ (.A1(_00314_),
    .A2(_09340_),
    .A3(_09135_),
    .A4(_09341_),
    .ZN(_09554_));
 OR4_X2 _35271_ (.A1(_00313_),
    .A2(_09340_),
    .A3(_09341_),
    .A4(_09343_),
    .ZN(_09555_));
 NAND4_X4 _35272_ (.A1(_09553_),
    .A2(_09042_),
    .A3(_09554_),
    .A4(_09555_),
    .ZN(_09556_));
 NAND2_X1 _35273_ (.A1(_09118_),
    .A2(_00312_),
    .ZN(_09557_));
 AOI21_X2 _35274_ (.A(_09039_),
    .B1(_09556_),
    .B2(_09557_),
    .ZN(_09558_));
 NOR3_X4 _35275_ (.A1(_09545_),
    .A2(fe_queue_o[99]),
    .A3(_09558_),
    .ZN(fe_queue_o[41]));
 NAND3_X1 _35276_ (.A1(_09323_),
    .A2(_00321_),
    .A3(_09217_),
    .ZN(_09559_));
 NOR2_X1 _35277_ (.A1(_09075_),
    .A2(_00327_),
    .ZN(_09560_));
 AND3_X1 _35278_ (.A1(_09128_),
    .A2(\icache.data_set_select_mux.data_i [462]),
    .A3(_09144_),
    .ZN(_09561_));
 NOR4_X1 _35279_ (.A1(_09254_),
    .A2(_09200_),
    .A3(_09497_),
    .A4(_00326_),
    .ZN(_09562_));
 NOR3_X1 _35280_ (.A1(_09560_),
    .A2(_09561_),
    .A3(_09562_),
    .ZN(_09563_));
 OR4_X2 _35281_ (.A1(_00325_),
    .A2(_09206_),
    .A3(_09202_),
    .A4(_09315_),
    .ZN(_09564_));
 OR4_X1 _35282_ (.A1(_00324_),
    .A2(_09144_),
    .A3(_09200_),
    .A4(_09099_),
    .ZN(_09565_));
 AND3_X1 _35283_ (.A1(_09563_),
    .A2(_09564_),
    .A3(_09565_),
    .ZN(_09566_));
 OR2_X2 _35284_ (.A1(_09152_),
    .A2(_00323_),
    .ZN(_09567_));
 OR4_X2 _35285_ (.A1(_00322_),
    .A2(_09145_),
    .A3(_09210_),
    .A4(_09080_),
    .ZN(_09568_));
 NAND3_X4 _35286_ (.A1(_09566_),
    .A2(_09567_),
    .A3(_09568_),
    .ZN(_09569_));
 OAI211_X1 _35287_ (.A(_09177_),
    .B(_09559_),
    .C1(_09569_),
    .C2(_09056_),
    .ZN(_09570_));
 BUF_X4 _35288_ (.A(_09040_),
    .Z(_09571_));
 NOR2_X1 _35289_ (.A1(_09571_),
    .A2(_00320_),
    .ZN(_09572_));
 NOR2_X1 _35290_ (.A1(_09572_),
    .A2(net1389),
    .ZN(_09573_));
 NOR2_X1 _35291_ (.A1(_09075_),
    .A2(_00335_),
    .ZN(_09574_));
 AND3_X1 _35292_ (.A1(_09064_),
    .A2(\icache.data_set_select_mux.data_i [494]),
    .A3(_09068_),
    .ZN(_09575_));
 NOR4_X1 _35293_ (.A1(_09079_),
    .A2(_09084_),
    .A3(_09054_),
    .A4(_00334_),
    .ZN(_09576_));
 NOR3_X1 _35294_ (.A1(_09574_),
    .A2(_09575_),
    .A3(_09576_),
    .ZN(_09577_));
 OR4_X1 _35295_ (.A1(_00333_),
    .A2(_09079_),
    .A3(_09054_),
    .A4(_09048_),
    .ZN(_09578_));
 OR4_X1 _35296_ (.A1(_00332_),
    .A2(_09068_),
    .A3(_09084_),
    .A4(_09099_),
    .ZN(_09579_));
 AND3_X1 _35297_ (.A1(_09577_),
    .A2(_09578_),
    .A3(_09579_),
    .ZN(_09580_));
 OR2_X1 _35298_ (.A1(_09152_),
    .A2(_00331_),
    .ZN(_09581_));
 NAND2_X4 _35299_ (.A1(_09580_),
    .A2(_09581_),
    .ZN(_09582_));
 NOR4_X2 _35300_ (.A1(_09354_),
    .A2(_09098_),
    .A3(_00330_),
    .A4(_09207_),
    .ZN(_09583_));
 NOR4_X2 _35301_ (.A1(_09354_),
    .A2(_09124_),
    .A3(_09141_),
    .A4(_00329_),
    .ZN(_09584_));
 NOR3_X4 _35302_ (.A1(_09582_),
    .A2(_09583_),
    .A3(_09584_),
    .ZN(_09585_));
 MUX2_X1 _35303_ (.A(_00328_),
    .B(_09585_),
    .S(_09571_),
    .Z(_09586_));
 BUF_X4 _35304_ (.A(net1389),
    .Z(_09587_));
 AOI221_X4 _35305_ (.A(_08644_),
    .B1(_09570_),
    .B2(_09573_),
    .C1(_09586_),
    .C2(_09587_),
    .ZN(fe_queue_o[42]));
 NAND4_X2 _35306_ (.A1(_09148_),
    .A2(_00339_),
    .A3(_09259_),
    .A4(_09172_),
    .ZN(_09588_));
 NAND3_X2 _35307_ (.A1(_09197_),
    .A2(\icache.data_set_select_mux.data_i [463]),
    .A3(_09198_),
    .ZN(_09589_));
 OAI21_X4 _35308_ (.A(_09589_),
    .B1(_09195_),
    .B2(_00343_),
    .ZN(_09590_));
 NOR4_X2 _35309_ (.A1(_09267_),
    .A2(_09207_),
    .A3(_09313_),
    .A4(_00342_),
    .ZN(_09591_));
 NOR4_X2 _35310_ (.A1(_09332_),
    .A2(_09138_),
    .A3(_09316_),
    .A4(_00341_),
    .ZN(_09592_));
 NOR3_X4 _35311_ (.A1(_09590_),
    .A2(_09591_),
    .A3(_09592_),
    .ZN(_09593_));
 OAI21_X2 _35312_ (.A(_09593_),
    .B1(_00340_),
    .B2(_09337_),
    .ZN(_09594_));
 OAI21_X4 _35313_ (.A(_09588_),
    .B1(_09594_),
    .B2(_09103_),
    .ZN(_09595_));
 OR4_X4 _35314_ (.A1(_00338_),
    .A2(_09340_),
    .A3(_09135_),
    .A4(_09258_),
    .ZN(_09596_));
 OR4_X2 _35315_ (.A1(_00337_),
    .A2(_09146_),
    .A3(_09258_),
    .A4(_09343_),
    .ZN(_09597_));
 NAND4_X4 _35316_ (.A1(_09595_),
    .A2(_09194_),
    .A3(_09596_),
    .A4(_09597_),
    .ZN(_09598_));
 NAND2_X1 _35317_ (.A1(_09220_),
    .A2(_00336_),
    .ZN(_09599_));
 AOI21_X1 _35318_ (.A(_09121_),
    .B1(_09598_),
    .B2(_09599_),
    .ZN(_09600_));
 NAND3_X1 _35319_ (.A1(_09128_),
    .A2(\icache.data_set_select_mux.data_i [495]),
    .A3(_09378_),
    .ZN(_09601_));
 OAI21_X1 _35320_ (.A(_09601_),
    .B1(_09075_),
    .B2(_00351_),
    .ZN(_09602_));
 NOR4_X1 _35321_ (.A1(_09206_),
    .A2(_09084_),
    .A3(_09497_),
    .A4(_00350_),
    .ZN(_09603_));
 NOR4_X2 _35322_ (.A1(_09079_),
    .A2(_09497_),
    .A3(_09048_),
    .A4(_00349_),
    .ZN(_09604_));
 NOR4_X2 _35323_ (.A1(_09602_),
    .A2(_09311_),
    .A3(_09603_),
    .A4(_09604_),
    .ZN(_09605_));
 AND4_X1 _35324_ (.A1(_00348_),
    .A2(_09136_),
    .A3(_09112_),
    .A4(_09109_),
    .ZN(_09606_));
 OAI221_X2 _35325_ (.A(_09061_),
    .B1(_00347_),
    .B2(_09152_),
    .C1(_09605_),
    .C2(_09606_),
    .ZN(_09607_));
 NAND4_X1 _35326_ (.A1(_09110_),
    .A2(_09343_),
    .A3(_00346_),
    .A4(_09150_),
    .ZN(_09608_));
 NAND2_X2 _35327_ (.A1(_09607_),
    .A2(_09608_),
    .ZN(_09609_));
 MUX2_X2 _35328_ (.A(_00345_),
    .B(_09609_),
    .S(_09057_),
    .Z(_09610_));
 MUX2_X1 _35329_ (.A(_00344_),
    .B(_09610_),
    .S(_09178_),
    .Z(_09611_));
 AOI211_X2 _35330_ (.A(_09348_),
    .B(_09600_),
    .C1(_09611_),
    .C2(_09308_),
    .ZN(fe_queue_o[43]));
 NOR2_X2 _35331_ (.A1(_09195_),
    .A2(_00359_),
    .ZN(_09612_));
 AND3_X1 _35332_ (.A1(_09197_),
    .A2(\icache.data_set_select_mux.data_i [464]),
    .A3(_09198_),
    .ZN(_09613_));
 NOR4_X4 _35333_ (.A1(_09124_),
    .A2(_09201_),
    .A3(_09203_),
    .A4(_00358_),
    .ZN(_09614_));
 NOR3_X4 _35334_ (.A1(_09612_),
    .A2(_09613_),
    .A3(_09614_),
    .ZN(_09615_));
 OR4_X4 _35335_ (.A1(_00357_),
    .A2(_09207_),
    .A3(_09203_),
    .A4(_09208_),
    .ZN(_09616_));
 OR4_X1 _35336_ (.A1(_00356_),
    .A2(_09198_),
    .A3(_09210_),
    .A4(_09211_),
    .ZN(_09617_));
 NOR2_X2 _35337_ (.A1(_09152_),
    .A2(_00355_),
    .ZN(_09618_));
 NOR2_X4 _35338_ (.A1(_09618_),
    .A2(_09060_),
    .ZN(_09619_));
 AND4_X2 _35339_ (.A1(_09615_),
    .A2(_09616_),
    .A3(_09617_),
    .A4(_09619_),
    .ZN(_09620_));
 AND4_X1 _35340_ (.A1(_00354_),
    .A2(_09217_),
    .A3(_09114_),
    .A4(_09115_),
    .ZN(_09621_));
 OAI221_X2 _35341_ (.A(_09194_),
    .B1(_00353_),
    .B2(_09058_),
    .C1(_09620_),
    .C2(_09621_),
    .ZN(_09622_));
 NAND2_X1 _35342_ (.A1(_09220_),
    .A2(_00352_),
    .ZN(_09623_));
 AOI21_X2 _35343_ (.A(_09587_),
    .B1(_09622_),
    .B2(_09623_),
    .ZN(_09624_));
 NAND3_X2 _35344_ (.A1(_09329_),
    .A2(\icache.data_set_select_mux.data_i [496]),
    .A3(_09230_),
    .ZN(_09625_));
 OAI21_X4 _35345_ (.A(_09625_),
    .B1(_09077_),
    .B2(_00367_),
    .ZN(_09626_));
 NOR4_X2 _35346_ (.A1(_09239_),
    .A2(_09267_),
    .A3(_09166_),
    .A4(_00366_),
    .ZN(_09627_));
 NOR4_X2 _35347_ (.A1(_09227_),
    .A2(_09088_),
    .A3(_09141_),
    .A4(_00365_),
    .ZN(_09628_));
 NOR3_X4 _35348_ (.A1(_09626_),
    .A2(_09627_),
    .A3(_09628_),
    .ZN(_09629_));
 OR4_X2 _35349_ (.A1(_00364_),
    .A2(_09271_),
    .A3(_09432_),
    .A4(_09272_),
    .ZN(_09630_));
 OR2_X2 _35350_ (.A1(_09106_),
    .A2(_00363_),
    .ZN(_09631_));
 NAND3_X4 _35351_ (.A1(_09629_),
    .A2(_09630_),
    .A3(_09631_),
    .ZN(_09632_));
 NOR4_X2 _35352_ (.A1(_09276_),
    .A2(_09426_),
    .A3(_00362_),
    .A4(_09125_),
    .ZN(_09633_));
 NOR4_X2 _35353_ (.A1(_09237_),
    .A2(_09240_),
    .A3(_09241_),
    .A4(_00361_),
    .ZN(_09634_));
 NOR3_X4 _35354_ (.A1(_09632_),
    .A2(_09633_),
    .A3(_09634_),
    .ZN(_09635_));
 MUX2_X1 _35355_ (.A(_00360_),
    .B(_09635_),
    .S(_09280_),
    .Z(_09636_));
 AOI211_X2 _35356_ (.A(_09348_),
    .B(_09624_),
    .C1(_09223_),
    .C2(_09636_),
    .ZN(fe_queue_o[44]));
 AND3_X1 _35357_ (.A1(_09129_),
    .A2(\icache.data_set_select_mux.data_i [465]),
    .A3(_09385_),
    .ZN(_09637_));
 NOR4_X2 _35358_ (.A1(_09332_),
    .A2(_09432_),
    .A3(_09313_),
    .A4(_00374_),
    .ZN(_09638_));
 NOR4_X1 _35359_ (.A1(_09140_),
    .A2(_09316_),
    .A3(_00375_),
    .A4(_09149_),
    .ZN(_09639_));
 NOR3_X2 _35360_ (.A1(_09637_),
    .A2(_09638_),
    .A3(_09639_),
    .ZN(_09640_));
 NOR2_X4 _35361_ (.A1(_09436_),
    .A2(_00371_),
    .ZN(_09641_));
 NOR2_X4 _35362_ (.A1(_09641_),
    .A2(_09214_),
    .ZN(_09642_));
 OR4_X4 _35363_ (.A1(_00373_),
    .A2(_09238_),
    .A3(_09203_),
    .A4(_09208_),
    .ZN(_09643_));
 OR4_X1 _35364_ (.A1(_00372_),
    .A2(_09145_),
    .A3(_09210_),
    .A4(_09211_),
    .ZN(_09644_));
 AND4_X2 _35365_ (.A1(_09640_),
    .A2(_09642_),
    .A3(_09643_),
    .A4(_09644_),
    .ZN(_09645_));
 AND4_X1 _35366_ (.A1(_00370_),
    .A2(_09217_),
    .A3(_09114_),
    .A4(_09150_),
    .ZN(_09646_));
 OAI221_X2 _35367_ (.A(_09194_),
    .B1(_00369_),
    .B2(_09057_),
    .C1(_09645_),
    .C2(_09646_),
    .ZN(_09647_));
 NAND2_X1 _35368_ (.A1(_09220_),
    .A2(_00368_),
    .ZN(_09648_));
 AOI21_X1 _35369_ (.A(_09587_),
    .B1(_09647_),
    .B2(_09648_),
    .ZN(_09649_));
 NAND3_X2 _35370_ (.A1(_09329_),
    .A2(\icache.data_set_select_mux.data_i [497]),
    .A3(_09230_),
    .ZN(_09650_));
 OAI21_X4 _35371_ (.A(_09650_),
    .B1(_09077_),
    .B2(_00383_),
    .ZN(_09651_));
 NOR4_X2 _35372_ (.A1(_09239_),
    .A2(_09267_),
    .A3(_09166_),
    .A4(_00382_),
    .ZN(_09652_));
 NOR4_X2 _35373_ (.A1(_09227_),
    .A2(_09088_),
    .A3(_09141_),
    .A4(_00381_),
    .ZN(_09653_));
 NOR3_X4 _35374_ (.A1(_09651_),
    .A2(_09652_),
    .A3(_09653_),
    .ZN(_09654_));
 OR4_X2 _35375_ (.A1(_00380_),
    .A2(_09271_),
    .A3(_09432_),
    .A4(_09272_),
    .ZN(_09655_));
 OR2_X2 _35376_ (.A1(_09106_),
    .A2(_00379_),
    .ZN(_09656_));
 NAND3_X4 _35377_ (.A1(_09654_),
    .A2(_09655_),
    .A3(_09656_),
    .ZN(_09657_));
 NOR4_X2 _35378_ (.A1(_09276_),
    .A2(_09426_),
    .A3(_00378_),
    .A4(_09125_),
    .ZN(_09658_));
 NOR4_X2 _35379_ (.A1(_09237_),
    .A2(_09240_),
    .A3(_09241_),
    .A4(_00377_),
    .ZN(_09659_));
 NOR3_X4 _35380_ (.A1(_09657_),
    .A2(_09658_),
    .A3(_09659_),
    .ZN(_09660_));
 MUX2_X1 _35381_ (.A(_00376_),
    .B(_09660_),
    .S(_09280_),
    .Z(_09661_));
 AOI211_X2 _35382_ (.A(_09348_),
    .B(_09649_),
    .C1(_09223_),
    .C2(_09661_),
    .ZN(fe_queue_o[45]));
 NOR2_X1 _35383_ (.A1(_09076_),
    .A2(_00391_),
    .ZN(_09662_));
 AND3_X1 _35384_ (.A1(_09128_),
    .A2(\icache.data_set_select_mux.data_i [466]),
    .A3(_09378_),
    .ZN(_09663_));
 NOR4_X1 _35385_ (.A1(_09254_),
    .A2(_09231_),
    .A3(_09202_),
    .A4(_00390_),
    .ZN(_09664_));
 NOR3_X1 _35386_ (.A1(_09662_),
    .A2(_09663_),
    .A3(_09664_),
    .ZN(_09665_));
 OR4_X2 _35387_ (.A1(_00389_),
    .A2(_09254_),
    .A3(_09312_),
    .A4(_09315_),
    .ZN(_09666_));
 OR4_X1 _35388_ (.A1(_00388_),
    .A2(_09378_),
    .A3(_09200_),
    .A4(_09100_),
    .ZN(_09667_));
 AND3_X2 _35389_ (.A1(_09665_),
    .A2(_09666_),
    .A3(_09667_),
    .ZN(_09668_));
 OR2_X2 _35390_ (.A1(_09436_),
    .A2(_00387_),
    .ZN(_09669_));
 OR4_X4 _35391_ (.A1(_00386_),
    .A2(_09198_),
    .A3(_09201_),
    .A4(_09238_),
    .ZN(_09670_));
 NAND3_X2 _35392_ (.A1(_09668_),
    .A2(_09669_),
    .A3(_09670_),
    .ZN(_09671_));
 NOR4_X1 _35393_ (.A1(_09122_),
    .A2(_09341_),
    .A3(_09343_),
    .A4(_00385_),
    .ZN(_09672_));
 OAI21_X1 _35394_ (.A(_09041_),
    .B1(_09671_),
    .B2(_09672_),
    .ZN(_09673_));
 NOR2_X1 _35395_ (.A1(_09571_),
    .A2(_00384_),
    .ZN(_09674_));
 NOR2_X1 _35396_ (.A1(_09674_),
    .A2(net1389),
    .ZN(_09675_));
 NOR2_X1 _35397_ (.A1(_09074_),
    .A2(_00399_),
    .ZN(_09676_));
 AND3_X1 _35398_ (.A1(_09063_),
    .A2(\icache.data_set_select_mux.data_i [498]),
    .A3(_09067_),
    .ZN(_09677_));
 NOR4_X1 _35399_ (.A1(_09044_),
    .A2(_09082_),
    .A3(_09052_),
    .A4(_00398_),
    .ZN(_09678_));
 NOR3_X1 _35400_ (.A1(_09676_),
    .A2(_09677_),
    .A3(_09678_),
    .ZN(_09679_));
 OR4_X1 _35401_ (.A1(_00397_),
    .A2(_09044_),
    .A3(_09052_),
    .A4(_09047_),
    .ZN(_09680_));
 OR4_X1 _35402_ (.A1(_00396_),
    .A2(_09067_),
    .A3(_09082_),
    .A4(_09043_),
    .ZN(_09681_));
 AND3_X1 _35403_ (.A1(_09679_),
    .A2(_09680_),
    .A3(_09681_),
    .ZN(_09682_));
 MUX2_X2 _35404_ (.A(_00395_),
    .B(_09682_),
    .S(_09104_),
    .Z(_09683_));
 MUX2_X2 _35405_ (.A(_00394_),
    .B(_09683_),
    .S(_09061_),
    .Z(_09684_));
 OR4_X1 _35406_ (.A1(_00393_),
    .A2(_09185_),
    .A3(_09123_),
    .A4(_09112_),
    .ZN(_09685_));
 AND2_X2 _35407_ (.A1(_09684_),
    .A2(_09685_),
    .ZN(_09686_));
 MUX2_X1 _35408_ (.A(_00392_),
    .B(_09686_),
    .S(_09571_),
    .Z(_09687_));
 AOI221_X4 _35409_ (.A(_08644_),
    .B1(_09673_),
    .B2(_09675_),
    .C1(_09687_),
    .C2(_09587_),
    .ZN(fe_queue_o[46]));
 BUF_X16 _35410_ (.A(_08643_),
    .Z(_09688_));
 NOR2_X1 _35411_ (.A1(_09076_),
    .A2(_00407_),
    .ZN(_09689_));
 AND3_X1 _35412_ (.A1(_09065_),
    .A2(\icache.data_set_select_mux.data_i [467]),
    .A3(_09069_),
    .ZN(_09690_));
 NOR4_X1 _35413_ (.A1(_09080_),
    .A2(_09085_),
    .A3(_09090_),
    .A4(_00406_),
    .ZN(_09691_));
 NOR3_X1 _35414_ (.A1(_09689_),
    .A2(_09690_),
    .A3(_09691_),
    .ZN(_09692_));
 OR4_X1 _35415_ (.A1(_00405_),
    .A2(_09136_),
    .A3(_09090_),
    .A4(_09092_),
    .ZN(_09693_));
 OR4_X2 _35416_ (.A1(_00404_),
    .A2(_09185_),
    .A3(_09097_),
    .A4(_09186_),
    .ZN(_09694_));
 AND3_X2 _35417_ (.A1(_09692_),
    .A2(_09693_),
    .A3(_09694_),
    .ZN(_09695_));
 OR2_X4 _35418_ (.A1(_09106_),
    .A2(_00403_),
    .ZN(_09696_));
 OR4_X1 _35419_ (.A1(_00402_),
    .A2(_09096_),
    .A3(_09232_),
    .A4(_09255_),
    .ZN(_09697_));
 NAND3_X1 _35420_ (.A1(_09695_),
    .A2(_09696_),
    .A3(_09697_),
    .ZN(_09698_));
 NOR4_X1 _35421_ (.A1(_09147_),
    .A2(_09259_),
    .A3(_09126_),
    .A4(_00401_),
    .ZN(_09699_));
 OAI21_X1 _35422_ (.A(_09245_),
    .B1(_09698_),
    .B2(_09699_),
    .ZN(_09700_));
 OR2_X1 _35423_ (.A1(_09177_),
    .A2(_00400_),
    .ZN(_09701_));
 AND3_X1 _35424_ (.A1(_09700_),
    .A2(_09262_),
    .A3(_09701_),
    .ZN(_09702_));
 NAND3_X2 _35425_ (.A1(_09329_),
    .A2(\icache.data_set_select_mux.data_i [499]),
    .A3(_09230_),
    .ZN(_09703_));
 OAI21_X4 _35426_ (.A(_09703_),
    .B1(_09133_),
    .B2(_00415_),
    .ZN(_09704_));
 NOR4_X2 _35427_ (.A1(_09239_),
    .A2(_09267_),
    .A3(_09166_),
    .A4(_00414_),
    .ZN(_09705_));
 NOR4_X2 _35428_ (.A1(_09227_),
    .A2(_09088_),
    .A3(_09141_),
    .A4(_00413_),
    .ZN(_09706_));
 NOR3_X4 _35429_ (.A1(_09704_),
    .A2(_09705_),
    .A3(_09706_),
    .ZN(_09707_));
 OR4_X2 _35430_ (.A1(_00412_),
    .A2(_09271_),
    .A3(_09432_),
    .A4(_09272_),
    .ZN(_09708_));
 OR2_X1 _35431_ (.A1(_09436_),
    .A2(_00411_),
    .ZN(_09709_));
 NAND3_X4 _35432_ (.A1(_09707_),
    .A2(_09708_),
    .A3(_09709_),
    .ZN(_09710_));
 NOR4_X1 _35433_ (.A1(_09276_),
    .A2(_09426_),
    .A3(_00410_),
    .A4(_09125_),
    .ZN(_09711_));
 NOR4_X1 _35434_ (.A1(_09237_),
    .A2(_09240_),
    .A3(_09241_),
    .A4(_00409_),
    .ZN(_09712_));
 NOR3_X2 _35435_ (.A1(_09710_),
    .A2(_09711_),
    .A3(_09712_),
    .ZN(_09713_));
 MUX2_X1 _35436_ (.A(_00408_),
    .B(_09713_),
    .S(_09280_),
    .Z(_09714_));
 AOI211_X2 _35437_ (.A(_09688_),
    .B(_09702_),
    .C1(_09223_),
    .C2(_09714_),
    .ZN(fe_queue_o[47]));
 AND3_X1 _35438_ (.A1(_09059_),
    .A2(_00426_),
    .A3(_09091_),
    .ZN(_09715_));
 NOR2_X1 _35439_ (.A1(_09076_),
    .A2(_00431_),
    .ZN(_09716_));
 AND3_X1 _35440_ (.A1(_09128_),
    .A2(\icache.data_set_select_mux.data_i [500]),
    .A3(_09378_),
    .ZN(_09717_));
 NOR4_X1 _35441_ (.A1(_09254_),
    .A2(_09200_),
    .A3(_09497_),
    .A4(_00430_),
    .ZN(_09718_));
 NOR3_X1 _35442_ (.A1(_09716_),
    .A2(_09717_),
    .A3(_09718_),
    .ZN(_09719_));
 OR4_X4 _35443_ (.A1(_00429_),
    .A2(_09206_),
    .A3(_09202_),
    .A4(_09315_),
    .ZN(_09720_));
 OR4_X1 _35444_ (.A1(_00428_),
    .A2(_09378_),
    .A3(_09200_),
    .A4(_09100_),
    .ZN(_09721_));
 AND3_X1 _35445_ (.A1(_09719_),
    .A2(_09720_),
    .A3(_09721_),
    .ZN(_09722_));
 NOR4_X1 _35446_ (.A1(_09131_),
    .A2(_00427_),
    .A3(_09316_),
    .A4(_09149_),
    .ZN(_09723_));
 NOR2_X1 _35447_ (.A1(_09214_),
    .A2(_09723_),
    .ZN(_09724_));
 AOI21_X4 _35448_ (.A(_09715_),
    .B1(_09722_),
    .B2(_09724_),
    .ZN(_09725_));
 NOR4_X2 _35449_ (.A1(_09122_),
    .A2(_09258_),
    .A3(_09343_),
    .A4(_00425_),
    .ZN(_09726_));
 OAI21_X4 _35450_ (.A(_09041_),
    .B1(_09725_),
    .B2(_09726_),
    .ZN(_09727_));
 NOR2_X1 _35451_ (.A1(_09571_),
    .A2(_00424_),
    .ZN(_09728_));
 NOR2_X1 _35452_ (.A1(_09728_),
    .A2(_09038_),
    .ZN(_09729_));
 NAND3_X1 _35453_ (.A1(_09065_),
    .A2(\icache.data_set_select_mux.data_i [468]),
    .A3(_09130_),
    .ZN(_09730_));
 OAI21_X2 _35454_ (.A(_09730_),
    .B1(_09076_),
    .B2(_00423_),
    .ZN(_09731_));
 NOR4_X2 _35455_ (.A1(_09136_),
    .A2(_09097_),
    .A3(_09312_),
    .A4(_00422_),
    .ZN(_09732_));
 NOR4_X2 _35456_ (.A1(_09123_),
    .A2(_09090_),
    .A3(_09092_),
    .A4(_00421_),
    .ZN(_09733_));
 NOR3_X4 _35457_ (.A1(_09731_),
    .A2(_09732_),
    .A3(_09733_),
    .ZN(_09734_));
 OR4_X1 _35458_ (.A1(_00420_),
    .A2(_09130_),
    .A3(_09231_),
    .A4(_09100_),
    .ZN(_09735_));
 OR2_X1 _35459_ (.A1(_09105_),
    .A2(_00419_),
    .ZN(_09736_));
 NAND3_X2 _35460_ (.A1(_09734_),
    .A2(_09735_),
    .A3(_09736_),
    .ZN(_09737_));
 NOR4_X4 _35461_ (.A1(_09354_),
    .A2(_09098_),
    .A3(_00418_),
    .A4(_09207_),
    .ZN(_09738_));
 NOR4_X1 _35462_ (.A1(_09070_),
    .A2(_09124_),
    .A3(_09334_),
    .A4(_00417_),
    .ZN(_09739_));
 NOR3_X2 _35463_ (.A1(_09737_),
    .A2(_09738_),
    .A3(_09739_),
    .ZN(_09740_));
 MUX2_X1 _35464_ (.A(_00416_),
    .B(_09740_),
    .S(_09571_),
    .Z(_09741_));
 AOI221_X4 _35465_ (.A(_08644_),
    .B1(_09727_),
    .B2(_09729_),
    .C1(_09741_),
    .C2(_09039_),
    .ZN(fe_queue_o[48]));
 NAND3_X2 _35466_ (.A1(_09323_),
    .A2(_00441_),
    .A3(_09217_),
    .ZN(_09742_));
 NOR2_X1 _35467_ (.A1(_09075_),
    .A2(_00447_),
    .ZN(_09743_));
 AND3_X1 _35468_ (.A1(_09064_),
    .A2(\icache.data_set_select_mux.data_i [501]),
    .A3(_09144_),
    .ZN(_09744_));
 NOR4_X1 _35469_ (.A1(_09254_),
    .A2(_09200_),
    .A3(_09497_),
    .A4(_00446_),
    .ZN(_09745_));
 NOR3_X1 _35470_ (.A1(_09743_),
    .A2(_09744_),
    .A3(_09745_),
    .ZN(_09746_));
 OR4_X2 _35471_ (.A1(_00445_),
    .A2(_09206_),
    .A3(_09202_),
    .A4(_09315_),
    .ZN(_09747_));
 OR4_X1 _35472_ (.A1(_00444_),
    .A2(_09144_),
    .A3(_09084_),
    .A4(_09099_),
    .ZN(_09748_));
 AND3_X2 _35473_ (.A1(_09746_),
    .A2(_09747_),
    .A3(_09748_),
    .ZN(_09749_));
 OR2_X2 _35474_ (.A1(_09152_),
    .A2(_00443_),
    .ZN(_09750_));
 OR4_X4 _35475_ (.A1(_00442_),
    .A2(_09145_),
    .A3(_09210_),
    .A4(_09080_),
    .ZN(_09751_));
 NAND3_X4 _35476_ (.A1(_09749_),
    .A2(_09750_),
    .A3(_09751_),
    .ZN(_09752_));
 OAI211_X4 _35477_ (.A(_09177_),
    .B(_09742_),
    .C1(_09752_),
    .C2(_09056_),
    .ZN(_09753_));
 NOR2_X1 _35478_ (.A1(_09571_),
    .A2(_00440_),
    .ZN(_09754_));
 NOR2_X1 _35479_ (.A1(_09754_),
    .A2(_09038_),
    .ZN(_09755_));
 NAND3_X1 _35480_ (.A1(_09065_),
    .A2(\icache.data_set_select_mux.data_i [469]),
    .A3(_09130_),
    .ZN(_09756_));
 OAI21_X2 _35481_ (.A(_09756_),
    .B1(_09076_),
    .B2(_00439_),
    .ZN(_09757_));
 NOR4_X2 _35482_ (.A1(_09136_),
    .A2(_09097_),
    .A3(_09312_),
    .A4(_00438_),
    .ZN(_09758_));
 NOR4_X2 _35483_ (.A1(_09123_),
    .A2(_09090_),
    .A3(_09092_),
    .A4(_00437_),
    .ZN(_09759_));
 NOR3_X4 _35484_ (.A1(_09757_),
    .A2(_09758_),
    .A3(_09759_),
    .ZN(_09760_));
 OR4_X1 _35485_ (.A1(_00436_),
    .A2(_09130_),
    .A3(_09231_),
    .A4(_09100_),
    .ZN(_09761_));
 OR2_X1 _35486_ (.A1(_09105_),
    .A2(_00435_),
    .ZN(_09762_));
 NAND3_X2 _35487_ (.A1(_09760_),
    .A2(_09761_),
    .A3(_09762_),
    .ZN(_09763_));
 NOR4_X4 _35488_ (.A1(_09354_),
    .A2(_09098_),
    .A3(_00434_),
    .A4(_09207_),
    .ZN(_09764_));
 NOR4_X1 _35489_ (.A1(_09070_),
    .A2(_09124_),
    .A3(_09334_),
    .A4(_00433_),
    .ZN(_09765_));
 NOR3_X1 _35490_ (.A1(_09763_),
    .A2(_09764_),
    .A3(_09765_),
    .ZN(_09766_));
 MUX2_X1 _35491_ (.A(_00432_),
    .B(_09766_),
    .S(_09571_),
    .Z(_09767_));
 AOI221_X4 _35492_ (.A(_08644_),
    .B1(_09753_),
    .B2(_09755_),
    .C1(_09767_),
    .C2(_09262_),
    .ZN(fe_queue_o[49]));
 AND3_X1 _35493_ (.A1(_09197_),
    .A2(\icache.data_set_select_mux.data_i [470]),
    .A3(_09385_),
    .ZN(_09768_));
 NOR4_X2 _35494_ (.A1(_09332_),
    .A2(_09432_),
    .A3(_09313_),
    .A4(_00454_),
    .ZN(_09769_));
 NOR4_X1 _35495_ (.A1(_09140_),
    .A2(_09316_),
    .A3(_00455_),
    .A4(_09149_),
    .ZN(_09770_));
 NOR3_X2 _35496_ (.A1(_09768_),
    .A2(_09769_),
    .A3(_09770_),
    .ZN(_09771_));
 NOR2_X2 _35497_ (.A1(_09436_),
    .A2(_00451_),
    .ZN(_09772_));
 NOR2_X2 _35498_ (.A1(_09772_),
    .A2(_09214_),
    .ZN(_09773_));
 OR4_X2 _35499_ (.A1(_00453_),
    .A2(_09238_),
    .A3(_09109_),
    .A4(_09208_),
    .ZN(_09774_));
 OR4_X1 _35500_ (.A1(_00452_),
    .A2(_09145_),
    .A3(_09210_),
    .A4(_09211_),
    .ZN(_09775_));
 AND4_X1 _35501_ (.A1(_09771_),
    .A2(_09773_),
    .A3(_09774_),
    .A4(_09775_),
    .ZN(_09776_));
 AND4_X1 _35502_ (.A1(_00450_),
    .A2(_09358_),
    .A3(_09114_),
    .A4(_09150_),
    .ZN(_09777_));
 OAI221_X2 _35503_ (.A(_09194_),
    .B1(_00449_),
    .B2(_09057_),
    .C1(_09776_),
    .C2(_09777_),
    .ZN(_09778_));
 NAND2_X2 _35504_ (.A1(net1264),
    .A2(_00448_),
    .ZN(_09779_));
 AOI21_X4 _35505_ (.A(_09587_),
    .B1(_09778_),
    .B2(_09779_),
    .ZN(_09780_));
 NOR2_X1 _35506_ (.A1(_09074_),
    .A2(_00463_),
    .ZN(_09781_));
 AND3_X1 _35507_ (.A1(_09063_),
    .A2(\icache.data_set_select_mux.data_i [502]),
    .A3(_09067_),
    .ZN(_09782_));
 NOR4_X1 _35508_ (.A1(_09045_),
    .A2(_09083_),
    .A3(_09053_),
    .A4(_00462_),
    .ZN(_09783_));
 NOR3_X1 _35509_ (.A1(_09781_),
    .A2(_09782_),
    .A3(_09783_),
    .ZN(_09784_));
 OR4_X2 _35510_ (.A1(_00461_),
    .A2(_09045_),
    .A3(_09053_),
    .A4(_09047_),
    .ZN(_09785_));
 OR4_X1 _35511_ (.A1(_00460_),
    .A2(_09067_),
    .A3(_09083_),
    .A4(_09043_),
    .ZN(_09786_));
 AND3_X1 _35512_ (.A1(_09784_),
    .A2(_09785_),
    .A3(_09786_),
    .ZN(_09787_));
 MUX2_X1 _35513_ (.A(_00459_),
    .B(_09787_),
    .S(_09105_),
    .Z(_09788_));
 MUX2_X2 _35514_ (.A(_00458_),
    .B(_09788_),
    .S(_09061_),
    .Z(_09789_));
 OR4_X1 _35515_ (.A1(_00457_),
    .A2(_09354_),
    .A3(_09081_),
    .A4(_09113_),
    .ZN(_09790_));
 AND2_X2 _35516_ (.A1(_09789_),
    .A2(_09790_),
    .ZN(_09791_));
 MUX2_X1 _35517_ (.A(_00456_),
    .B(_09791_),
    .S(_09178_),
    .Z(_09792_));
 AOI211_X2 _35518_ (.A(_09688_),
    .B(_09780_),
    .C1(_09792_),
    .C2(_09308_),
    .ZN(fe_queue_o[50]));
 AND3_X1 _35519_ (.A1(_09059_),
    .A2(_00474_),
    .A3(_09091_),
    .ZN(_09793_));
 NOR2_X1 _35520_ (.A1(_09075_),
    .A2(_00479_),
    .ZN(_09794_));
 AND3_X1 _35521_ (.A1(_09128_),
    .A2(\icache.data_set_select_mux.data_i [503]),
    .A3(_09144_),
    .ZN(_09795_));
 NOR4_X1 _35522_ (.A1(_09254_),
    .A2(_09200_),
    .A3(_09497_),
    .A4(_00478_),
    .ZN(_09796_));
 NOR3_X1 _35523_ (.A1(_09794_),
    .A2(_09795_),
    .A3(_09796_),
    .ZN(_09797_));
 OR4_X1 _35524_ (.A1(_00477_),
    .A2(_09206_),
    .A3(_09202_),
    .A4(_09315_),
    .ZN(_09798_));
 OR4_X1 _35525_ (.A1(_00476_),
    .A2(_09378_),
    .A3(_09200_),
    .A4(_09099_),
    .ZN(_09799_));
 AND3_X1 _35526_ (.A1(_09797_),
    .A2(_09798_),
    .A3(_09799_),
    .ZN(_09800_));
 NOR4_X1 _35527_ (.A1(_09131_),
    .A2(_00475_),
    .A3(_09316_),
    .A4(_09149_),
    .ZN(_09801_));
 NOR2_X1 _35528_ (.A1(_09214_),
    .A2(_09801_),
    .ZN(_09802_));
 AOI21_X4 _35529_ (.A(_09793_),
    .B1(_09800_),
    .B2(_09802_),
    .ZN(_09803_));
 NOR4_X1 _35530_ (.A1(_09122_),
    .A2(_09258_),
    .A3(_09343_),
    .A4(_00473_),
    .ZN(_09804_));
 OAI21_X2 _35531_ (.A(_09041_),
    .B1(_09803_),
    .B2(_09804_),
    .ZN(_09805_));
 NOR2_X1 _35532_ (.A1(_09040_),
    .A2(_00472_),
    .ZN(_09806_));
 NOR2_X1 _35533_ (.A1(_09806_),
    .A2(_09038_),
    .ZN(_09807_));
 NAND3_X2 _35534_ (.A1(_09065_),
    .A2(\icache.data_set_select_mux.data_i [471]),
    .A3(_09130_),
    .ZN(_09808_));
 OAI21_X4 _35535_ (.A(_09808_),
    .B1(_09076_),
    .B2(_00471_),
    .ZN(_09809_));
 NOR4_X2 _35536_ (.A1(_09123_),
    .A2(_09097_),
    .A3(_09312_),
    .A4(_00470_),
    .ZN(_09810_));
 NOR4_X2 _35537_ (.A1(_09123_),
    .A2(_09312_),
    .A3(_09315_),
    .A4(_00469_),
    .ZN(_09811_));
 NOR3_X4 _35538_ (.A1(_09809_),
    .A2(_09810_),
    .A3(_09811_),
    .ZN(_09812_));
 OR4_X1 _35539_ (.A1(_00468_),
    .A2(_09130_),
    .A3(_09231_),
    .A4(_09100_),
    .ZN(_09813_));
 OR2_X1 _35540_ (.A1(_09105_),
    .A2(_00467_),
    .ZN(_09814_));
 NAND3_X2 _35541_ (.A1(_09812_),
    .A2(_09813_),
    .A3(_09814_),
    .ZN(_09815_));
 NOR4_X4 _35542_ (.A1(_09354_),
    .A2(_09098_),
    .A3(_00466_),
    .A4(_09207_),
    .ZN(_09816_));
 NOR4_X1 _35543_ (.A1(_09070_),
    .A2(_09124_),
    .A3(_09334_),
    .A4(_00465_),
    .ZN(_09817_));
 NOR3_X1 _35544_ (.A1(_09815_),
    .A2(_09816_),
    .A3(_09817_),
    .ZN(_09818_));
 MUX2_X1 _35545_ (.A(_00464_),
    .B(_09818_),
    .S(_09571_),
    .Z(_09819_));
 AOI221_X4 _35546_ (.A(_08644_),
    .B1(_09805_),
    .B2(_09807_),
    .C1(_09819_),
    .C2(_09262_),
    .ZN(fe_queue_o[51]));
 NOR2_X2 _35547_ (.A1(_09195_),
    .A2(_00487_),
    .ZN(_09820_));
 AND3_X1 _35548_ (.A1(_09197_),
    .A2(\icache.data_set_select_mux.data_i [472]),
    .A3(_09198_),
    .ZN(_09821_));
 NOR4_X2 _35549_ (.A1(_09124_),
    .A2(_09201_),
    .A3(_09203_),
    .A4(_00486_),
    .ZN(_09822_));
 NOR3_X4 _35550_ (.A1(_09820_),
    .A2(_09821_),
    .A3(_09822_),
    .ZN(_09823_));
 OR4_X4 _35551_ (.A1(_00485_),
    .A2(_09207_),
    .A3(_09203_),
    .A4(_09208_),
    .ZN(_09824_));
 OR4_X1 _35552_ (.A1(_00484_),
    .A2(_09198_),
    .A3(_09210_),
    .A4(_09211_),
    .ZN(_09825_));
 NOR2_X2 _35553_ (.A1(_09152_),
    .A2(_00483_),
    .ZN(_09826_));
 NOR2_X4 _35554_ (.A1(_09826_),
    .A2(_09060_),
    .ZN(_09827_));
 AND4_X2 _35555_ (.A1(_09823_),
    .A2(_09824_),
    .A3(_09825_),
    .A4(_09827_),
    .ZN(_09828_));
 AND4_X1 _35556_ (.A1(_00482_),
    .A2(_09358_),
    .A3(_09126_),
    .A4(_09150_),
    .ZN(_09829_));
 OAI221_X2 _35557_ (.A(_09245_),
    .B1(_00481_),
    .B2(_09057_),
    .C1(_09828_),
    .C2(_09829_),
    .ZN(_09830_));
 NAND2_X2 _35558_ (.A1(net1264),
    .A2(_00480_),
    .ZN(_09831_));
 AOI21_X2 _35559_ (.A(_09587_),
    .B1(_09830_),
    .B2(_09831_),
    .ZN(_09832_));
 NOR2_X1 _35560_ (.A1(_09162_),
    .A2(_00493_),
    .ZN(_09833_));
 NAND3_X1 _35561_ (.A1(_09129_),
    .A2(\icache.data_set_select_mux.data_i [504]),
    .A3(_09385_),
    .ZN(_09834_));
 OAI21_X2 _35562_ (.A(_09834_),
    .B1(_09195_),
    .B2(_00495_),
    .ZN(_09835_));
 NOR4_X2 _35563_ (.A1(_09227_),
    .A2(_09098_),
    .A3(_09138_),
    .A4(_00494_),
    .ZN(_09836_));
 NOR3_X4 _35564_ (.A1(_09833_),
    .A2(_09835_),
    .A3(_09836_),
    .ZN(_09837_));
 OR4_X2 _35565_ (.A1(_00492_),
    .A2(_09271_),
    .A3(_09432_),
    .A4(_09272_),
    .ZN(_09838_));
 OR2_X2 _35566_ (.A1(_09436_),
    .A2(_00491_),
    .ZN(_09839_));
 NAND3_X4 _35567_ (.A1(_09837_),
    .A2(_09838_),
    .A3(_09839_),
    .ZN(_09840_));
 NOR4_X2 _35568_ (.A1(_09276_),
    .A2(_09426_),
    .A3(_00490_),
    .A4(_09341_),
    .ZN(_09841_));
 NOR4_X2 _35569_ (.A1(_09237_),
    .A2(_09240_),
    .A3(_09241_),
    .A4(_00489_),
    .ZN(_09842_));
 NOR3_X4 _35570_ (.A1(_09840_),
    .A2(_09841_),
    .A3(_09842_),
    .ZN(_09843_));
 MUX2_X1 _35571_ (.A(_00488_),
    .B(_09843_),
    .S(_09280_),
    .Z(_09844_));
 AOI211_X2 _35572_ (.A(_09688_),
    .B(_09832_),
    .C1(_09223_),
    .C2(_09844_),
    .ZN(fe_queue_o[52]));
 NAND3_X1 _35573_ (.A1(_09129_),
    .A2(\icache.data_set_select_mux.data_i [473]),
    .A3(_09385_),
    .ZN(_09845_));
 OAI21_X2 _35574_ (.A(_09845_),
    .B1(_09195_),
    .B2(_00503_),
    .ZN(_09846_));
 NOR4_X2 _35575_ (.A1(_09255_),
    .A2(_09201_),
    .A3(_09203_),
    .A4(_00502_),
    .ZN(_09847_));
 NOR4_X2 _35576_ (.A1(_09255_),
    .A2(_09313_),
    .A3(_09208_),
    .A4(_00501_),
    .ZN(_09848_));
 NOR4_X4 _35577_ (.A1(_09846_),
    .A2(_09311_),
    .A3(_09847_),
    .A4(_09848_),
    .ZN(_09849_));
 AND4_X1 _35578_ (.A1(_00500_),
    .A2(_09258_),
    .A3(_09113_),
    .A4(_09110_),
    .ZN(_09850_));
 OAI221_X2 _35579_ (.A(_09062_),
    .B1(_00499_),
    .B2(_09153_),
    .C1(_09849_),
    .C2(_09850_),
    .ZN(_09851_));
 NAND4_X4 _35580_ (.A1(_09111_),
    .A2(_09114_),
    .A3(_00498_),
    .A4(_09115_),
    .ZN(_09852_));
 AOI21_X4 _35581_ (.A(_09056_),
    .B1(_09851_),
    .B2(_09852_),
    .ZN(_09853_));
 AND3_X1 _35582_ (.A1(_09323_),
    .A2(_00497_),
    .A3(_09111_),
    .ZN(_09854_));
 NOR3_X2 _35583_ (.A1(_09853_),
    .A2(_09220_),
    .A3(_09854_),
    .ZN(_09855_));
 NOR2_X1 _35584_ (.A1(_09042_),
    .A2(_00496_),
    .ZN(_09856_));
 NOR3_X4 _35585_ (.A1(_09855_),
    .A2(_09121_),
    .A3(_09856_),
    .ZN(_09857_));
 NAND4_X2 _35586_ (.A1(_09148_),
    .A2(_00507_),
    .A3(_09259_),
    .A4(_09172_),
    .ZN(_09858_));
 NAND3_X2 _35587_ (.A1(_09129_),
    .A2(\icache.data_set_select_mux.data_i [505]),
    .A3(_09131_),
    .ZN(_09859_));
 OAI21_X4 _35588_ (.A(_09859_),
    .B1(_09133_),
    .B2(_00511_),
    .ZN(_09860_));
 NOR4_X2 _35589_ (.A1(_09086_),
    .A2(_09332_),
    .A3(_09138_),
    .A4(_00510_),
    .ZN(_09861_));
 NOR4_X2 _35590_ (.A1(_09137_),
    .A2(_09140_),
    .A3(_09334_),
    .A4(_00509_),
    .ZN(_09862_));
 NOR3_X4 _35591_ (.A1(_09860_),
    .A2(_09861_),
    .A3(_09862_),
    .ZN(_09863_));
 OAI21_X2 _35592_ (.A(_09863_),
    .B1(_00508_),
    .B2(_09337_),
    .ZN(_09864_));
 OAI21_X4 _35593_ (.A(_09858_),
    .B1(_09864_),
    .B2(_09103_),
    .ZN(_09865_));
 OR4_X2 _35594_ (.A1(_00506_),
    .A2(_09340_),
    .A3(_09135_),
    .A4(_09341_),
    .ZN(_09866_));
 OR4_X2 _35595_ (.A1(_00505_),
    .A2(_09340_),
    .A3(_09341_),
    .A4(_09343_),
    .ZN(_09867_));
 NAND4_X4 _35596_ (.A1(_09865_),
    .A2(_09178_),
    .A3(_09866_),
    .A4(_09867_),
    .ZN(_09868_));
 NAND2_X1 _35597_ (.A1(_09118_),
    .A2(_00504_),
    .ZN(_09869_));
 AOI21_X2 _35598_ (.A(_09039_),
    .B1(_09868_),
    .B2(_09869_),
    .ZN(_09870_));
 NOR3_X4 _35599_ (.A1(_09857_),
    .A2(fe_queue_o[99]),
    .A3(_09870_),
    .ZN(fe_queue_o[53]));
 AND3_X1 _35600_ (.A1(_09197_),
    .A2(\icache.data_set_select_mux.data_i [474]),
    .A3(_09385_),
    .ZN(_09871_));
 NOR4_X2 _35601_ (.A1(_09332_),
    .A2(_09201_),
    .A3(_09313_),
    .A4(_00518_),
    .ZN(_09872_));
 NOR4_X1 _35602_ (.A1(_09140_),
    .A2(_09316_),
    .A3(_00519_),
    .A4(_09211_),
    .ZN(_09873_));
 NOR3_X2 _35603_ (.A1(_09871_),
    .A2(_09872_),
    .A3(_09873_),
    .ZN(_09874_));
 NOR2_X4 _35604_ (.A1(_09436_),
    .A2(_00515_),
    .ZN(_09875_));
 NOR2_X2 _35605_ (.A1(_09875_),
    .A2(_09214_),
    .ZN(_09876_));
 OR4_X2 _35606_ (.A1(_00517_),
    .A2(_09238_),
    .A3(_09109_),
    .A4(_09208_),
    .ZN(_09877_));
 OR4_X1 _35607_ (.A1(_00516_),
    .A2(_09145_),
    .A3(_09210_),
    .A4(_09211_),
    .ZN(_09878_));
 AND4_X2 _35608_ (.A1(_09874_),
    .A2(_09876_),
    .A3(_09877_),
    .A4(_09878_),
    .ZN(_09879_));
 AND4_X1 _35609_ (.A1(_00514_),
    .A2(_09358_),
    .A3(_09126_),
    .A4(_09150_),
    .ZN(_09880_));
 OAI221_X2 _35610_ (.A(_09245_),
    .B1(_00513_),
    .B2(_09057_),
    .C1(_09879_),
    .C2(_09880_),
    .ZN(_09881_));
 NAND2_X2 _35611_ (.A1(net1264),
    .A2(_00512_),
    .ZN(_09882_));
 AOI21_X1 _35612_ (.A(_09587_),
    .B1(_09881_),
    .B2(_09882_),
    .ZN(_09883_));
 NAND3_X2 _35613_ (.A1(_09329_),
    .A2(\icache.data_set_select_mux.data_i [506]),
    .A3(_09230_),
    .ZN(_09884_));
 OAI21_X4 _35614_ (.A(_09884_),
    .B1(_09133_),
    .B2(_00527_),
    .ZN(_09885_));
 NOR4_X2 _35615_ (.A1(_09239_),
    .A2(_09267_),
    .A3(_09166_),
    .A4(_00526_),
    .ZN(_09886_));
 NOR4_X2 _35616_ (.A1(_09227_),
    .A2(_09088_),
    .A3(_09141_),
    .A4(_00525_),
    .ZN(_09887_));
 NOR3_X4 _35617_ (.A1(_09885_),
    .A2(_09886_),
    .A3(_09887_),
    .ZN(_09888_));
 OR4_X2 _35618_ (.A1(_00524_),
    .A2(_09271_),
    .A3(_09432_),
    .A4(_09272_),
    .ZN(_09889_));
 OR2_X1 _35619_ (.A1(_09436_),
    .A2(_00523_),
    .ZN(_09890_));
 NAND3_X4 _35620_ (.A1(_09888_),
    .A2(_09889_),
    .A3(_09890_),
    .ZN(_09891_));
 NOR4_X2 _35621_ (.A1(_09276_),
    .A2(_09426_),
    .A3(_00522_),
    .A4(_09341_),
    .ZN(_09892_));
 NOR4_X2 _35622_ (.A1(_09122_),
    .A2(_09240_),
    .A3(_09241_),
    .A4(_00521_),
    .ZN(_09893_));
 NOR3_X4 _35623_ (.A1(_09891_),
    .A2(_09892_),
    .A3(_09893_),
    .ZN(_09894_));
 MUX2_X1 _35624_ (.A(_00520_),
    .B(_09894_),
    .S(_09280_),
    .Z(_09895_));
 AOI211_X2 _35625_ (.A(_09688_),
    .B(_09883_),
    .C1(_09223_),
    .C2(_09895_),
    .ZN(fe_queue_o[54]));
 NAND3_X1 _35626_ (.A1(_09323_),
    .A2(_00529_),
    .A3(_09217_),
    .ZN(_09896_));
 NOR2_X1 _35627_ (.A1(_09075_),
    .A2(_00535_),
    .ZN(_09897_));
 AND3_X1 _35628_ (.A1(_09064_),
    .A2(\icache.data_set_select_mux.data_i [475]),
    .A3(_09144_),
    .ZN(_09898_));
 NOR4_X1 _35629_ (.A1(_09254_),
    .A2(_09200_),
    .A3(_09497_),
    .A4(_00534_),
    .ZN(_09899_));
 NOR3_X1 _35630_ (.A1(_09897_),
    .A2(_09898_),
    .A3(_09899_),
    .ZN(_09900_));
 OR4_X1 _35631_ (.A1(_00533_),
    .A2(_09206_),
    .A3(_09202_),
    .A4(_09315_),
    .ZN(_09901_));
 OR4_X1 _35632_ (.A1(_00532_),
    .A2(_09144_),
    .A3(_09084_),
    .A4(_09099_),
    .ZN(_09902_));
 AND3_X1 _35633_ (.A1(_09900_),
    .A2(_09901_),
    .A3(_09902_),
    .ZN(_09903_));
 OR2_X2 _35634_ (.A1(_09152_),
    .A2(_00531_),
    .ZN(_09904_));
 OR4_X4 _35635_ (.A1(_00530_),
    .A2(_09145_),
    .A3(_09085_),
    .A4(_09080_),
    .ZN(_09905_));
 NAND3_X4 _35636_ (.A1(_09903_),
    .A2(_09904_),
    .A3(_09905_),
    .ZN(_09906_));
 OAI211_X1 _35637_ (.A(_09177_),
    .B(_09896_),
    .C1(_09906_),
    .C2(_09056_),
    .ZN(_09907_));
 NOR2_X1 _35638_ (.A1(_09040_),
    .A2(_00528_),
    .ZN(_09908_));
 NOR2_X1 _35639_ (.A1(_09908_),
    .A2(net1389),
    .ZN(_09909_));
 NAND3_X1 _35640_ (.A1(_09128_),
    .A2(\icache.data_set_select_mux.data_i [507]),
    .A3(_09130_),
    .ZN(_09910_));
 OAI21_X2 _35641_ (.A(_09910_),
    .B1(_09076_),
    .B2(_00543_),
    .ZN(_09911_));
 NOR4_X2 _35642_ (.A1(_09123_),
    .A2(_09097_),
    .A3(_09312_),
    .A4(_00542_),
    .ZN(_09912_));
 NOR4_X2 _35643_ (.A1(_09123_),
    .A2(_09312_),
    .A3(_09315_),
    .A4(_00541_),
    .ZN(_09913_));
 NOR3_X4 _35644_ (.A1(_09911_),
    .A2(_09912_),
    .A3(_09913_),
    .ZN(_09914_));
 OR4_X1 _35645_ (.A1(_00540_),
    .A2(_09130_),
    .A3(_09231_),
    .A4(_09100_),
    .ZN(_09915_));
 OR2_X2 _35646_ (.A1(_09105_),
    .A2(_00539_),
    .ZN(_09916_));
 NAND3_X2 _35647_ (.A1(_09914_),
    .A2(_09915_),
    .A3(_09916_),
    .ZN(_09917_));
 NOR4_X4 _35648_ (.A1(_09354_),
    .A2(_09098_),
    .A3(_00538_),
    .A4(_09207_),
    .ZN(_09918_));
 NOR4_X1 _35649_ (.A1(_09070_),
    .A2(_09124_),
    .A3(_09334_),
    .A4(_00537_),
    .ZN(_09919_));
 NOR3_X1 _35650_ (.A1(_09917_),
    .A2(_09918_),
    .A3(_09919_),
    .ZN(_09920_));
 MUX2_X1 _35651_ (.A(_00536_),
    .B(_09920_),
    .S(_09571_),
    .Z(_09921_));
 AOI221_X4 _35652_ (.A(_08643_),
    .B1(_09907_),
    .B2(_09909_),
    .C1(_09921_),
    .C2(_09587_),
    .ZN(fe_queue_o[55]));
 NAND3_X2 _35653_ (.A1(_09066_),
    .A2(\icache.data_set_select_mux.data_i [508]),
    .A3(_09070_),
    .ZN(_09922_));
 OAI21_X4 _35654_ (.A(_09922_),
    .B1(_09077_),
    .B2(_00559_),
    .ZN(_09923_));
 NOR4_X1 _35655_ (.A1(_09135_),
    .A2(_09137_),
    .A3(_09091_),
    .A4(_00558_),
    .ZN(_09924_));
 NOR4_X2 _35656_ (.A1(_09081_),
    .A2(_09091_),
    .A3(_09093_),
    .A4(_00557_),
    .ZN(_09925_));
 OR3_X4 _35657_ (.A1(_09923_),
    .A2(_09924_),
    .A3(_09925_),
    .ZN(_09926_));
 NOR4_X4 _35658_ (.A1(_09147_),
    .A2(_09148_),
    .A3(_00556_),
    .A4(_09150_),
    .ZN(_09927_));
 OAI21_X2 _35659_ (.A(_09062_),
    .B1(_09153_),
    .B2(_00555_),
    .ZN(_09928_));
 NOR3_X4 _35660_ (.A1(_09926_),
    .A2(_09927_),
    .A3(_09928_),
    .ZN(_09929_));
 AND3_X1 _35661_ (.A1(_09156_),
    .A2(_00554_),
    .A3(_09111_),
    .ZN(_09930_));
 OAI221_X2 _35662_ (.A(_09042_),
    .B1(_00553_),
    .B2(_09058_),
    .C1(_09929_),
    .C2(_09930_),
    .ZN(_09931_));
 NAND2_X1 _35663_ (.A1(_09118_),
    .A2(_00552_),
    .ZN(_09932_));
 AOI21_X2 _35664_ (.A(_09039_),
    .B1(_09931_),
    .B2(_09932_),
    .ZN(_09933_));
 AND3_X1 _35665_ (.A1(_09197_),
    .A2(\icache.data_set_select_mux.data_i [476]),
    .A3(_09145_),
    .ZN(_09934_));
 NOR4_X2 _35666_ (.A1(_09201_),
    .A2(_09136_),
    .A3(_09087_),
    .A4(_00550_),
    .ZN(_09935_));
 NOR4_X1 _35667_ (.A1(_09109_),
    .A2(_09112_),
    .A3(_00551_),
    .A4(_09186_),
    .ZN(_09936_));
 OR3_X2 _35668_ (.A1(_09934_),
    .A2(_09935_),
    .A3(_09936_),
    .ZN(_09937_));
 NOR4_X1 _35669_ (.A1(_09258_),
    .A2(_09110_),
    .A3(_09113_),
    .A4(_00549_),
    .ZN(_09938_));
 NOR4_X1 _35670_ (.A1(_09146_),
    .A2(_09135_),
    .A3(_00548_),
    .A4(_09101_),
    .ZN(_09939_));
 NOR3_X2 _35671_ (.A1(_09937_),
    .A2(_09938_),
    .A3(_09939_),
    .ZN(_09940_));
 OR4_X2 _35672_ (.A1(_00547_),
    .A2(_09354_),
    .A3(_09101_),
    .A4(_09113_),
    .ZN(_09941_));
 INV_X4 _35673_ (.A(_00546_),
    .ZN(_09942_));
 OAI211_X4 _35674_ (.A(_09115_),
    .B(_09217_),
    .C1(_09148_),
    .C2(_09942_),
    .ZN(_09943_));
 NAND3_X4 _35675_ (.A1(_09940_),
    .A2(_09941_),
    .A3(_09943_),
    .ZN(_09944_));
 NAND3_X1 _35676_ (.A1(_09323_),
    .A2(_00545_),
    .A3(_09111_),
    .ZN(_09945_));
 NAND3_X2 _35677_ (.A1(_09944_),
    .A2(_09194_),
    .A3(_09945_),
    .ZN(_09946_));
 OR2_X1 _35678_ (.A1(_09041_),
    .A2(_00544_),
    .ZN(_09947_));
 AND3_X1 _35679_ (.A1(_09946_),
    .A2(_09039_),
    .A3(_09947_),
    .ZN(_09948_));
 NOR3_X4 _35680_ (.A1(_09933_),
    .A2(fe_queue_o[99]),
    .A3(_09948_),
    .ZN(fe_queue_o[56]));
 AND3_X1 _35681_ (.A1(_09197_),
    .A2(\icache.data_set_select_mux.data_i [477]),
    .A3(_09385_),
    .ZN(_09949_));
 NOR4_X2 _35682_ (.A1(_09332_),
    .A2(_09201_),
    .A3(_09313_),
    .A4(_00566_),
    .ZN(_09950_));
 NOR4_X1 _35683_ (.A1(_09140_),
    .A2(_09316_),
    .A3(_00567_),
    .A4(_09211_),
    .ZN(_09951_));
 NOR3_X2 _35684_ (.A1(_09949_),
    .A2(_09950_),
    .A3(_09951_),
    .ZN(_09952_));
 NOR2_X2 _35685_ (.A1(_09436_),
    .A2(_00563_),
    .ZN(_09953_));
 NOR2_X1 _35686_ (.A1(_09953_),
    .A2(_09214_),
    .ZN(_09954_));
 OR4_X4 _35687_ (.A1(_00565_),
    .A2(_09238_),
    .A3(_09109_),
    .A4(_09208_),
    .ZN(_09955_));
 OR4_X1 _35688_ (.A1(_00564_),
    .A2(_09145_),
    .A3(_09210_),
    .A4(_09211_),
    .ZN(_09956_));
 AND4_X2 _35689_ (.A1(_09952_),
    .A2(_09954_),
    .A3(_09955_),
    .A4(_09956_),
    .ZN(_09957_));
 AND4_X1 _35690_ (.A1(_00562_),
    .A2(_09358_),
    .A3(_09126_),
    .A4(_09150_),
    .ZN(_09958_));
 OAI221_X2 _35691_ (.A(_09245_),
    .B1(_00561_),
    .B2(_09057_),
    .C1(_09957_),
    .C2(_09958_),
    .ZN(_09959_));
 NAND2_X2 _35692_ (.A1(net1264),
    .A2(_00560_),
    .ZN(_09960_));
 AOI21_X1 _35693_ (.A(_09587_),
    .B1(_09959_),
    .B2(_09960_),
    .ZN(_09961_));
 NAND3_X1 _35694_ (.A1(_09329_),
    .A2(\icache.data_set_select_mux.data_i [509]),
    .A3(_09230_),
    .ZN(_09962_));
 OAI21_X1 _35695_ (.A(_09962_),
    .B1(_09133_),
    .B2(_00575_),
    .ZN(_09963_));
 NOR4_X4 _35696_ (.A1(_09239_),
    .A2(_09267_),
    .A3(_09138_),
    .A4(_00574_),
    .ZN(_09964_));
 NOR4_X4 _35697_ (.A1(_09137_),
    .A2(_09088_),
    .A3(_09141_),
    .A4(_00573_),
    .ZN(_09965_));
 NOR3_X2 _35698_ (.A1(_09963_),
    .A2(_09964_),
    .A3(_09965_),
    .ZN(_09966_));
 OR4_X2 _35699_ (.A1(_00572_),
    .A2(_09271_),
    .A3(_09432_),
    .A4(_09272_),
    .ZN(_09967_));
 OR2_X2 _35700_ (.A1(_09436_),
    .A2(_00571_),
    .ZN(_09968_));
 NAND3_X4 _35701_ (.A1(_09966_),
    .A2(_09967_),
    .A3(_09968_),
    .ZN(_09969_));
 NOR4_X1 _35702_ (.A1(_09276_),
    .A2(_09426_),
    .A3(_00570_),
    .A4(_09341_),
    .ZN(_09970_));
 NOR4_X1 _35703_ (.A1(_09122_),
    .A2(_09125_),
    .A3(_09343_),
    .A4(_00569_),
    .ZN(_09971_));
 NOR3_X2 _35704_ (.A1(_09969_),
    .A2(_09970_),
    .A3(_09971_),
    .ZN(_09972_));
 MUX2_X1 _35705_ (.A(_00568_),
    .B(_09972_),
    .S(_09280_),
    .Z(_09973_));
 AOI211_X2 _35706_ (.A(_09688_),
    .B(_09961_),
    .C1(_09308_),
    .C2(_09973_),
    .ZN(fe_queue_o[57]));
 AND3_X1 _35707_ (.A1(_09059_),
    .A2(\icache.data_set_select_mux.data_i [382]),
    .A3(_09070_),
    .ZN(_09974_));
 AOI21_X4 _35708_ (.A(_09974_),
    .B1(\icache.data_set_select_mux.data_i [446]),
    .B2(_09073_),
    .ZN(_09975_));
 NAND3_X2 _35709_ (.A1(_09156_),
    .A2(\icache.data_set_select_mux.data_i [126]),
    .A3(_09217_),
    .ZN(_09976_));
 NAND3_X2 _35710_ (.A1(_09323_),
    .A2(\icache.data_set_select_mux.data_i [318]),
    .A3(_09237_),
    .ZN(_09977_));
 NAND3_X4 _35711_ (.A1(_09975_),
    .A2(_09976_),
    .A3(_09977_),
    .ZN(_09978_));
 NAND3_X1 _35712_ (.A1(_09066_),
    .A2(\icache.data_set_select_mux.data_i [254]),
    .A3(_09358_),
    .ZN(_09979_));
 NAND3_X1 _35713_ (.A1(_09066_),
    .A2(\icache.data_set_select_mux.data_i [510]),
    .A3(_09122_),
    .ZN(_09980_));
 NAND3_X2 _35714_ (.A1(_09323_),
    .A2(\icache.data_set_select_mux.data_i [62]),
    .A3(_09358_),
    .ZN(_09981_));
 NAND3_X1 _35715_ (.A1(_09072_),
    .A2(\icache.data_set_select_mux.data_i [190]),
    .A3(_09358_),
    .ZN(_09982_));
 NAND4_X1 _35716_ (.A1(_09979_),
    .A2(_09980_),
    .A3(_09981_),
    .A4(_09982_),
    .ZN(_09983_));
 OAI21_X1 _35717_ (.A(net1389),
    .B1(_09978_),
    .B2(_09983_),
    .ZN(_09984_));
 NAND3_X1 _35718_ (.A1(_09066_),
    .A2(\icache.data_set_select_mux.data_i [222]),
    .A3(_09217_),
    .ZN(_09985_));
 NAND3_X2 _35719_ (.A1(_09156_),
    .A2(net1266),
    .A3(_09358_),
    .ZN(_09986_));
 NAND3_X2 _35720_ (.A1(_09156_),
    .A2(\icache.data_set_select_mux.data_i [350]),
    .A3(_09122_),
    .ZN(_09987_));
 NAND3_X2 _35721_ (.A1(_09323_),
    .A2(\icache.data_set_select_mux.data_i [30]),
    .A3(_09358_),
    .ZN(_09988_));
 NAND4_X4 _35722_ (.A1(_09985_),
    .A2(_09986_),
    .A3(_09987_),
    .A4(_09988_),
    .ZN(_09989_));
 NAND3_X1 _35723_ (.A1(_09066_),
    .A2(\icache.data_set_select_mux.data_i [478]),
    .A3(_09122_),
    .ZN(_09990_));
 NAND3_X1 _35724_ (.A1(_09072_),
    .A2(\icache.data_set_select_mux.data_i [158]),
    .A3(_09110_),
    .ZN(_09991_));
 NAND3_X4 _35725_ (.A1(_09049_),
    .A2(\icache.data_set_select_mux.data_i [286]),
    .A3(_09340_),
    .ZN(_09992_));
 NAND3_X1 _35726_ (.A1(_09072_),
    .A2(\icache.data_set_select_mux.data_i [414]),
    .A3(_09340_),
    .ZN(_09993_));
 NAND4_X2 _35727_ (.A1(_09990_),
    .A2(_09991_),
    .A3(_09992_),
    .A4(_09993_),
    .ZN(_09994_));
 OAI21_X2 _35728_ (.A(_09262_),
    .B1(_09989_),
    .B2(_09994_),
    .ZN(_09995_));
 AOI21_X2 _35729_ (.A(_09220_),
    .B1(_09984_),
    .B2(_09995_),
    .ZN(_09996_));
 MUX2_X2 _35730_ (.A(\icache.final_data_mux.data_i [94]),
    .B(\icache.final_data_mux.data_i [126]),
    .S(net1390),
    .Z(_09997_));
 AND2_X1 _35731_ (.A1(_09997_),
    .A2(net1264),
    .ZN(_09998_));
 OAI21_X4 _35732_ (.A(_08647_),
    .B1(_09996_),
    .B2(_09998_),
    .ZN(_09999_));
 AND3_X1 _35733_ (.A1(_08641_),
    .A2(_08660_),
    .A3(\bp_fe_pc_gen_1.pc_v_if2_r ),
    .ZN(_10000_));
 INV_X1 _35734_ (.A(_10000_),
    .ZN(_10001_));
 OAI21_X4 _35735_ (.A(_09999_),
    .B1(\bp_fe_pc_gen_1.pc_if2_r [1]),
    .B2(_10001_),
    .ZN(fe_queue_o[58]));
 AND3_X1 _35736_ (.A1(_09064_),
    .A2(\icache.data_set_select_mux.data_i [255]),
    .A3(_09497_),
    .ZN(_10002_));
 AND3_X1 _35737_ (.A1(_09072_),
    .A2(\icache.data_set_select_mux.data_i [191]),
    .A3(_09054_),
    .ZN(_10003_));
 OR2_X1 _35738_ (.A1(_10002_),
    .A2(_10003_),
    .ZN(_10004_));
 AOI221_X4 _35739_ (.A(_10004_),
    .B1(\icache.data_set_select_mux.data_i [127]),
    .B2(_09060_),
    .C1(\icache.data_set_select_mux.data_i [63]),
    .C2(_09056_),
    .ZN(_10005_));
 AND3_X1 _35740_ (.A1(_09072_),
    .A2(\icache.data_set_select_mux.data_i [447]),
    .A3(_09069_),
    .ZN(_10006_));
 AOI221_X4 _35741_ (.A(_10006_),
    .B1(_09161_),
    .B2(\icache.data_set_select_mux.data_i [319]),
    .C1(\icache.data_set_select_mux.data_i [511]),
    .C2(_09394_),
    .ZN(_10007_));
 NAND3_X1 _35742_ (.A1(_09156_),
    .A2(\icache.data_set_select_mux.data_i [383]),
    .A3(_09147_),
    .ZN(_10008_));
 NAND4_X4 _35743_ (.A1(_10005_),
    .A2(_10007_),
    .A3(_09245_),
    .A4(_10008_),
    .ZN(_10009_));
 OR2_X1 _35744_ (.A1(_09177_),
    .A2(\icache.final_data_mux.data_i [127]),
    .ZN(_10010_));
 AND3_X1 _35745_ (.A1(_10009_),
    .A2(_09587_),
    .A3(_10010_),
    .ZN(_10011_));
 AND3_X1 _35746_ (.A1(_09072_),
    .A2(\icache.data_set_select_mux.data_i [159]),
    .A3(_09087_),
    .ZN(_10012_));
 AOI221_X4 _35747_ (.A(_10012_),
    .B1(_09056_),
    .B2(\icache.data_set_select_mux.data_i [31]),
    .C1(\icache.data_set_select_mux.data_i [223]),
    .C2(_09311_),
    .ZN(_10013_));
 NAND3_X1 _35748_ (.A1(_09066_),
    .A2(\icache.data_set_select_mux.data_i [479]),
    .A3(_09146_),
    .ZN(_10014_));
 NAND3_X1 _35749_ (.A1(_09072_),
    .A2(\icache.data_set_select_mux.data_i [415]),
    .A3(_09146_),
    .ZN(_10015_));
 NAND3_X4 _35750_ (.A1(_09059_),
    .A2(\icache.data_set_select_mux.data_i [351]),
    .A3(_09146_),
    .ZN(_10016_));
 AND3_X1 _35751_ (.A1(_10014_),
    .A2(_10015_),
    .A3(_10016_),
    .ZN(_10017_));
 AOI22_X4 _35752_ (.A1(_09161_),
    .A2(\icache.data_set_select_mux.data_i [287]),
    .B1(_09214_),
    .B2(net1265),
    .ZN(_10018_));
 NAND4_X4 _35753_ (.A1(_10013_),
    .A2(_09041_),
    .A3(_10017_),
    .A4(_10018_),
    .ZN(_10019_));
 OR2_X1 _35754_ (.A1(_09177_),
    .A2(\icache.final_data_mux.data_i [95]),
    .ZN(_10020_));
 AND3_X1 _35755_ (.A1(_10019_),
    .A2(_09262_),
    .A3(_10020_),
    .ZN(_10021_));
 OAI21_X1 _35756_ (.A(_08647_),
    .B1(_10011_),
    .B2(_10021_),
    .ZN(_10022_));
 NAND3_X4 _35757_ (.A1(_09006_),
    .A2(_09008_),
    .A3(_08640_),
    .ZN(_10023_));
 NAND2_X4 _35758_ (.A1(_10022_),
    .A2(_10023_),
    .ZN(fe_queue_o[59]));
 INV_X1 _35759_ (.A(\bp_fe_pc_gen_1.icache_pc_gen_i [0]),
    .ZN(_10024_));
 AOI21_X4 _35760_ (.A(_10000_),
    .B1(_08647_),
    .B2(_10024_),
    .ZN(fe_queue_o[60]));
 MUX2_X2 _35761_ (.A(\bp_fe_pc_gen_1.icache_pc_gen_i [1]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [1]),
    .S(_09688_),
    .Z(fe_queue_o[61]));
 MUX2_X2 _35762_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [11]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [2]),
    .S(_09688_),
    .Z(fe_queue_o[62]));
 MUX2_X2 _35763_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [12]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [3]),
    .S(_09688_),
    .Z(fe_queue_o[63]));
 MUX2_X2 _35764_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [13]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [4]),
    .S(_09688_),
    .Z(fe_queue_o[64]));
 MUX2_X2 _35765_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [14]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [5]),
    .S(_09688_),
    .Z(fe_queue_o[65]));
 BUF_X8 _35766_ (.A(_08643_),
    .Z(_10025_));
 MUX2_X2 _35767_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [15]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [6]),
    .S(_10025_),
    .Z(fe_queue_o[66]));
 MUX2_X2 _35768_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [16]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [7]),
    .S(_10025_),
    .Z(fe_queue_o[67]));
 MUX2_X2 _35769_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [17]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [8]),
    .S(_10025_),
    .Z(fe_queue_o[68]));
 MUX2_X2 _35770_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [18]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [9]),
    .S(_10025_),
    .Z(fe_queue_o[69]));
 MUX2_X2 _35771_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [19]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [10]),
    .S(_10025_),
    .Z(fe_queue_o[70]));
 MUX2_X2 _35772_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [20]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [11]),
    .S(_10025_),
    .Z(fe_queue_o[71]));
 MUX2_X2 _35773_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [21]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [12]),
    .S(_10025_),
    .Z(fe_queue_o[72]));
 MUX2_X2 _35774_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [22]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [13]),
    .S(_10025_),
    .Z(fe_queue_o[73]));
 MUX2_X2 _35775_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [23]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [14]),
    .S(_10025_),
    .Z(fe_queue_o[74]));
 MUX2_X2 _35776_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [24]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [15]),
    .S(_10025_),
    .Z(fe_queue_o[75]));
 BUF_X8 _35777_ (.A(_08643_),
    .Z(_10026_));
 MUX2_X2 _35778_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [25]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [16]),
    .S(_10026_),
    .Z(fe_queue_o[76]));
 MUX2_X2 _35779_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [26]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [17]),
    .S(_10026_),
    .Z(fe_queue_o[77]));
 MUX2_X2 _35780_ (.A(\bp_fe_pc_gen_1.icache_pc_gen_i [18]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [18]),
    .S(_10026_),
    .Z(fe_queue_o[78]));
 MUX2_X2 _35781_ (.A(\bp_fe_pc_gen_1.icache_pc_gen_i [19]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [19]),
    .S(_10026_),
    .Z(fe_queue_o[79]));
 MUX2_X2 _35782_ (.A(\bp_fe_pc_gen_1.icache_pc_gen_i [20]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [20]),
    .S(_10026_),
    .Z(fe_queue_o[80]));
 MUX2_X2 _35783_ (.A(\bp_fe_pc_gen_1.icache_pc_gen_i [21]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [21]),
    .S(_10026_),
    .Z(fe_queue_o[81]));
 MUX2_X2 _35784_ (.A(\bp_fe_pc_gen_1.icache_pc_gen_i [22]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [22]),
    .S(_10026_),
    .Z(fe_queue_o[82]));
 MUX2_X2 _35785_ (.A(\bp_fe_pc_gen_1.icache_pc_gen_i [23]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [23]),
    .S(_10026_),
    .Z(fe_queue_o[83]));
 MUX2_X2 _35786_ (.A(\bp_fe_pc_gen_1.icache_pc_gen_i [24]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [24]),
    .S(_10026_),
    .Z(fe_queue_o[84]));
 MUX2_X2 _35787_ (.A(\bp_fe_pc_gen_1.icache_pc_gen_i [25]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [25]),
    .S(_10026_),
    .Z(fe_queue_o[85]));
 BUF_X8 _35788_ (.A(_08643_),
    .Z(_10027_));
 MUX2_X2 _35789_ (.A(\bp_fe_pc_gen_1.icache_pc_gen_i [26]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [26]),
    .S(_10027_),
    .Z(fe_queue_o[86]));
 MUX2_X2 _35790_ (.A(\bp_fe_pc_gen_1.icache_pc_gen_i [27]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [27]),
    .S(_10027_),
    .Z(fe_queue_o[87]));
 MUX2_X2 _35791_ (.A(\bp_fe_pc_gen_1.icache_pc_gen_i [28]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [28]),
    .S(_10027_),
    .Z(fe_queue_o[88]));
 MUX2_X2 _35792_ (.A(\bp_fe_pc_gen_1.icache_pc_gen_i [29]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [29]),
    .S(_10027_),
    .Z(fe_queue_o[89]));
 MUX2_X2 _35793_ (.A(\bp_fe_pc_gen_1.icache_pc_gen_i [30]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [30]),
    .S(_10027_),
    .Z(fe_queue_o[90]));
 MUX2_X2 _35794_ (.A(\bp_fe_pc_gen_1.icache_pc_gen_i [31]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [31]),
    .S(_10027_),
    .Z(fe_queue_o[91]));
 MUX2_X2 _35795_ (.A(\bp_fe_pc_gen_1.icache_pc_gen_i [32]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [32]),
    .S(_10027_),
    .Z(fe_queue_o[92]));
 MUX2_X2 _35796_ (.A(\bp_fe_pc_gen_1.icache_pc_gen_i [33]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [33]),
    .S(_10027_),
    .Z(fe_queue_o[93]));
 MUX2_X2 _35797_ (.A(\bp_fe_pc_gen_1.icache_pc_gen_i [34]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [34]),
    .S(_10027_),
    .Z(fe_queue_o[94]));
 MUX2_X2 _35798_ (.A(\bp_fe_pc_gen_1.icache_pc_gen_i [35]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [35]),
    .S(_10027_),
    .Z(fe_queue_o[95]));
 MUX2_X2 _35799_ (.A(\bp_fe_pc_gen_1.icache_pc_gen_i [36]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [36]),
    .S(_08644_),
    .Z(fe_queue_o[96]));
 MUX2_X2 _35800_ (.A(\bp_fe_pc_gen_1.icache_pc_gen_i [37]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [37]),
    .S(_08644_),
    .Z(fe_queue_o[97]));
 MUX2_X2 _35801_ (.A(\bp_fe_pc_gen_1.icache_pc_gen_i [38]),
    .B(\bp_fe_pc_gen_1.pc_if2_r [38]),
    .S(_08644_),
    .Z(fe_queue_o[98]));
 XNOR2_X1 _35802_ (.A(_08981_),
    .B(\itlb.vtag_cam.mem [105]),
    .ZN(_10028_));
 AOI221_X2 _35803_ (.A(_10028_),
    .B1(\itlb.vtag_cam.mem [81]),
    .B2(_08784_),
    .C1(\itlb.vtag_cam.mem [89]),
    .C2(_08853_),
    .ZN(_10029_));
 XOR2_X2 _35804_ (.A(_08901_),
    .B(\itlb.vtag_cam.mem [95]),
    .Z(_10030_));
 OR2_X1 _35805_ (.A1(_08917_),
    .A2(\itlb.vtag_cam.mem [97]),
    .ZN(_10031_));
 NOR2_X4 _35806_ (.A1(_08808_),
    .A2(_08811_),
    .ZN(_10032_));
 BUF_X8 _35807_ (.A(_10032_),
    .Z(_10033_));
 NAND2_X2 _35808_ (.A1(_10033_),
    .A2(\itlb.vtag_cam.mem [84]),
    .ZN(_10034_));
 NAND4_X4 _35809_ (.A1(_10029_),
    .A2(_10030_),
    .A3(_10031_),
    .A4(_10034_),
    .ZN(_10035_));
 NOR2_X4 _35810_ (.A1(_08856_),
    .A2(_08859_),
    .ZN(_10036_));
 INV_X1 _35811_ (.A(_10036_),
    .ZN(_10037_));
 INV_X1 _35812_ (.A(\itlb.vtag_cam.mem [90]),
    .ZN(_10038_));
 OAI22_X2 _35813_ (.A1(_10037_),
    .A2(_10038_),
    .B1(\itlb.vtag_cam.mem [85]),
    .B2(_08821_),
    .ZN(_10039_));
 INV_X1 _35814_ (.A(\itlb.vtag_cam.mem [100]),
    .ZN(_10040_));
 NOR2_X4 _35815_ (.A1(_08936_),
    .A2(_08939_),
    .ZN(_10041_));
 BUF_X8 _35816_ (.A(_10041_),
    .Z(_10042_));
 INV_X2 _35817_ (.A(_10042_),
    .ZN(_10043_));
 AOI221_X2 _35818_ (.A(_10039_),
    .B1(\itlb.vtag_cam.mem [85]),
    .B2(_08822_),
    .C1(_10040_),
    .C2(_10043_),
    .ZN(_10044_));
 NOR2_X1 _35819_ (.A1(_08997_),
    .A2(\itlb.vtag_cam.mem [107]),
    .ZN(_10045_));
 NOR2_X4 _35820_ (.A1(_08920_),
    .A2(_08923_),
    .ZN(_10046_));
 OAI22_X1 _35821_ (.A1(_10043_),
    .A2(_10040_),
    .B1(\itlb.vtag_cam.mem [98]),
    .B2(_10046_),
    .ZN(_10047_));
 AOI211_X2 _35822_ (.A(_10045_),
    .B(_10047_),
    .C1(\itlb.vtag_cam.mem [98]),
    .C2(_10046_),
    .ZN(_10048_));
 AND2_X1 _35823_ (.A1(_08933_),
    .A2(\itlb.vtag_cam.mem [99]),
    .ZN(_10049_));
 NOR2_X4 _35824_ (.A1(_08825_),
    .A2(_08828_),
    .ZN(_10050_));
 NOR2_X4 _35825_ (.A1(_08841_),
    .A2(_08844_),
    .ZN(_10051_));
 AOI221_X2 _35826_ (.A(_10049_),
    .B1(\itlb.vtag_cam.mem [86]),
    .B2(_10050_),
    .C1(\itlb.vtag_cam.mem [88]),
    .C2(_10051_),
    .ZN(_10052_));
 NOR2_X4 _35827_ (.A1(_08871_),
    .A2(_08874_),
    .ZN(_10053_));
 NOR2_X4 _35828_ (.A1(_08888_),
    .A2(_08891_),
    .ZN(_10054_));
 OAI22_X2 _35829_ (.A1(\itlb.vtag_cam.mem [92]),
    .A2(_10053_),
    .B1(_10054_),
    .B2(\itlb.vtag_cam.mem [94]),
    .ZN(_10055_));
 AOI221_X2 _35830_ (.A(_10055_),
    .B1(_10038_),
    .B2(_10037_),
    .C1(\itlb.vtag_cam.mem [107]),
    .C2(_08997_),
    .ZN(_10056_));
 NAND4_X4 _35831_ (.A1(_10044_),
    .A2(_10048_),
    .A3(_10052_),
    .A4(_10056_),
    .ZN(_10057_));
 NOR2_X4 _35832_ (.A1(_08904_),
    .A2(_08907_),
    .ZN(_10058_));
 BUF_X8 _35833_ (.A(_10058_),
    .Z(_10059_));
 AOI22_X2 _35834_ (.A1(\itlb.vtag_cam.mem [93]),
    .A2(_08885_),
    .B1(_10059_),
    .B2(\itlb.vtag_cam.mem [96]),
    .ZN(_10060_));
 BUF_X8 _35835_ (.A(_10054_),
    .Z(_10061_));
 NAND2_X1 _35836_ (.A1(_10061_),
    .A2(\itlb.vtag_cam.mem [94]),
    .ZN(_10062_));
 OAI211_X2 _35837_ (.A(_10060_),
    .B(_10062_),
    .C1(\itlb.vtag_cam.mem [93]),
    .C2(_08885_),
    .ZN(_10063_));
 BUF_X8 _35838_ (.A(_10053_),
    .Z(_10064_));
 AOI22_X1 _35839_ (.A1(\itlb.vtag_cam.mem [92]),
    .A2(_10064_),
    .B1(_08949_),
    .B2(\itlb.vtag_cam.mem [101]),
    .ZN(_10065_));
 NAND2_X1 _35840_ (.A1(_08917_),
    .A2(\itlb.vtag_cam.mem [97]),
    .ZN(_10066_));
 OAI211_X2 _35841_ (.A(_10065_),
    .B(_10066_),
    .C1(\itlb.vtag_cam.mem [96]),
    .C2(_10059_),
    .ZN(_10067_));
 NOR4_X4 _35842_ (.A1(_10035_),
    .A2(_10057_),
    .A3(_10063_),
    .A4(_10067_),
    .ZN(_10068_));
 INV_X1 _35843_ (.A(\itlb.vtag_cam.valid [4]),
    .ZN(_10069_));
 NOR2_X4 _35844_ (.A1(_08329_),
    .A2(reset_i),
    .ZN(_10070_));
 INV_X8 _35845_ (.A(_10070_),
    .ZN(_10071_));
 NOR2_X2 _35846_ (.A1(_08985_),
    .A2(_08988_),
    .ZN(_10072_));
 BUF_X8 _35847_ (.A(_10072_),
    .Z(_10073_));
 AOI211_X1 _35848_ (.A(_10069_),
    .B(_10071_),
    .C1(_10073_),
    .C2(\itlb.vtag_cam.mem [106]),
    .ZN(_10074_));
 OAI221_X1 _35849_ (.A(_10074_),
    .B1(\itlb.vtag_cam.mem [84]),
    .B2(_10033_),
    .C1(\itlb.vtag_cam.mem [99]),
    .C2(_08933_),
    .ZN(_10075_));
 NOR2_X4 _35850_ (.A1(_08789_),
    .A2(_08793_),
    .ZN(_10076_));
 BUF_X8 _35851_ (.A(_10076_),
    .Z(_10077_));
 AND2_X1 _35852_ (.A1(_10077_),
    .A2(\itlb.vtag_cam.mem [82]),
    .ZN(_10078_));
 NOR2_X4 _35853_ (.A1(_08969_),
    .A2(_08972_),
    .ZN(_10079_));
 BUF_X8 _35854_ (.A(_10079_),
    .Z(_10080_));
 NOR2_X1 _35855_ (.A1(_10080_),
    .A2(\itlb.vtag_cam.mem [104]),
    .ZN(_10081_));
 OAI22_X1 _35856_ (.A1(\itlb.vtag_cam.mem [82]),
    .A2(_10077_),
    .B1(_10073_),
    .B2(\itlb.vtag_cam.mem [106]),
    .ZN(_10082_));
 NOR4_X1 _35857_ (.A1(_10075_),
    .A2(_10078_),
    .A3(_10081_),
    .A4(_10082_),
    .ZN(_10083_));
 NOR2_X1 _35858_ (.A1(_08949_),
    .A2(\itlb.vtag_cam.mem [101]),
    .ZN(_10084_));
 NAND2_X1 _35859_ (.A1(_08838_),
    .A2(\itlb.vtag_cam.mem [87]),
    .ZN(_10085_));
 OAI21_X1 _35860_ (.A(_10085_),
    .B1(_08805_),
    .B2(\itlb.vtag_cam.mem [83]),
    .ZN(_10086_));
 AOI211_X2 _35861_ (.A(_10084_),
    .B(_10086_),
    .C1(\itlb.vtag_cam.mem [83]),
    .C2(_08805_),
    .ZN(_10087_));
 INV_X8 _35862_ (.A(_08868_),
    .ZN(_10088_));
 INV_X1 _35863_ (.A(\itlb.vtag_cam.mem [91]),
    .ZN(_10089_));
 NOR2_X4 _35864_ (.A1(_08952_),
    .A2(_08955_),
    .ZN(_10090_));
 BUF_X8 _35865_ (.A(_10090_),
    .Z(_10091_));
 AOI22_X1 _35866_ (.A1(_10088_),
    .A2(_10089_),
    .B1(_10091_),
    .B2(\itlb.vtag_cam.mem [102]),
    .ZN(_10092_));
 NAND2_X1 _35867_ (.A1(_10080_),
    .A2(\itlb.vtag_cam.mem [104]),
    .ZN(_10093_));
 OAI211_X1 _35868_ (.A(_10092_),
    .B(_10093_),
    .C1(\itlb.vtag_cam.mem [102]),
    .C2(_10091_),
    .ZN(_10094_));
 OAI22_X1 _35869_ (.A1(_10088_),
    .A2(_10089_),
    .B1(\itlb.vtag_cam.mem [103]),
    .B2(_08966_),
    .ZN(_10095_));
 AND2_X1 _35870_ (.A1(_08966_),
    .A2(\itlb.vtag_cam.mem [103]),
    .ZN(_10096_));
 NOR2_X1 _35871_ (.A1(_08838_),
    .A2(\itlb.vtag_cam.mem [87]),
    .ZN(_10097_));
 NOR4_X1 _35872_ (.A1(_10094_),
    .A2(_10095_),
    .A3(_10096_),
    .A4(_10097_),
    .ZN(_10098_));
 OAI22_X2 _35873_ (.A1(_08853_),
    .A2(\itlb.vtag_cam.mem [89]),
    .B1(\itlb.vtag_cam.mem [81]),
    .B2(_08784_),
    .ZN(_10099_));
 BUF_X8 _35874_ (.A(_10050_),
    .Z(_10100_));
 BUF_X8 _35875_ (.A(_10051_),
    .Z(_10101_));
 OAI22_X2 _35876_ (.A1(\itlb.vtag_cam.mem [86]),
    .A2(_10100_),
    .B1(_10101_),
    .B2(\itlb.vtag_cam.mem [88]),
    .ZN(_10102_));
 NOR2_X2 _35877_ (.A1(_10099_),
    .A2(_10102_),
    .ZN(_10103_));
 AND4_X1 _35878_ (.A1(_10083_),
    .A2(_10087_),
    .A3(_10098_),
    .A4(_10103_),
    .ZN(_10104_));
 AND2_X1 _35879_ (.A1(_10068_),
    .A2(_10104_),
    .ZN(_10105_));
 INV_X1 _35880_ (.A(_08916_),
    .ZN(_10106_));
 INV_X1 _35881_ (.A(\itlb.vtag_cam.mem [43]),
    .ZN(_10107_));
 AOI22_X4 _35882_ (.A1(_10106_),
    .A2(_10107_),
    .B1(_08933_),
    .B2(\itlb.vtag_cam.mem [45]),
    .ZN(_10108_));
 NAND2_X1 _35883_ (.A1(_08885_),
    .A2(\itlb.vtag_cam.mem [39]),
    .ZN(_10109_));
 OAI211_X1 _35884_ (.A(_10108_),
    .B(_10109_),
    .C1(\itlb.vtag_cam.mem [50]),
    .C2(_10080_),
    .ZN(_10110_));
 AOI22_X1 _35885_ (.A1(\itlb.vtag_cam.mem [30]),
    .A2(_10033_),
    .B1(_10080_),
    .B2(\itlb.vtag_cam.mem [50]),
    .ZN(_10111_));
 NAND2_X1 _35886_ (.A1(_10077_),
    .A2(\itlb.vtag_cam.mem [28]),
    .ZN(_10112_));
 OAI211_X1 _35887_ (.A(_10111_),
    .B(_10112_),
    .C1(\itlb.vtag_cam.mem [52]),
    .C2(_10073_),
    .ZN(_10113_));
 NOR2_X1 _35888_ (.A1(_10110_),
    .A2(_10113_),
    .ZN(_10114_));
 XOR2_X2 _35889_ (.A(_08804_),
    .B(\itlb.vtag_cam.mem [29]),
    .Z(_10115_));
 INV_X1 _35890_ (.A(\itlb.vtag_cam.mem [51]),
    .ZN(_10116_));
 INV_X4 _35891_ (.A(_08982_),
    .ZN(_10117_));
 OAI221_X2 _35892_ (.A(_10115_),
    .B1(\itlb.vtag_cam.mem [27]),
    .B2(_08784_),
    .C1(_10116_),
    .C2(_10117_),
    .ZN(_10118_));
 OAI22_X2 _35893_ (.A1(\itlb.vtag_cam.mem [41]),
    .A2(_08901_),
    .B1(_10042_),
    .B2(\itlb.vtag_cam.mem [46]),
    .ZN(_10119_));
 AND2_X1 _35894_ (.A1(_08900_),
    .A2(\itlb.vtag_cam.mem [41]),
    .ZN(_10120_));
 AOI21_X4 _35895_ (.A(\itlb.vtag_cam.mem [35]),
    .B1(net211),
    .B2(_08851_),
    .ZN(_10121_));
 NOR4_X4 _35896_ (.A1(_10118_),
    .A2(_10119_),
    .A3(_10120_),
    .A4(_10121_),
    .ZN(_10122_));
 INV_X2 _35897_ (.A(_08948_),
    .ZN(_10123_));
 INV_X1 _35898_ (.A(\itlb.vtag_cam.mem [47]),
    .ZN(_10124_));
 AOI22_X1 _35899_ (.A1(_10123_),
    .A2(_10124_),
    .B1(_10073_),
    .B2(\itlb.vtag_cam.mem [52]),
    .ZN(_10125_));
 NAND2_X1 _35900_ (.A1(_10061_),
    .A2(\itlb.vtag_cam.mem [40]),
    .ZN(_10126_));
 OAI211_X1 _35901_ (.A(_10125_),
    .B(_10126_),
    .C1(\itlb.vtag_cam.mem [32]),
    .C2(_10100_),
    .ZN(_10127_));
 NOR2_X1 _35902_ (.A1(_10061_),
    .A2(\itlb.vtag_cam.mem [40]),
    .ZN(_10128_));
 OAI22_X1 _35903_ (.A1(\itlb.vtag_cam.mem [34]),
    .A2(_10101_),
    .B1(_08885_),
    .B2(\itlb.vtag_cam.mem [39]),
    .ZN(_10129_));
 NOR3_X1 _35904_ (.A1(_10127_),
    .A2(_10128_),
    .A3(_10129_),
    .ZN(_10130_));
 OR2_X1 _35905_ (.A1(_10076_),
    .A2(\itlb.vtag_cam.mem [28]),
    .ZN(_10131_));
 NOR2_X1 _35906_ (.A1(_08821_),
    .A2(\itlb.vtag_cam.mem [31]),
    .ZN(_10132_));
 NAND2_X1 _35907_ (.A1(_08821_),
    .A2(\itlb.vtag_cam.mem [31]),
    .ZN(_10133_));
 OAI21_X1 _35908_ (.A(_10133_),
    .B1(\itlb.vtag_cam.mem [30]),
    .B2(_10032_),
    .ZN(_10134_));
 AOI211_X1 _35909_ (.A(_10132_),
    .B(_10134_),
    .C1(\itlb.vtag_cam.mem [35]),
    .C2(_08852_),
    .ZN(_10135_));
 NAND2_X1 _35910_ (.A1(_10064_),
    .A2(\itlb.vtag_cam.mem [38]),
    .ZN(_10136_));
 AOI22_X1 _35911_ (.A1(\itlb.vtag_cam.mem [43]),
    .A2(_08916_),
    .B1(_08949_),
    .B2(\itlb.vtag_cam.mem [47]),
    .ZN(_10137_));
 AND4_X1 _35912_ (.A1(_10131_),
    .A2(_10135_),
    .A3(_10136_),
    .A4(_10137_),
    .ZN(_10138_));
 AND4_X2 _35913_ (.A1(_10114_),
    .A2(_10122_),
    .A3(_10130_),
    .A4(_10138_),
    .ZN(_10139_));
 OAI22_X2 _35914_ (.A1(\itlb.vtag_cam.mem [45]),
    .A2(_08932_),
    .B1(_08965_),
    .B2(\itlb.vtag_cam.mem [49]),
    .ZN(_10140_));
 AOI221_X1 _35915_ (.A(_10140_),
    .B1(\itlb.vtag_cam.mem [32]),
    .B2(_10050_),
    .C1(\itlb.vtag_cam.mem [34]),
    .C2(_10051_),
    .ZN(_10141_));
 NAND2_X1 _35916_ (.A1(_08966_),
    .A2(\itlb.vtag_cam.mem [49]),
    .ZN(_10142_));
 OR2_X1 _35917_ (.A1(_10058_),
    .A2(\itlb.vtag_cam.mem [42]),
    .ZN(_10143_));
 NOR2_X1 _35918_ (.A1(_10053_),
    .A2(\itlb.vtag_cam.mem [38]),
    .ZN(_10144_));
 AOI21_X1 _35919_ (.A(_10144_),
    .B1(\itlb.vtag_cam.mem [42]),
    .B2(_10059_),
    .ZN(_10145_));
 AND4_X1 _35920_ (.A1(_10141_),
    .A2(_10142_),
    .A3(_10143_),
    .A4(_10145_),
    .ZN(_10146_));
 XOR2_X1 _35921_ (.A(_08997_),
    .B(\itlb.vtag_cam.mem [53]),
    .Z(_10147_));
 XOR2_X1 _35922_ (.A(_10046_),
    .B(\itlb.vtag_cam.mem [44]),
    .Z(_10148_));
 XOR2_X1 _35923_ (.A(_10091_),
    .B(\itlb.vtag_cam.mem [48]),
    .Z(_10149_));
 XOR2_X2 _35924_ (.A(_10036_),
    .B(\itlb.vtag_cam.mem [36]),
    .Z(_10150_));
 AND4_X1 _35925_ (.A1(_10147_),
    .A2(_10148_),
    .A3(_10149_),
    .A4(_10150_),
    .ZN(_10151_));
 NOR2_X1 _35926_ (.A1(_08837_),
    .A2(\itlb.vtag_cam.mem [33]),
    .ZN(_10152_));
 OAI211_X1 _35927_ (.A(\itlb.vtag_cam.valid [6]),
    .B(_10070_),
    .C1(_08868_),
    .C2(\itlb.vtag_cam.mem [37]),
    .ZN(_10153_));
 AOI211_X1 _35928_ (.A(_10152_),
    .B(_10153_),
    .C1(\itlb.vtag_cam.mem [37]),
    .C2(_08868_),
    .ZN(_10154_));
 AOI22_X1 _35929_ (.A1(\itlb.vtag_cam.mem [33]),
    .A2(_08838_),
    .B1(_10042_),
    .B2(\itlb.vtag_cam.mem [46]),
    .ZN(_10155_));
 AOI22_X1 _35930_ (.A1(_10117_),
    .A2(_10116_),
    .B1(_08784_),
    .B2(\itlb.vtag_cam.mem [27]),
    .ZN(_10156_));
 AND3_X2 _35931_ (.A1(_10154_),
    .A2(_10155_),
    .A3(_10156_),
    .ZN(_10157_));
 AND3_X2 _35932_ (.A1(_10146_),
    .A2(_10151_),
    .A3(_10157_),
    .ZN(_10158_));
 AOI21_X4 _35933_ (.A(_10105_),
    .B1(_10139_),
    .B2(_10158_),
    .ZN(_10159_));
 XOR2_X2 _35934_ (.A(_08965_),
    .B(\itlb.vtag_cam.mem [22]),
    .Z(_10160_));
 INV_X1 _35935_ (.A(\itlb.vtag_cam.mem [17]),
    .ZN(_10161_));
 INV_X4 _35936_ (.A(_10046_),
    .ZN(_10162_));
 OAI221_X2 _35937_ (.A(_10160_),
    .B1(\itlb.vtag_cam.mem [0]),
    .B2(_08784_),
    .C1(_10161_),
    .C2(_10162_),
    .ZN(_10163_));
 INV_X4 _35938_ (.A(_10091_),
    .ZN(_10164_));
 INV_X1 _35939_ (.A(\itlb.vtag_cam.mem [21]),
    .ZN(_10165_));
 AOI22_X1 _35940_ (.A1(_10164_),
    .A2(_10165_),
    .B1(_10054_),
    .B2(\itlb.vtag_cam.mem [13]),
    .ZN(_10166_));
 AOI22_X1 _35941_ (.A1(\itlb.vtag_cam.mem [1]),
    .A2(_10076_),
    .B1(_08948_),
    .B2(\itlb.vtag_cam.mem [20]),
    .ZN(_10167_));
 NAND2_X1 _35942_ (.A1(_10166_),
    .A2(_10167_),
    .ZN(_10168_));
 NAND2_X1 _35943_ (.A1(_10058_),
    .A2(\itlb.vtag_cam.mem [15]),
    .ZN(_10169_));
 OAI221_X2 _35944_ (.A(_10169_),
    .B1(\itlb.vtag_cam.mem [7]),
    .B2(_10051_),
    .C1(\itlb.vtag_cam.mem [16]),
    .C2(_08917_),
    .ZN(_10170_));
 INV_X4 _35945_ (.A(_10032_),
    .ZN(_10171_));
 INV_X1 _35946_ (.A(\itlb.vtag_cam.mem [3]),
    .ZN(_10172_));
 AOI22_X1 _35947_ (.A1(_10171_),
    .A2(_10172_),
    .B1(_10053_),
    .B2(\itlb.vtag_cam.mem [11]),
    .ZN(_10173_));
 NAND2_X1 _35948_ (.A1(_10051_),
    .A2(\itlb.vtag_cam.mem [7]),
    .ZN(_10174_));
 OAI211_X1 _35949_ (.A(_10173_),
    .B(_10174_),
    .C1(\itlb.vtag_cam.mem [11]),
    .C2(_10053_),
    .ZN(_10175_));
 NOR4_X1 _35950_ (.A1(_10163_),
    .A2(_10168_),
    .A3(_10170_),
    .A4(_10175_),
    .ZN(_10176_));
 OAI22_X1 _35951_ (.A1(\itlb.vtag_cam.mem [13]),
    .A2(_10054_),
    .B1(_08948_),
    .B2(\itlb.vtag_cam.mem [20]),
    .ZN(_10177_));
 INV_X1 _35952_ (.A(\itlb.vtag_cam.mem [25]),
    .ZN(_10178_));
 INV_X4 _35953_ (.A(_10072_),
    .ZN(_10179_));
 AOI221_X1 _35954_ (.A(_10177_),
    .B1(\itlb.vtag_cam.mem [5]),
    .B2(_10050_),
    .C1(_10178_),
    .C2(_10179_),
    .ZN(_10180_));
 XOR2_X2 _35955_ (.A(_08852_),
    .B(\itlb.vtag_cam.mem [8]),
    .Z(_10181_));
 OR3_X1 _35956_ (.A1(_08985_),
    .A2(_10178_),
    .A3(_08988_),
    .ZN(_10182_));
 INV_X1 _35957_ (.A(\itlb.vtag_cam.mem [18]),
    .ZN(_10183_));
 OR3_X1 _35958_ (.A1(_08928_),
    .A2(_10183_),
    .A3(_08931_),
    .ZN(_10184_));
 AND4_X1 _35959_ (.A1(_10180_),
    .A2(_10181_),
    .A3(_10182_),
    .A4(_10184_),
    .ZN(_10185_));
 XOR2_X2 _35960_ (.A(_08997_),
    .B(\itlb.vtag_cam.mem [26]),
    .Z(_10186_));
 OAI221_X2 _35961_ (.A(_10186_),
    .B1(\itlb.vtag_cam.mem [1]),
    .B2(_10076_),
    .C1(\itlb.vtag_cam.mem [24]),
    .C2(_08982_),
    .ZN(_10187_));
 AND2_X1 _35962_ (.A1(_08917_),
    .A2(\itlb.vtag_cam.mem [16]),
    .ZN(_10188_));
 NOR3_X1 _35963_ (.A1(_08808_),
    .A2(_10172_),
    .A3(_08811_),
    .ZN(_10189_));
 XNOR2_X1 _35964_ (.A(_08822_),
    .B(\itlb.vtag_cam.mem [4]),
    .ZN(_10190_));
 NOR4_X1 _35965_ (.A1(_10187_),
    .A2(_10188_),
    .A3(_10189_),
    .A4(_10190_),
    .ZN(_10191_));
 AND3_X2 _35966_ (.A1(_10176_),
    .A2(_10185_),
    .A3(_10191_),
    .ZN(_10192_));
 INV_X4 _35967_ (.A(_08933_),
    .ZN(_10193_));
 BUF_X8 _35968_ (.A(_10036_),
    .Z(_10194_));
 AOI22_X2 _35969_ (.A1(_10193_),
    .A2(_10183_),
    .B1(_10194_),
    .B2(\itlb.vtag_cam.mem [9]),
    .ZN(_10195_));
 OAI221_X2 _35970_ (.A(_10195_),
    .B1(\itlb.vtag_cam.mem [15]),
    .B2(_10058_),
    .C1(_10165_),
    .C2(_10164_),
    .ZN(_10196_));
 OAI22_X2 _35971_ (.A1(\itlb.vtag_cam.mem [5]),
    .A2(_10050_),
    .B1(_08885_),
    .B2(\itlb.vtag_cam.mem [12]),
    .ZN(_10197_));
 AND2_X1 _35972_ (.A1(_08885_),
    .A2(\itlb.vtag_cam.mem [12]),
    .ZN(_10198_));
 NOR2_X1 _35973_ (.A1(_10194_),
    .A2(\itlb.vtag_cam.mem [9]),
    .ZN(_10199_));
 NOR4_X4 _35974_ (.A1(_10196_),
    .A2(_10197_),
    .A3(_10198_),
    .A4(_10199_),
    .ZN(_10200_));
 NAND2_X1 _35975_ (.A1(_08838_),
    .A2(\itlb.vtag_cam.mem [6]),
    .ZN(_10201_));
 OAI21_X1 _35976_ (.A(_10201_),
    .B1(_08805_),
    .B2(\itlb.vtag_cam.mem [2]),
    .ZN(_10202_));
 NAND2_X1 _35977_ (.A1(_08900_),
    .A2(\itlb.vtag_cam.mem [14]),
    .ZN(_10203_));
 OAI21_X1 _35978_ (.A(_10203_),
    .B1(\itlb.vtag_cam.mem [6]),
    .B2(_08838_),
    .ZN(_10204_));
 XNOR2_X1 _35979_ (.A(_10079_),
    .B(\itlb.vtag_cam.mem [23]),
    .ZN(_10205_));
 BUF_X4 _35980_ (.A(_10070_),
    .Z(_10206_));
 OAI211_X2 _35981_ (.A(\itlb.vtag_cam.valid [7]),
    .B(_10206_),
    .C1(_08900_),
    .C2(\itlb.vtag_cam.mem [14]),
    .ZN(_10207_));
 NOR4_X1 _35982_ (.A1(_10202_),
    .A2(_10204_),
    .A3(_10205_),
    .A4(_10207_),
    .ZN(_10208_));
 XOR2_X1 _35983_ (.A(_08868_),
    .B(\itlb.vtag_cam.mem [10]),
    .Z(_10209_));
 AOI22_X1 _35984_ (.A1(_08804_),
    .A2(\itlb.vtag_cam.mem [2]),
    .B1(\itlb.vtag_cam.mem [0]),
    .B2(_08784_),
    .ZN(_10210_));
 XOR2_X1 _35985_ (.A(_10042_),
    .B(\itlb.vtag_cam.mem [19]),
    .Z(_10211_));
 AOI22_X4 _35986_ (.A1(_10162_),
    .A2(_10161_),
    .B1(_08981_),
    .B2(\itlb.vtag_cam.mem [24]),
    .ZN(_10212_));
 AND4_X1 _35987_ (.A1(_10209_),
    .A2(_10210_),
    .A3(_10211_),
    .A4(_10212_),
    .ZN(_10213_));
 AND3_X2 _35988_ (.A1(_10200_),
    .A2(_10208_),
    .A3(_10213_),
    .ZN(_10214_));
 OAI22_X1 _35989_ (.A1(\itlb.vtag_cam.mem [65]),
    .A2(_10064_),
    .B1(_10061_),
    .B2(\itlb.vtag_cam.mem [67]),
    .ZN(_10215_));
 NAND3_X2 _35990_ (.A1(net210),
    .A2(\itlb.vtag_cam.mem [62]),
    .A3(_08851_),
    .ZN(_10216_));
 OR2_X1 _35991_ (.A1(_08822_),
    .A2(\itlb.vtag_cam.mem [58]),
    .ZN(_10217_));
 OR2_X1 _35992_ (.A1(_10073_),
    .A2(\itlb.vtag_cam.mem [79]),
    .ZN(_10218_));
 NAND2_X1 _35993_ (.A1(_10061_),
    .A2(\itlb.vtag_cam.mem [67]),
    .ZN(_10219_));
 NAND4_X1 _35994_ (.A1(_10216_),
    .A2(_10217_),
    .A3(_10218_),
    .A4(_10219_),
    .ZN(_10220_));
 AOI211_X1 _35995_ (.A(_10215_),
    .B(_10220_),
    .C1(\itlb.vtag_cam.mem [61]),
    .C2(_10101_),
    .ZN(_10221_));
 INV_X1 _35996_ (.A(\itlb.vtag_cam.mem [72]),
    .ZN(_10222_));
 AOI22_X2 _35997_ (.A1(_10193_),
    .A2(_10222_),
    .B1(_08965_),
    .B2(\itlb.vtag_cam.mem [76]),
    .ZN(_10223_));
 OAI221_X2 _35998_ (.A(_10223_),
    .B1(\itlb.vtag_cam.mem [76]),
    .B2(_08966_),
    .C1(_08853_),
    .C2(\itlb.vtag_cam.mem [62]),
    .ZN(_10224_));
 AOI22_X2 _35999_ (.A1(\itlb.vtag_cam.mem [70]),
    .A2(_08917_),
    .B1(_10073_),
    .B2(\itlb.vtag_cam.mem [79]),
    .ZN(_10225_));
 OAI221_X2 _36000_ (.A(_10225_),
    .B1(\itlb.vtag_cam.mem [59]),
    .B2(_10050_),
    .C1(\itlb.vtag_cam.mem [74]),
    .C2(_08949_),
    .ZN(_10226_));
 NOR2_X1 _36001_ (.A1(_10224_),
    .A2(_10226_),
    .ZN(_10227_));
 NAND2_X1 _36002_ (.A1(_10221_),
    .A2(_10227_),
    .ZN(_10228_));
 NAND2_X1 _36003_ (.A1(_10100_),
    .A2(\itlb.vtag_cam.mem [59]),
    .ZN(_10229_));
 AOI22_X4 _36004_ (.A1(\itlb.vtag_cam.mem [58]),
    .A2(_08822_),
    .B1(_10059_),
    .B2(\itlb.vtag_cam.mem [69]),
    .ZN(_10230_));
 OAI211_X2 _36005_ (.A(_10229_),
    .B(_10230_),
    .C1(_08805_),
    .C2(\itlb.vtag_cam.mem [56]),
    .ZN(_10231_));
 INV_X1 _36006_ (.A(\itlb.vtag_cam.mem [54]),
    .ZN(_10232_));
 INV_X8 _36007_ (.A(_08783_),
    .ZN(_10233_));
 AOI22_X2 _36008_ (.A1(_08805_),
    .A2(\itlb.vtag_cam.mem [56]),
    .B1(_10232_),
    .B2(_10233_),
    .ZN(_10234_));
 OAI221_X2 _36009_ (.A(_10234_),
    .B1(_10232_),
    .B2(_10233_),
    .C1(\itlb.vtag_cam.mem [57]),
    .C2(_10033_),
    .ZN(_10235_));
 OAI22_X1 _36010_ (.A1(\itlb.vtag_cam.mem [55]),
    .A2(_10077_),
    .B1(_10080_),
    .B2(\itlb.vtag_cam.mem [77]),
    .ZN(_10236_));
 OAI22_X2 _36011_ (.A1(\itlb.vtag_cam.mem [69]),
    .A2(_10059_),
    .B1(_08917_),
    .B2(\itlb.vtag_cam.mem [70]),
    .ZN(_10237_));
 NOR2_X1 _36012_ (.A1(_10236_),
    .A2(_10237_),
    .ZN(_10238_));
 XOR2_X2 _36013_ (.A(_08837_),
    .B(\itlb.vtag_cam.mem [60]),
    .Z(_10239_));
 OR2_X1 _36014_ (.A1(_08885_),
    .A2(\itlb.vtag_cam.mem [66]),
    .ZN(_10240_));
 NAND2_X1 _36015_ (.A1(_08949_),
    .A2(\itlb.vtag_cam.mem [74]),
    .ZN(_10241_));
 NAND4_X2 _36016_ (.A1(_10238_),
    .A2(_10239_),
    .A3(_10240_),
    .A4(_10241_),
    .ZN(_10242_));
 NOR4_X4 _36017_ (.A1(_10228_),
    .A2(_10231_),
    .A3(_10235_),
    .A4(_10242_),
    .ZN(_10243_));
 AOI22_X2 _36018_ (.A1(\itlb.vtag_cam.mem [57]),
    .A2(_10033_),
    .B1(_08884_),
    .B2(\itlb.vtag_cam.mem [66]),
    .ZN(_10244_));
 OAI221_X2 _36019_ (.A(_10244_),
    .B1(\itlb.vtag_cam.mem [61]),
    .B2(_10101_),
    .C1(_10222_),
    .C2(_10193_),
    .ZN(_10245_));
 XNOR2_X2 _36020_ (.A(_10194_),
    .B(\itlb.vtag_cam.mem [63]),
    .ZN(_10246_));
 AND2_X1 _36021_ (.A1(_10077_),
    .A2(\itlb.vtag_cam.mem [55]),
    .ZN(_10247_));
 INV_X1 _36022_ (.A(\itlb.vtag_cam.valid [5]),
    .ZN(_10248_));
 OR3_X1 _36023_ (.A1(_08329_),
    .A2(_08516_),
    .A3(_10248_),
    .ZN(_10249_));
 NOR4_X1 _36024_ (.A1(_10245_),
    .A2(_10246_),
    .A3(_10247_),
    .A4(_10249_),
    .ZN(_10250_));
 XNOR2_X1 _36025_ (.A(_08997_),
    .B(\itlb.vtag_cam.mem [80]),
    .ZN(_10251_));
 XNOR2_X1 _36026_ (.A(_10042_),
    .B(\itlb.vtag_cam.mem [73]),
    .ZN(_10252_));
 NOR2_X1 _36027_ (.A1(_10251_),
    .A2(_10252_),
    .ZN(_10253_));
 NOR2_X1 _36028_ (.A1(_08901_),
    .A2(\itlb.vtag_cam.mem [68]),
    .ZN(_10254_));
 INV_X1 _36029_ (.A(\itlb.vtag_cam.mem [68]),
    .ZN(_10255_));
 OR3_X1 _36030_ (.A1(_08896_),
    .A2(_10255_),
    .A3(_08899_),
    .ZN(_10256_));
 OAI21_X1 _36031_ (.A(_10256_),
    .B1(\itlb.vtag_cam.mem [78]),
    .B2(_08982_),
    .ZN(_10257_));
 AOI211_X2 _36032_ (.A(_10254_),
    .B(_10257_),
    .C1(\itlb.vtag_cam.mem [78]),
    .C2(_08982_),
    .ZN(_10258_));
 XOR2_X1 _36033_ (.A(_10046_),
    .B(\itlb.vtag_cam.mem [71]),
    .Z(_10259_));
 XOR2_X1 _36034_ (.A(_10091_),
    .B(\itlb.vtag_cam.mem [75]),
    .Z(_10260_));
 XOR2_X1 _36035_ (.A(_08868_),
    .B(\itlb.vtag_cam.mem [64]),
    .Z(_10261_));
 AOI22_X1 _36036_ (.A1(\itlb.vtag_cam.mem [65]),
    .A2(_10064_),
    .B1(_10080_),
    .B2(\itlb.vtag_cam.mem [77]),
    .ZN(_10262_));
 AND4_X1 _36037_ (.A1(_10259_),
    .A2(_10260_),
    .A3(_10261_),
    .A4(_10262_),
    .ZN(_10263_));
 AND4_X4 _36038_ (.A1(_10250_),
    .A2(_10253_),
    .A3(_10258_),
    .A4(_10263_),
    .ZN(_10264_));
 AOI22_X4 _36039_ (.A1(_10192_),
    .A2(_10214_),
    .B1(_10243_),
    .B2(_10264_),
    .ZN(_10265_));
 AND2_X4 _36040_ (.A1(_10159_),
    .A2(_10265_),
    .ZN(_10266_));
 NOR2_X1 _36041_ (.A1(_10100_),
    .A2(\itlb.vtag_cam.mem [113]),
    .ZN(_10267_));
 INV_X4 _36042_ (.A(_08997_),
    .ZN(_10268_));
 INV_X1 _36043_ (.A(\itlb.vtag_cam.mem [134]),
    .ZN(_10269_));
 OAI22_X1 _36044_ (.A1(_10268_),
    .A2(_10269_),
    .B1(\itlb.vtag_cam.mem [127]),
    .B2(_10042_),
    .ZN(_10270_));
 AOI211_X4 _36045_ (.A(_10267_),
    .B(_10270_),
    .C1(\itlb.vtag_cam.mem [127]),
    .C2(_10042_),
    .ZN(_10271_));
 INV_X1 _36046_ (.A(\itlb.vtag_cam.mem [118]),
    .ZN(_10272_));
 AOI22_X1 _36047_ (.A1(_08804_),
    .A2(\itlb.vtag_cam.mem [110]),
    .B1(_10272_),
    .B2(_10088_),
    .ZN(_10273_));
 NAND2_X1 _36048_ (.A1(_08821_),
    .A2(\itlb.vtag_cam.mem [112]),
    .ZN(_10274_));
 OAI211_X1 _36049_ (.A(_10273_),
    .B(_10274_),
    .C1(\itlb.vtag_cam.mem [110]),
    .C2(_08804_),
    .ZN(_10275_));
 NOR2_X1 _36050_ (.A1(_08783_),
    .A2(\itlb.vtag_cam.mem [108]),
    .ZN(_10276_));
 AOI21_X1 _36051_ (.A(_10276_),
    .B1(\itlb.vtag_cam.mem [132]),
    .B2(_08981_),
    .ZN(_10277_));
 OAI221_X1 _36052_ (.A(_10277_),
    .B1(_10272_),
    .B2(_10088_),
    .C1(\itlb.vtag_cam.mem [132]),
    .C2(_08981_),
    .ZN(_10278_));
 NOR2_X1 _36053_ (.A1(_10275_),
    .A2(_10278_),
    .ZN(_10279_));
 INV_X1 _36054_ (.A(\itlb.vtag_cam.mem [125]),
    .ZN(_10280_));
 OAI22_X1 _36055_ (.A1(_10162_),
    .A2(_10280_),
    .B1(\itlb.vtag_cam.mem [129]),
    .B2(_10090_),
    .ZN(_10281_));
 AOI221_X1 _36056_ (.A(_10281_),
    .B1(\itlb.vtag_cam.mem [124]),
    .B2(_08916_),
    .C1(\itlb.vtag_cam.mem [129]),
    .C2(_10091_),
    .ZN(_10282_));
 INV_X2 _36057_ (.A(_10054_),
    .ZN(_10283_));
 INV_X1 _36058_ (.A(\itlb.vtag_cam.mem [121]),
    .ZN(_10284_));
 AOI22_X2 _36059_ (.A1(_10283_),
    .A2(_10284_),
    .B1(_08784_),
    .B2(\itlb.vtag_cam.mem [108]),
    .ZN(_10285_));
 AOI22_X1 _36060_ (.A1(_10162_),
    .A2(_10280_),
    .B1(_10050_),
    .B2(\itlb.vtag_cam.mem [113]),
    .ZN(_10286_));
 AND4_X1 _36061_ (.A1(_10279_),
    .A2(_10282_),
    .A3(_10285_),
    .A4(_10286_),
    .ZN(_10287_));
 OR2_X1 _36062_ (.A1(_08852_),
    .A2(\itlb.vtag_cam.mem [116]),
    .ZN(_10288_));
 OAI221_X2 _36063_ (.A(_10288_),
    .B1(\itlb.vtag_cam.mem [109]),
    .B2(_10076_),
    .C1(\itlb.vtag_cam.mem [117]),
    .C2(_10194_),
    .ZN(_10289_));
 NOR2_X1 _36064_ (.A1(_08884_),
    .A2(\itlb.vtag_cam.mem [120]),
    .ZN(_10290_));
 AOI21_X1 _36065_ (.A(_10290_),
    .B1(\itlb.vtag_cam.mem [131]),
    .B2(_10079_),
    .ZN(_10291_));
 NAND2_X1 _36066_ (.A1(_08948_),
    .A2(\itlb.vtag_cam.mem [128]),
    .ZN(_10292_));
 OAI211_X1 _36067_ (.A(_10291_),
    .B(_10292_),
    .C1(\itlb.vtag_cam.mem [124]),
    .C2(_08917_),
    .ZN(_10293_));
 XOR2_X2 _36068_ (.A(_10073_),
    .B(\itlb.vtag_cam.mem [133]),
    .Z(_10294_));
 OAI221_X2 _36069_ (.A(_10294_),
    .B1(\itlb.vtag_cam.mem [128]),
    .B2(_08948_),
    .C1(\itlb.vtag_cam.mem [131]),
    .C2(_10079_),
    .ZN(_10295_));
 INV_X1 _36070_ (.A(\itlb.vtag_cam.mem [111]),
    .ZN(_10296_));
 AOI22_X1 _36071_ (.A1(_10171_),
    .A2(_10296_),
    .B1(_10053_),
    .B2(\itlb.vtag_cam.mem [119]),
    .ZN(_10297_));
 NAND2_X1 _36072_ (.A1(_08884_),
    .A2(\itlb.vtag_cam.mem [120]),
    .ZN(_10298_));
 OAI211_X1 _36073_ (.A(_10297_),
    .B(_10298_),
    .C1(\itlb.vtag_cam.mem [119]),
    .C2(_10053_),
    .ZN(_10299_));
 NOR4_X1 _36074_ (.A1(_10289_),
    .A2(_10293_),
    .A3(_10295_),
    .A4(_10299_),
    .ZN(_10300_));
 AND2_X1 _36075_ (.A1(_10287_),
    .A2(_10300_),
    .ZN(_10301_));
 INV_X1 _36076_ (.A(\itlb.vtag_cam.valid [3]),
    .ZN(_10302_));
 NOR3_X1 _36077_ (.A1(_08329_),
    .A2(_08516_),
    .A3(_10302_),
    .ZN(_10303_));
 OAI21_X1 _36078_ (.A(_10303_),
    .B1(_08966_),
    .B2(\itlb.vtag_cam.mem [130]),
    .ZN(_10304_));
 AOI221_X4 _36079_ (.A(_10304_),
    .B1(\itlb.vtag_cam.mem [130]),
    .B2(_08966_),
    .C1(_10269_),
    .C2(_10268_),
    .ZN(_10305_));
 XOR2_X2 _36080_ (.A(_08837_),
    .B(\itlb.vtag_cam.mem [114]),
    .Z(_10306_));
 OAI221_X2 _36081_ (.A(_10306_),
    .B1(_10296_),
    .B2(_10171_),
    .C1(\itlb.vtag_cam.mem [122]),
    .C2(_08901_),
    .ZN(_10307_));
 XOR2_X2 _36082_ (.A(_08933_),
    .B(\itlb.vtag_cam.mem [126]),
    .Z(_10308_));
 OAI221_X2 _36083_ (.A(_10308_),
    .B1(_10284_),
    .B2(_10283_),
    .C1(\itlb.vtag_cam.mem [123]),
    .C2(_10059_),
    .ZN(_10309_));
 AOI22_X2 _36084_ (.A1(_08853_),
    .A2(\itlb.vtag_cam.mem [116]),
    .B1(\itlb.vtag_cam.mem [109]),
    .B2(_10076_),
    .ZN(_10310_));
 AOI22_X2 _36085_ (.A1(\itlb.vtag_cam.mem [115]),
    .A2(_10101_),
    .B1(_10194_),
    .B2(\itlb.vtag_cam.mem [117]),
    .ZN(_10311_));
 NAND2_X2 _36086_ (.A1(_10310_),
    .A2(_10311_),
    .ZN(_10312_));
 NOR2_X1 _36087_ (.A1(_10051_),
    .A2(\itlb.vtag_cam.mem [115]),
    .ZN(_10313_));
 AOI21_X1 _36088_ (.A(_10313_),
    .B1(\itlb.vtag_cam.mem [123]),
    .B2(_10059_),
    .ZN(_10314_));
 NAND2_X1 _36089_ (.A1(_08901_),
    .A2(\itlb.vtag_cam.mem [122]),
    .ZN(_10315_));
 OAI211_X2 _36090_ (.A(_10314_),
    .B(_10315_),
    .C1(\itlb.vtag_cam.mem [112]),
    .C2(_08822_),
    .ZN(_10316_));
 NOR4_X4 _36091_ (.A1(_10307_),
    .A2(_10309_),
    .A3(_10312_),
    .A4(_10316_),
    .ZN(_10317_));
 AND4_X1 _36092_ (.A1(_10271_),
    .A2(_10301_),
    .A3(_10305_),
    .A4(_10317_),
    .ZN(_10318_));
 AND2_X1 _36093_ (.A1(_10192_),
    .A2(_10214_),
    .ZN(_10319_));
 NOR2_X2 _36094_ (.A1(_10318_),
    .A2(_10319_),
    .ZN(_10320_));
 AND2_X1 _36095_ (.A1(_10243_),
    .A2(_10264_),
    .ZN(_10321_));
 NOR2_X1 _36096_ (.A1(_10042_),
    .A2(\itlb.vtag_cam.mem [181]),
    .ZN(_10322_));
 AOI21_X1 _36097_ (.A(_10322_),
    .B1(\itlb.vtag_cam.mem [168]),
    .B2(_08838_),
    .ZN(_10323_));
 AOI22_X1 _36098_ (.A1(\itlb.vtag_cam.mem [181]),
    .A2(_10042_),
    .B1(_08965_),
    .B2(\itlb.vtag_cam.mem [184]),
    .ZN(_10324_));
 INV_X1 _36099_ (.A(\itlb.vtag_cam.mem [185]),
    .ZN(_10325_));
 INV_X4 _36100_ (.A(_10080_),
    .ZN(_10326_));
 OAI221_X1 _36101_ (.A(_10324_),
    .B1(\itlb.vtag_cam.mem [168]),
    .B2(_08838_),
    .C1(_10325_),
    .C2(_10326_),
    .ZN(_10327_));
 AND2_X1 _36102_ (.A1(_10101_),
    .A2(\itlb.vtag_cam.mem [169]),
    .ZN(_10328_));
 NOR2_X1 _36103_ (.A1(_10064_),
    .A2(\itlb.vtag_cam.mem [173]),
    .ZN(_10329_));
 INV_X4 _36104_ (.A(_08822_),
    .ZN(_10330_));
 INV_X1 _36105_ (.A(\itlb.vtag_cam.mem [166]),
    .ZN(_10331_));
 OAI22_X2 _36106_ (.A1(_10330_),
    .A2(_10331_),
    .B1(_08933_),
    .B2(\itlb.vtag_cam.mem [180]),
    .ZN(_10332_));
 NOR4_X1 _36107_ (.A1(_10327_),
    .A2(_10328_),
    .A3(_10329_),
    .A4(_10332_),
    .ZN(_10333_));
 XOR2_X1 _36108_ (.A(_08901_),
    .B(\itlb.vtag_cam.mem [176]),
    .Z(_10334_));
 NOR2_X1 _36109_ (.A1(_08966_),
    .A2(\itlb.vtag_cam.mem [184]),
    .ZN(_10335_));
 INV_X1 _36110_ (.A(\itlb.vtag_cam.mem [172]),
    .ZN(_10336_));
 OAI22_X1 _36111_ (.A1(_10088_),
    .A2(_10336_),
    .B1(_08982_),
    .B2(\itlb.vtag_cam.mem [186]),
    .ZN(_10337_));
 AOI211_X1 _36112_ (.A(_10335_),
    .B(_10337_),
    .C1(\itlb.vtag_cam.mem [186]),
    .C2(_08982_),
    .ZN(_10338_));
 AND4_X1 _36113_ (.A1(_10323_),
    .A2(_10333_),
    .A3(_10334_),
    .A4(_10338_),
    .ZN(_10339_));
 INV_X1 _36114_ (.A(\itlb.vtag_cam.mem [162]),
    .ZN(_10340_));
 OAI22_X1 _36115_ (.A1(_08853_),
    .A2(\itlb.vtag_cam.mem [170]),
    .B1(_10340_),
    .B2(_10233_),
    .ZN(_10341_));
 AOI221_X4 _36116_ (.A(_10341_),
    .B1(\itlb.vtag_cam.mem [170]),
    .B2(_08853_),
    .C1(_10336_),
    .C2(_10088_),
    .ZN(_10342_));
 OAI211_X1 _36117_ (.A(\itlb.vtag_cam.valid [1]),
    .B(_10206_),
    .C1(_08805_),
    .C2(\itlb.vtag_cam.mem [164]),
    .ZN(_10343_));
 AOI221_X4 _36118_ (.A(_10343_),
    .B1(_10340_),
    .B2(_10233_),
    .C1(\itlb.vtag_cam.mem [164]),
    .C2(_08805_),
    .ZN(_10344_));
 NAND3_X1 _36119_ (.A1(_10339_),
    .A2(_10342_),
    .A3(_10344_),
    .ZN(_10345_));
 INV_X1 _36120_ (.A(\itlb.vtag_cam.mem [188]),
    .ZN(_10346_));
 OAI22_X1 _36121_ (.A1(_10268_),
    .A2(_10346_),
    .B1(_10091_),
    .B2(\itlb.vtag_cam.mem [183]),
    .ZN(_10347_));
 INV_X1 _36122_ (.A(\itlb.vtag_cam.mem [179]),
    .ZN(_10348_));
 AOI221_X1 _36123_ (.A(_10347_),
    .B1(_10348_),
    .B2(_10162_),
    .C1(\itlb.vtag_cam.mem [183]),
    .C2(_10091_),
    .ZN(_10349_));
 INV_X2 _36124_ (.A(_10058_),
    .ZN(_10350_));
 INV_X1 _36125_ (.A(\itlb.vtag_cam.mem [177]),
    .ZN(_10351_));
 OAI22_X2 _36126_ (.A1(_10350_),
    .A2(_10351_),
    .B1(_08884_),
    .B2(\itlb.vtag_cam.mem [174]),
    .ZN(_10352_));
 AOI221_X1 _36127_ (.A(_10352_),
    .B1(\itlb.vtag_cam.mem [174]),
    .B2(_08884_),
    .C1(_10346_),
    .C2(_10268_),
    .ZN(_10353_));
 OAI22_X1 _36128_ (.A1(_10162_),
    .A2(_10348_),
    .B1(_08916_),
    .B2(\itlb.vtag_cam.mem [178]),
    .ZN(_10354_));
 AOI221_X1 _36129_ (.A(_10354_),
    .B1(\itlb.vtag_cam.mem [165]),
    .B2(_10032_),
    .C1(\itlb.vtag_cam.mem [178]),
    .C2(_08916_),
    .ZN(_10355_));
 NOR2_X1 _36130_ (.A1(_10073_),
    .A2(\itlb.vtag_cam.mem [187]),
    .ZN(_10356_));
 OAI22_X1 _36131_ (.A1(\itlb.vtag_cam.mem [175]),
    .A2(_10061_),
    .B1(_08949_),
    .B2(\itlb.vtag_cam.mem [182]),
    .ZN(_10357_));
 AOI211_X2 _36132_ (.A(_10356_),
    .B(_10357_),
    .C1(\itlb.vtag_cam.mem [167]),
    .C2(_10100_),
    .ZN(_10358_));
 AND4_X1 _36133_ (.A1(_10349_),
    .A2(_10353_),
    .A3(_10355_),
    .A4(_10358_),
    .ZN(_10359_));
 OAI22_X1 _36134_ (.A1(\itlb.vtag_cam.mem [169]),
    .A2(_10101_),
    .B1(_10059_),
    .B2(\itlb.vtag_cam.mem [177]),
    .ZN(_10360_));
 AOI22_X2 _36135_ (.A1(_10326_),
    .A2(_10325_),
    .B1(_08949_),
    .B2(\itlb.vtag_cam.mem [182]),
    .ZN(_10361_));
 OAI221_X2 _36136_ (.A(_10361_),
    .B1(\itlb.vtag_cam.mem [165]),
    .B2(_10033_),
    .C1(\itlb.vtag_cam.mem [171]),
    .C2(_10194_),
    .ZN(_10362_));
 AOI211_X2 _36137_ (.A(_10360_),
    .B(_10362_),
    .C1(_10331_),
    .C2(_10330_),
    .ZN(_10363_));
 NOR2_X1 _36138_ (.A1(_10100_),
    .A2(\itlb.vtag_cam.mem [167]),
    .ZN(_10364_));
 AOI21_X1 _36139_ (.A(_10364_),
    .B1(\itlb.vtag_cam.mem [175]),
    .B2(_10061_),
    .ZN(_10365_));
 XOR2_X1 _36140_ (.A(_10077_),
    .B(\itlb.vtag_cam.mem [163]),
    .Z(_10366_));
 AOI22_X1 _36141_ (.A1(\itlb.vtag_cam.mem [173]),
    .A2(_10064_),
    .B1(_10073_),
    .B2(\itlb.vtag_cam.mem [187]),
    .ZN(_10367_));
 AOI22_X2 _36142_ (.A1(\itlb.vtag_cam.mem [171]),
    .A2(_10194_),
    .B1(_08933_),
    .B2(\itlb.vtag_cam.mem [180]),
    .ZN(_10368_));
 AND4_X1 _36143_ (.A1(_10365_),
    .A2(_10366_),
    .A3(_10367_),
    .A4(_10368_),
    .ZN(_10369_));
 NAND3_X2 _36144_ (.A1(_10359_),
    .A2(_10363_),
    .A3(_10369_),
    .ZN(_10370_));
 NOR2_X2 _36145_ (.A1(_10345_),
    .A2(_10370_),
    .ZN(_10371_));
 NOR2_X2 _36146_ (.A1(_10321_),
    .A2(_10371_),
    .ZN(_10372_));
 NAND2_X4 _36147_ (.A1(_10320_),
    .A2(_10372_),
    .ZN(_10373_));
 XOR2_X2 _36148_ (.A(_10091_),
    .B(\itlb.vtag_cam.mem [156]),
    .Z(_10374_));
 INV_X1 _36149_ (.A(\itlb.vtag_cam.valid [2]),
    .ZN(_10375_));
 NOR3_X4 _36150_ (.A1(_08329_),
    .A2(_08516_),
    .A3(_10375_),
    .ZN(_10376_));
 OAI211_X1 _36151_ (.A(_10374_),
    .B(_10376_),
    .C1(\itlb.vtag_cam.mem [159]),
    .C2(_08982_),
    .ZN(_10377_));
 XNOR2_X1 _36152_ (.A(_08901_),
    .B(\itlb.vtag_cam.mem [149]),
    .ZN(_10378_));
 XNOR2_X1 _36153_ (.A(_08838_),
    .B(\itlb.vtag_cam.mem [141]),
    .ZN(_10379_));
 NOR3_X1 _36154_ (.A1(_10377_),
    .A2(_10378_),
    .A3(_10379_),
    .ZN(_10380_));
 INV_X2 _36155_ (.A(_08965_),
    .ZN(_10381_));
 INV_X1 _36156_ (.A(\itlb.vtag_cam.mem [157]),
    .ZN(_10382_));
 AOI22_X2 _36157_ (.A1(_10381_),
    .A2(_10382_),
    .B1(_08981_),
    .B2(\itlb.vtag_cam.mem [159]),
    .ZN(_10383_));
 OAI221_X2 _36158_ (.A(_10383_),
    .B1(_10382_),
    .B2(_10381_),
    .C1(\itlb.vtag_cam.mem [161]),
    .C2(_08997_),
    .ZN(_10384_));
 NAND2_X1 _36159_ (.A1(_08997_),
    .A2(\itlb.vtag_cam.mem [161]),
    .ZN(_10385_));
 OAI21_X1 _36160_ (.A(_10385_),
    .B1(\itlb.vtag_cam.mem [154]),
    .B2(_10041_),
    .ZN(_10386_));
 AND2_X1 _36161_ (.A1(_10041_),
    .A2(\itlb.vtag_cam.mem [154]),
    .ZN(_10387_));
 NOR2_X1 _36162_ (.A1(_08821_),
    .A2(\itlb.vtag_cam.mem [139]),
    .ZN(_10388_));
 NOR4_X1 _36163_ (.A1(_10384_),
    .A2(_10386_),
    .A3(_10387_),
    .A4(_10388_),
    .ZN(_10389_));
 XOR2_X1 _36164_ (.A(_08783_),
    .B(\itlb.vtag_cam.mem [135]),
    .Z(_10390_));
 AOI22_X1 _36165_ (.A1(_08804_),
    .A2(\itlb.vtag_cam.mem [137]),
    .B1(\itlb.vtag_cam.mem [152]),
    .B2(_10046_),
    .ZN(_10391_));
 AOI21_X1 _36166_ (.A(\itlb.vtag_cam.mem [137]),
    .B1(net212),
    .B2(_08803_),
    .ZN(_10392_));
 INV_X2 _36167_ (.A(\itlb.vtag_cam.mem [145]),
    .ZN(_10393_));
 OAI22_X1 _36168_ (.A1(_10088_),
    .A2(_10393_),
    .B1(_10046_),
    .B2(\itlb.vtag_cam.mem [152]),
    .ZN(_10394_));
 AOI211_X1 _36169_ (.A(_10392_),
    .B(_10394_),
    .C1(\itlb.vtag_cam.mem [139]),
    .C2(_08822_),
    .ZN(_10395_));
 AND4_X1 _36170_ (.A1(_10389_),
    .A2(_10390_),
    .A3(_10391_),
    .A4(_10395_),
    .ZN(_10396_));
 NOR2_X1 _36171_ (.A1(_10076_),
    .A2(\itlb.vtag_cam.mem [136]),
    .ZN(_10397_));
 AOI21_X1 _36172_ (.A(_10397_),
    .B1(\itlb.vtag_cam.mem [144]),
    .B2(_10194_),
    .ZN(_10398_));
 OAI221_X2 _36173_ (.A(_10398_),
    .B1(\itlb.vtag_cam.mem [144]),
    .B2(_10194_),
    .C1(\itlb.vtag_cam.mem [143]),
    .C2(_08852_),
    .ZN(_10399_));
 NOR2_X1 _36174_ (.A1(_08916_),
    .A2(\itlb.vtag_cam.mem [151]),
    .ZN(_10400_));
 AOI21_X1 _36175_ (.A(_10400_),
    .B1(\itlb.vtag_cam.mem [155]),
    .B2(_08948_),
    .ZN(_10401_));
 NAND2_X1 _36176_ (.A1(_10079_),
    .A2(\itlb.vtag_cam.mem [158]),
    .ZN(_10402_));
 OAI211_X1 _36177_ (.A(_10401_),
    .B(_10402_),
    .C1(\itlb.vtag_cam.mem [147]),
    .C2(_08885_),
    .ZN(_10403_));
 AOI22_X2 _36178_ (.A1(\itlb.vtag_cam.mem [146]),
    .A2(_10053_),
    .B1(_08884_),
    .B2(\itlb.vtag_cam.mem [147]),
    .ZN(_10404_));
 INV_X1 _36179_ (.A(\itlb.vtag_cam.mem [150]),
    .ZN(_10405_));
 OAI221_X2 _36180_ (.A(_10404_),
    .B1(\itlb.vtag_cam.mem [138]),
    .B2(_10033_),
    .C1(_10405_),
    .C2(_10350_),
    .ZN(_10406_));
 INV_X1 _36181_ (.A(\itlb.vtag_cam.mem [142]),
    .ZN(_10407_));
 OR3_X1 _36182_ (.A1(_08841_),
    .A2(_10407_),
    .A3(_08844_),
    .ZN(_10408_));
 OAI21_X1 _36183_ (.A(_10407_),
    .B1(_08841_),
    .B2(_08844_),
    .ZN(_10409_));
 OAI211_X2 _36184_ (.A(_10408_),
    .B(_10409_),
    .C1(\itlb.vtag_cam.mem [146]),
    .C2(_10064_),
    .ZN(_10410_));
 NOR4_X1 _36185_ (.A1(_10399_),
    .A2(_10403_),
    .A3(_10406_),
    .A4(_10410_),
    .ZN(_10411_));
 AOI22_X2 _36186_ (.A1(_08852_),
    .A2(\itlb.vtag_cam.mem [143]),
    .B1(_10393_),
    .B2(_10088_),
    .ZN(_10412_));
 OAI221_X2 _36187_ (.A(_10412_),
    .B1(\itlb.vtag_cam.mem [158]),
    .B2(_10080_),
    .C1(\itlb.vtag_cam.mem [160]),
    .C2(_10073_),
    .ZN(_10413_));
 AOI22_X1 _36188_ (.A1(\itlb.vtag_cam.mem [136]),
    .A2(_10076_),
    .B1(_10050_),
    .B2(\itlb.vtag_cam.mem [140]),
    .ZN(_10414_));
 INV_X1 _36189_ (.A(\itlb.vtag_cam.mem [160]),
    .ZN(_10415_));
 OAI221_X1 _36190_ (.A(_10414_),
    .B1(\itlb.vtag_cam.mem [140]),
    .B2(_10050_),
    .C1(_10415_),
    .C2(_10179_),
    .ZN(_10416_));
 AOI22_X2 _36191_ (.A1(\itlb.vtag_cam.mem [138]),
    .A2(_10032_),
    .B1(_10054_),
    .B2(\itlb.vtag_cam.mem [148]),
    .ZN(_10417_));
 OAI221_X2 _36192_ (.A(_10417_),
    .B1(\itlb.vtag_cam.mem [148]),
    .B2(_10061_),
    .C1(\itlb.vtag_cam.mem [150]),
    .C2(_10058_),
    .ZN(_10418_));
 XOR2_X1 _36193_ (.A(_08933_),
    .B(\itlb.vtag_cam.mem [153]),
    .Z(_10419_));
 NAND2_X1 _36194_ (.A1(_08916_),
    .A2(\itlb.vtag_cam.mem [151]),
    .ZN(_10420_));
 OAI211_X1 _36195_ (.A(_10419_),
    .B(_10420_),
    .C1(\itlb.vtag_cam.mem [155]),
    .C2(_08949_),
    .ZN(_10421_));
 NOR4_X1 _36196_ (.A1(_10413_),
    .A2(_10416_),
    .A3(_10418_),
    .A4(_10421_),
    .ZN(_10422_));
 AND4_X2 _36197_ (.A1(_10380_),
    .A2(_10396_),
    .A3(_10411_),
    .A4(_10422_),
    .ZN(_10423_));
 AOI21_X4 _36198_ (.A(_10423_),
    .B1(_10139_),
    .B2(_10158_),
    .ZN(_10424_));
 INV_X1 _36199_ (.A(\itlb.vtag_cam.mem [189]),
    .ZN(_10425_));
 OAI22_X2 _36200_ (.A1(_10233_),
    .A2(_10425_),
    .B1(_08982_),
    .B2(\itlb.vtag_cam.mem [213]),
    .ZN(_10426_));
 AOI221_X2 _36201_ (.A(_10426_),
    .B1(\itlb.vtag_cam.mem [190]),
    .B2(_10077_),
    .C1(\itlb.vtag_cam.mem [213]),
    .C2(_08982_),
    .ZN(_10427_));
 AOI22_X1 _36202_ (.A1(\itlb.vtag_cam.mem [194]),
    .A2(_10100_),
    .B1(_10101_),
    .B2(\itlb.vtag_cam.mem [196]),
    .ZN(_10428_));
 OAI221_X1 _36203_ (.A(_10428_),
    .B1(\itlb.vtag_cam.mem [200]),
    .B2(_10064_),
    .C1(\itlb.vtag_cam.mem [202]),
    .C2(_10061_),
    .ZN(_10429_));
 NAND2_X1 _36204_ (.A1(_10033_),
    .A2(\itlb.vtag_cam.mem [192]),
    .ZN(_10430_));
 OAI21_X1 _36205_ (.A(_10430_),
    .B1(\itlb.vtag_cam.mem [212]),
    .B2(_10080_),
    .ZN(_10431_));
 AND2_X1 _36206_ (.A1(_10064_),
    .A2(\itlb.vtag_cam.mem [200]),
    .ZN(_10432_));
 NOR2_X1 _36207_ (.A1(_10101_),
    .A2(\itlb.vtag_cam.mem [196]),
    .ZN(_10433_));
 NOR4_X1 _36208_ (.A1(_10429_),
    .A2(_10431_),
    .A3(_10432_),
    .A4(_10433_),
    .ZN(_10434_));
 INV_X1 _36209_ (.A(\itlb.vtag_cam.mem [209]),
    .ZN(_10435_));
 AOI22_X1 _36210_ (.A1(_10123_),
    .A2(_10435_),
    .B1(_10059_),
    .B2(\itlb.vtag_cam.mem [204]),
    .ZN(_10436_));
 XOR2_X1 _36211_ (.A(_08933_),
    .B(\itlb.vtag_cam.mem [207]),
    .Z(_10437_));
 AND4_X1 _36212_ (.A1(_10427_),
    .A2(_10434_),
    .A3(_10436_),
    .A4(_10437_),
    .ZN(_10438_));
 XOR2_X1 _36213_ (.A(_08997_),
    .B(\itlb.vtag_cam.mem [215]),
    .Z(_10439_));
 INV_X1 _36214_ (.A(\itlb.vtag_cam.valid [0]),
    .ZN(_10440_));
 NOR3_X2 _36215_ (.A1(_08329_),
    .A2(_08516_),
    .A3(_10440_),
    .ZN(_10441_));
 OAI211_X1 _36216_ (.A(_10439_),
    .B(_10441_),
    .C1(\itlb.vtag_cam.mem [194]),
    .C2(_10100_),
    .ZN(_10442_));
 XNOR2_X1 _36217_ (.A(_10046_),
    .B(\itlb.vtag_cam.mem [206]),
    .ZN(_10443_));
 XNOR2_X1 _36218_ (.A(_10042_),
    .B(\itlb.vtag_cam.mem [208]),
    .ZN(_10444_));
 NOR3_X1 _36219_ (.A1(_10442_),
    .A2(_10443_),
    .A3(_10444_),
    .ZN(_10445_));
 AND2_X1 _36220_ (.A1(_10438_),
    .A2(_10445_),
    .ZN(_10446_));
 OAI22_X1 _36221_ (.A1(_08853_),
    .A2(\itlb.vtag_cam.mem [197]),
    .B1(\itlb.vtag_cam.mem [189]),
    .B2(_08784_),
    .ZN(_10447_));
 INV_X2 _36222_ (.A(\itlb.vtag_cam.mem [195]),
    .ZN(_10448_));
 INV_X2 _36223_ (.A(_08838_),
    .ZN(_10449_));
 AOI221_X4 _36224_ (.A(_10447_),
    .B1(_10448_),
    .B2(_10449_),
    .C1(\itlb.vtag_cam.mem [197]),
    .C2(_08853_),
    .ZN(_10450_));
 INV_X1 _36225_ (.A(\itlb.vtag_cam.mem [214]),
    .ZN(_10451_));
 AOI22_X1 _36226_ (.A1(_10179_),
    .A2(_10451_),
    .B1(_10080_),
    .B2(\itlb.vtag_cam.mem [212]),
    .ZN(_10452_));
 XOR2_X2 _36227_ (.A(_08805_),
    .B(\itlb.vtag_cam.mem [191]),
    .Z(_10453_));
 NAND3_X1 _36228_ (.A1(_10450_),
    .A2(_10452_),
    .A3(_10453_),
    .ZN(_10454_));
 INV_X2 _36229_ (.A(_08885_),
    .ZN(_10455_));
 INV_X1 _36230_ (.A(\itlb.vtag_cam.mem [201]),
    .ZN(_10456_));
 AOI22_X1 _36231_ (.A1(_10455_),
    .A2(_10456_),
    .B1(_10061_),
    .B2(\itlb.vtag_cam.mem [202]),
    .ZN(_10457_));
 OAI221_X1 _36232_ (.A(_10457_),
    .B1(\itlb.vtag_cam.mem [190]),
    .B2(_10077_),
    .C1(\itlb.vtag_cam.mem [204]),
    .C2(_10059_),
    .ZN(_10458_));
 XOR2_X2 _36233_ (.A(_10194_),
    .B(\itlb.vtag_cam.mem [198]),
    .Z(_10459_));
 OAI221_X2 _36234_ (.A(_10459_),
    .B1(\itlb.vtag_cam.mem [192]),
    .B2(_10033_),
    .C1(_10451_),
    .C2(_10179_),
    .ZN(_10460_));
 NOR3_X1 _36235_ (.A1(_10454_),
    .A2(_10458_),
    .A3(_10460_),
    .ZN(_10461_));
 XOR2_X2 _36236_ (.A(_08822_),
    .B(\itlb.vtag_cam.mem [193]),
    .Z(_10462_));
 INV_X1 _36237_ (.A(\itlb.vtag_cam.mem [210]),
    .ZN(_10463_));
 OAI221_X1 _36238_ (.A(_10462_),
    .B1(_10456_),
    .B2(_10455_),
    .C1(_10463_),
    .C2(_10164_),
    .ZN(_10464_));
 XOR2_X1 _36239_ (.A(_08901_),
    .B(\itlb.vtag_cam.mem [203]),
    .Z(_10465_));
 OR2_X1 _36240_ (.A1(_08917_),
    .A2(\itlb.vtag_cam.mem [205]),
    .ZN(_10466_));
 AOI22_X1 _36241_ (.A1(\itlb.vtag_cam.mem [205]),
    .A2(_08917_),
    .B1(_08949_),
    .B2(\itlb.vtag_cam.mem [209]),
    .ZN(_10467_));
 AOI22_X2 _36242_ (.A1(\itlb.vtag_cam.mem [199]),
    .A2(_08868_),
    .B1(_08966_),
    .B2(\itlb.vtag_cam.mem [211]),
    .ZN(_10468_));
 NAND4_X1 _36243_ (.A1(_10465_),
    .A2(_10466_),
    .A3(_10467_),
    .A4(_10468_),
    .ZN(_10469_));
 OAI22_X1 _36244_ (.A1(\itlb.vtag_cam.mem [199]),
    .A2(_08868_),
    .B1(_10091_),
    .B2(\itlb.vtag_cam.mem [210]),
    .ZN(_10470_));
 OAI22_X1 _36245_ (.A1(_10449_),
    .A2(_10448_),
    .B1(_08966_),
    .B2(\itlb.vtag_cam.mem [211]),
    .ZN(_10471_));
 NOR4_X1 _36246_ (.A1(_10464_),
    .A2(_10469_),
    .A3(_10470_),
    .A4(_10471_),
    .ZN(_10472_));
 NAND3_X2 _36247_ (.A1(_10446_),
    .A2(_10461_),
    .A3(_10472_),
    .ZN(_10473_));
 NAND2_X1 _36248_ (.A1(_10068_),
    .A2(_10104_),
    .ZN(_10474_));
 AND2_X1 _36249_ (.A1(_10473_),
    .A2(_10474_),
    .ZN(_10475_));
 NAND2_X4 _36250_ (.A1(_10424_),
    .A2(_10475_),
    .ZN(_10476_));
 OAI211_X4 _36251_ (.A(_10266_),
    .B(_08037_),
    .C1(_10373_),
    .C2(_10476_),
    .ZN(_10477_));
 NOR2_X4 _36252_ (.A1(_10373_),
    .A2(_10476_),
    .ZN(_10478_));
 NOR2_X4 _36253_ (.A1(_10478_),
    .A2(_08480_),
    .ZN(\itlb.r_v_reg.N3 ));
 OR2_X1 _36254_ (.A1(\itlb.r_v_reg.N3 ),
    .A2(_10071_),
    .ZN(_10479_));
 INV_X4 _36255_ (.A(\itlb.plru.encoder.N1 ),
    .ZN(_10480_));
 OAI21_X1 _36256_ (.A(_10477_),
    .B1(_10479_),
    .B2(_10480_),
    .ZN(_06817_));
 OAI211_X1 _36257_ (.A(\itlb.plru.encoder.lru_i [1]),
    .B(_10206_),
    .C1(_10478_),
    .C2(_08480_),
    .ZN(_10481_));
 INV_X1 _36258_ (.A(\itlb.r_v_reg.N3 ),
    .ZN(_10482_));
 INV_X1 _36259_ (.A(_10159_),
    .ZN(_10483_));
 INV_X1 _36260_ (.A(_10265_),
    .ZN(_10484_));
 OAI21_X1 _36261_ (.A(_00576_),
    .B1(_10483_),
    .B2(_10484_),
    .ZN(_10485_));
 INV_X1 _36262_ (.A(_10266_),
    .ZN(_10486_));
 AND2_X2 _36263_ (.A1(_10320_),
    .A2(_10424_),
    .ZN(_10487_));
 OAI21_X1 _36264_ (.A(_10485_),
    .B1(_10486_),
    .B2(_10487_),
    .ZN(_10488_));
 OAI21_X1 _36265_ (.A(_10481_),
    .B1(_10482_),
    .B2(_10488_),
    .ZN(_06818_));
 NOR2_X1 _36266_ (.A1(_10487_),
    .A2(_10266_),
    .ZN(_10489_));
 INV_X1 _36267_ (.A(_10489_),
    .ZN(_10490_));
 INV_X1 _36268_ (.A(_00577_),
    .ZN(_10491_));
 OAI211_X1 _36269_ (.A(_10490_),
    .B(\itlb.r_v_reg.N3 ),
    .C1(_10491_),
    .C2(_10486_),
    .ZN(_10492_));
 OAI211_X1 _36270_ (.A(\itlb.plru.encoder.lru_i [2]),
    .B(_10206_),
    .C1(_10478_),
    .C2(_08480_),
    .ZN(_10493_));
 NAND2_X1 _36271_ (.A1(_10492_),
    .A2(_10493_),
    .ZN(_06819_));
 NAND3_X1 _36272_ (.A1(_10266_),
    .A2(_10320_),
    .A3(_10424_),
    .ZN(_10494_));
 NAND2_X1 _36273_ (.A1(_10494_),
    .A2(_00578_),
    .ZN(_10495_));
 INV_X1 _36274_ (.A(_10372_),
    .ZN(_10496_));
 NAND4_X1 _36275_ (.A1(_10266_),
    .A2(_10320_),
    .A3(_10496_),
    .A4(_10424_),
    .ZN(_10497_));
 NAND3_X1 _36276_ (.A1(\itlb.r_v_reg.N3 ),
    .A2(_10495_),
    .A3(_10497_),
    .ZN(_10498_));
 INV_X1 _36277_ (.A(\itlb.plru.encoder.lru_i [3]),
    .ZN(_10499_));
 OAI21_X1 _36278_ (.A(_10498_),
    .B1(_10479_),
    .B2(_10499_),
    .ZN(_06820_));
 OAI21_X1 _36279_ (.A(_00579_),
    .B1(_10486_),
    .B2(_10487_),
    .ZN(_10500_));
 OR2_X2 _36280_ (.A1(_10318_),
    .A2(_10319_),
    .ZN(_10501_));
 INV_X1 _36281_ (.A(_10424_),
    .ZN(_10502_));
 OAI211_X1 _36282_ (.A(_10266_),
    .B(_10373_),
    .C1(_10501_),
    .C2(_10502_),
    .ZN(_10503_));
 NAND3_X1 _36283_ (.A1(\itlb.r_v_reg.N3 ),
    .A2(_10500_),
    .A3(_10503_),
    .ZN(_10504_));
 OAI211_X1 _36284_ (.A(\itlb.plru.encoder.lru_i [4]),
    .B(_10206_),
    .C1(_10478_),
    .C2(_08480_),
    .ZN(_10505_));
 NAND2_X1 _36285_ (.A1(_10504_),
    .A2(_10505_),
    .ZN(_06821_));
 INV_X1 _36286_ (.A(_10487_),
    .ZN(_10506_));
 OAI21_X1 _36287_ (.A(_00580_),
    .B1(_10506_),
    .B2(_10266_),
    .ZN(_10507_));
 NAND3_X1 _36288_ (.A1(_10486_),
    .A2(_10496_),
    .A3(_10487_),
    .ZN(_10508_));
 NAND3_X1 _36289_ (.A1(_10507_),
    .A2(\itlb.r_v_reg.N3 ),
    .A3(_10508_),
    .ZN(_10509_));
 INV_X1 _36290_ (.A(\itlb.plru.encoder.lru_i [5]),
    .ZN(_10510_));
 OAI21_X1 _36291_ (.A(_10509_),
    .B1(_10479_),
    .B2(_10510_),
    .ZN(_06822_));
 OAI221_X2 _36292_ (.A(_10373_),
    .B1(_10483_),
    .B2(_10484_),
    .C1(_10501_),
    .C2(_10502_),
    .ZN(_10511_));
 OAI21_X1 _36293_ (.A(_00581_),
    .B1(_10487_),
    .B2(_10266_),
    .ZN(_10512_));
 NAND3_X1 _36294_ (.A1(\itlb.r_v_reg.N3 ),
    .A2(_10511_),
    .A3(_10512_),
    .ZN(_10513_));
 OAI211_X1 _36295_ (.A(\itlb.plru.encoder.lru_i [6]),
    .B(_10206_),
    .C1(_10478_),
    .C2(_08480_),
    .ZN(_10514_));
 NAND2_X1 _36296_ (.A1(_10513_),
    .A2(_10514_),
    .ZN(_06823_));
 BUF_X8 _36297_ (.A(_08551_),
    .Z(_10515_));
 AND2_X4 _36298_ (.A1(_08031_),
    .A2(_10206_),
    .ZN(_10516_));
 NAND3_X2 _36299_ (.A1(_10491_),
    .A2(\itlb.plru.encoder.lru_i [2]),
    .A3(\itlb.plru.encoder.lru_i [6]),
    .ZN(_10517_));
 OAI211_X4 _36300_ (.A(_10517_),
    .B(\itlb.plru.encoder.N1 ),
    .C1(\itlb.plru.encoder.lru_i [2]),
    .C2(_10510_),
    .ZN(_10518_));
 NAND2_X1 _36301_ (.A1(\itlb.plru.encoder.lru_i [1]),
    .A2(\itlb.plru.encoder.lru_i [4]),
    .ZN(_10519_));
 OAI211_X4 _36302_ (.A(_10519_),
    .B(_10480_),
    .C1(\itlb.plru.encoder.lru_i [1]),
    .C2(_10499_),
    .ZN(_10520_));
 NAND2_X1 _36303_ (.A1(_10480_),
    .A2(_00576_),
    .ZN(_10521_));
 NAND2_X1 _36304_ (.A1(\itlb.plru.encoder.N1 ),
    .A2(_00577_),
    .ZN(_10522_));
 NAND2_X2 _36305_ (.A1(_10521_),
    .A2(_10522_),
    .ZN(_10523_));
 AND4_X1 _36306_ (.A1(_10480_),
    .A2(_10518_),
    .A3(_10520_),
    .A4(_10523_),
    .ZN(_10524_));
 AND2_X1 _36307_ (.A1(_10516_),
    .A2(_10524_),
    .ZN(_10525_));
 BUF_X4 _36308_ (.A(_10525_),
    .Z(_10526_));
 BUF_X4 _36309_ (.A(_10526_),
    .Z(_10527_));
 MUX2_X1 _36310_ (.A(\itlb.vtag_cam.mem [162]),
    .B(_10515_),
    .S(_10527_),
    .Z(_06893_));
 BUF_X16 _36311_ (.A(_08555_),
    .Z(_10528_));
 MUX2_X1 _36312_ (.A(\itlb.vtag_cam.mem [163]),
    .B(_10528_),
    .S(_10527_),
    .Z(_06894_));
 BUF_X16 _36313_ (.A(_08558_),
    .Z(_10529_));
 MUX2_X1 _36314_ (.A(\itlb.vtag_cam.mem [164]),
    .B(_10529_),
    .S(_10527_),
    .Z(_06895_));
 BUF_X8 _36315_ (.A(_08561_),
    .Z(_10530_));
 MUX2_X1 _36316_ (.A(\itlb.vtag_cam.mem [165]),
    .B(_10530_),
    .S(_10527_),
    .Z(_06896_));
 BUF_X8 _36317_ (.A(_08564_),
    .Z(_10531_));
 MUX2_X1 _36318_ (.A(\itlb.vtag_cam.mem [166]),
    .B(_10531_),
    .S(_10527_),
    .Z(_06897_));
 BUF_X16 _36319_ (.A(_08567_),
    .Z(_10532_));
 MUX2_X1 _36320_ (.A(\itlb.vtag_cam.mem [167]),
    .B(_10532_),
    .S(_10527_),
    .Z(_06898_));
 BUF_X8 _36321_ (.A(_08571_),
    .Z(_10533_));
 MUX2_X1 _36322_ (.A(\itlb.vtag_cam.mem [168]),
    .B(_10533_),
    .S(_10527_),
    .Z(_06899_));
 BUF_X8 _36323_ (.A(_08575_),
    .Z(_10534_));
 MUX2_X1 _36324_ (.A(\itlb.vtag_cam.mem [169]),
    .B(_10534_),
    .S(_10527_),
    .Z(_06900_));
 BUF_X8 _36325_ (.A(_08578_),
    .Z(_10535_));
 MUX2_X1 _36326_ (.A(\itlb.vtag_cam.mem [170]),
    .B(_10535_),
    .S(_10527_),
    .Z(_06902_));
 BUF_X8 _36327_ (.A(_08581_),
    .Z(_10536_));
 BUF_X4 _36328_ (.A(_10526_),
    .Z(_10537_));
 MUX2_X1 _36329_ (.A(\itlb.vtag_cam.mem [171]),
    .B(_10536_),
    .S(_10537_),
    .Z(_06903_));
 BUF_X8 _36330_ (.A(_08584_),
    .Z(_10538_));
 MUX2_X1 _36331_ (.A(\itlb.vtag_cam.mem [172]),
    .B(_10538_),
    .S(_10537_),
    .Z(_06904_));
 BUF_X16 _36332_ (.A(_08588_),
    .Z(_10539_));
 MUX2_X1 _36333_ (.A(\itlb.vtag_cam.mem [173]),
    .B(_10539_),
    .S(_10537_),
    .Z(_06905_));
 BUF_X8 _36334_ (.A(_08591_),
    .Z(_10540_));
 MUX2_X1 _36335_ (.A(\itlb.vtag_cam.mem [174]),
    .B(_10540_),
    .S(_10537_),
    .Z(_06906_));
 BUF_X16 _36336_ (.A(_08594_),
    .Z(_10541_));
 MUX2_X1 _36337_ (.A(\itlb.vtag_cam.mem [175]),
    .B(_10541_),
    .S(_10537_),
    .Z(_06907_));
 BUF_X8 _36338_ (.A(_08597_),
    .Z(_10542_));
 MUX2_X1 _36339_ (.A(\itlb.vtag_cam.mem [176]),
    .B(_10542_),
    .S(_10537_),
    .Z(_06908_));
 BUF_X16 _36340_ (.A(_08600_),
    .Z(_10543_));
 MUX2_X1 _36341_ (.A(\itlb.vtag_cam.mem [177]),
    .B(_10543_),
    .S(_10537_),
    .Z(_06909_));
 BUF_X16 _36342_ (.A(_08604_),
    .Z(_10544_));
 MUX2_X1 _36343_ (.A(\itlb.vtag_cam.mem [178]),
    .B(_10544_),
    .S(_10537_),
    .Z(_06910_));
 BUF_X16 _36344_ (.A(_08608_),
    .Z(_10545_));
 MUX2_X1 _36345_ (.A(\itlb.vtag_cam.mem [179]),
    .B(_10545_),
    .S(_10537_),
    .Z(_06911_));
 BUF_X8 _36346_ (.A(_08611_),
    .Z(_10546_));
 MUX2_X1 _36347_ (.A(\itlb.vtag_cam.mem [180]),
    .B(_10546_),
    .S(_10537_),
    .Z(_06913_));
 BUF_X16 _36348_ (.A(_08614_),
    .Z(_10547_));
 MUX2_X1 _36349_ (.A(\itlb.vtag_cam.mem [181]),
    .B(_10547_),
    .S(_10526_),
    .Z(_06914_));
 BUF_X8 _36350_ (.A(_08617_),
    .Z(_10548_));
 MUX2_X1 _36351_ (.A(\itlb.vtag_cam.mem [182]),
    .B(_10548_),
    .S(_10526_),
    .Z(_06915_));
 BUF_X8 _36352_ (.A(_08620_),
    .Z(_10549_));
 MUX2_X1 _36353_ (.A(\itlb.vtag_cam.mem [183]),
    .B(_10549_),
    .S(_10526_),
    .Z(_06916_));
 BUF_X16 _36354_ (.A(_08623_),
    .Z(_10550_));
 MUX2_X1 _36355_ (.A(\itlb.vtag_cam.mem [184]),
    .B(_10550_),
    .S(_10526_),
    .Z(_06917_));
 BUF_X8 _36356_ (.A(_08626_),
    .Z(_10551_));
 MUX2_X1 _36357_ (.A(\itlb.vtag_cam.mem [185]),
    .B(_10551_),
    .S(_10526_),
    .Z(_06918_));
 BUF_X8 _36358_ (.A(_08629_),
    .Z(_10552_));
 MUX2_X1 _36359_ (.A(\itlb.vtag_cam.mem [186]),
    .B(_10552_),
    .S(_10526_),
    .Z(_06919_));
 BUF_X16 _36360_ (.A(_08632_),
    .Z(_10553_));
 MUX2_X1 _36361_ (.A(\itlb.vtag_cam.mem [187]),
    .B(_10553_),
    .S(_10526_),
    .Z(_06920_));
 BUF_X16 _36362_ (.A(_08635_),
    .Z(_10554_));
 MUX2_X1 _36363_ (.A(\itlb.vtag_cam.mem [188]),
    .B(_10554_),
    .S(_10526_),
    .Z(_06921_));
 INV_X1 _36364_ (.A(_00582_),
    .ZN(_10555_));
 NAND2_X4 _36365_ (.A1(_10516_),
    .A2(_10555_),
    .ZN(_10556_));
 NAND2_X2 _36366_ (.A1(_10518_),
    .A2(_10520_),
    .ZN(_10557_));
 INV_X2 _36367_ (.A(_10523_),
    .ZN(_10558_));
 NAND2_X4 _36368_ (.A1(_10557_),
    .A2(_10558_),
    .ZN(_10559_));
 NOR2_X4 _36369_ (.A1(_10556_),
    .A2(_10559_),
    .ZN(_10560_));
 BUF_X4 _36370_ (.A(_10560_),
    .Z(_10561_));
 MUX2_X1 _36371_ (.A(\itlb.vtag_cam.mem [27]),
    .B(_10515_),
    .S(_10561_),
    .Z(_06959_));
 MUX2_X1 _36372_ (.A(\itlb.vtag_cam.mem [28]),
    .B(_10528_),
    .S(_10561_),
    .Z(_06960_));
 MUX2_X1 _36373_ (.A(\itlb.vtag_cam.mem [29]),
    .B(_10529_),
    .S(_10561_),
    .Z(_06961_));
 MUX2_X1 _36374_ (.A(\itlb.vtag_cam.mem [30]),
    .B(_10530_),
    .S(_10561_),
    .Z(_06963_));
 MUX2_X1 _36375_ (.A(\itlb.vtag_cam.mem [31]),
    .B(_10531_),
    .S(_10561_),
    .Z(_06964_));
 MUX2_X1 _36376_ (.A(\itlb.vtag_cam.mem [32]),
    .B(_10532_),
    .S(_10561_),
    .Z(_06965_));
 MUX2_X1 _36377_ (.A(\itlb.vtag_cam.mem [33]),
    .B(_10533_),
    .S(_10561_),
    .Z(_06966_));
 MUX2_X1 _36378_ (.A(\itlb.vtag_cam.mem [34]),
    .B(_10534_),
    .S(_10561_),
    .Z(_06967_));
 MUX2_X1 _36379_ (.A(\itlb.vtag_cam.mem [35]),
    .B(_10535_),
    .S(_10561_),
    .Z(_06968_));
 MUX2_X1 _36380_ (.A(\itlb.vtag_cam.mem [36]),
    .B(_10536_),
    .S(_10561_),
    .Z(_06969_));
 BUF_X8 _36381_ (.A(_10560_),
    .Z(_10562_));
 MUX2_X1 _36382_ (.A(\itlb.vtag_cam.mem [37]),
    .B(_10538_),
    .S(_10562_),
    .Z(_06970_));
 MUX2_X1 _36383_ (.A(\itlb.vtag_cam.mem [38]),
    .B(_10539_),
    .S(_10562_),
    .Z(_06971_));
 MUX2_X1 _36384_ (.A(\itlb.vtag_cam.mem [39]),
    .B(_10540_),
    .S(_10562_),
    .Z(_06972_));
 MUX2_X1 _36385_ (.A(\itlb.vtag_cam.mem [40]),
    .B(_10541_),
    .S(_10562_),
    .Z(_06974_));
 MUX2_X1 _36386_ (.A(\itlb.vtag_cam.mem [41]),
    .B(_10542_),
    .S(_10562_),
    .Z(_06975_));
 MUX2_X1 _36387_ (.A(\itlb.vtag_cam.mem [42]),
    .B(_10543_),
    .S(_10562_),
    .Z(_06976_));
 MUX2_X1 _36388_ (.A(\itlb.vtag_cam.mem [43]),
    .B(_10544_),
    .S(_10562_),
    .Z(_06977_));
 MUX2_X1 _36389_ (.A(\itlb.vtag_cam.mem [44]),
    .B(_10545_),
    .S(_10562_),
    .Z(_06978_));
 MUX2_X1 _36390_ (.A(\itlb.vtag_cam.mem [45]),
    .B(_10546_),
    .S(_10562_),
    .Z(_06979_));
 MUX2_X1 _36391_ (.A(\itlb.vtag_cam.mem [46]),
    .B(_10547_),
    .S(_10562_),
    .Z(_06980_));
 MUX2_X1 _36392_ (.A(\itlb.vtag_cam.mem [47]),
    .B(_10548_),
    .S(_10560_),
    .Z(_06981_));
 MUX2_X1 _36393_ (.A(\itlb.vtag_cam.mem [48]),
    .B(_10549_),
    .S(_10560_),
    .Z(_06982_));
 MUX2_X1 _36394_ (.A(\itlb.vtag_cam.mem [49]),
    .B(_10550_),
    .S(_10560_),
    .Z(_06983_));
 MUX2_X1 _36395_ (.A(\itlb.vtag_cam.mem [50]),
    .B(_10551_),
    .S(_10560_),
    .Z(_06985_));
 MUX2_X1 _36396_ (.A(\itlb.vtag_cam.mem [51]),
    .B(_10552_),
    .S(_10560_),
    .Z(_06986_));
 MUX2_X1 _36397_ (.A(\itlb.vtag_cam.mem [52]),
    .B(_10553_),
    .S(_10560_),
    .Z(_06987_));
 MUX2_X1 _36398_ (.A(\itlb.vtag_cam.mem [53]),
    .B(_10554_),
    .S(_10560_),
    .Z(_06988_));
 BUF_X32 _36399_ (.A(_08551_),
    .Z(_10563_));
 NAND2_X4 _36400_ (.A1(_10516_),
    .A2(_10480_),
    .ZN(_10564_));
 NAND2_X4 _36401_ (.A1(_10557_),
    .A2(_10523_),
    .ZN(_10565_));
 OR2_X1 _36402_ (.A1(_10564_),
    .A2(_10565_),
    .ZN(_10566_));
 BUF_X4 _36403_ (.A(_10566_),
    .Z(_10567_));
 BUF_X4 _36404_ (.A(_10567_),
    .Z(_10568_));
 MUX2_X1 _36405_ (.A(_10563_),
    .B(\itlb.vtag_cam.mem [189]),
    .S(_10568_),
    .Z(_06922_));
 BUF_X16 _36406_ (.A(_08555_),
    .Z(_10569_));
 MUX2_X1 _36407_ (.A(_10569_),
    .B(\itlb.vtag_cam.mem [190]),
    .S(_10568_),
    .Z(_06924_));
 BUF_X16 _36408_ (.A(_08558_),
    .Z(_10570_));
 MUX2_X1 _36409_ (.A(_10570_),
    .B(\itlb.vtag_cam.mem [191]),
    .S(_10568_),
    .Z(_06925_));
 BUF_X16 _36410_ (.A(_08561_),
    .Z(_10571_));
 MUX2_X1 _36411_ (.A(_10571_),
    .B(\itlb.vtag_cam.mem [192]),
    .S(_10568_),
    .Z(_06926_));
 BUF_X32 _36412_ (.A(_08564_),
    .Z(_10572_));
 MUX2_X1 _36413_ (.A(_10572_),
    .B(\itlb.vtag_cam.mem [193]),
    .S(_10568_),
    .Z(_06927_));
 BUF_X16 _36414_ (.A(_08567_),
    .Z(_10573_));
 BUF_X4 _36415_ (.A(_10567_),
    .Z(_10574_));
 MUX2_X1 _36416_ (.A(_10573_),
    .B(\itlb.vtag_cam.mem [194]),
    .S(_10574_),
    .Z(_06928_));
 NOR3_X1 _36417_ (.A1(_10564_),
    .A2(_08571_),
    .A3(_10565_),
    .ZN(_10575_));
 AOI21_X1 _36418_ (.A(_10575_),
    .B1(_10448_),
    .B2(_10568_),
    .ZN(_06929_));
 BUF_X8 _36419_ (.A(_08575_),
    .Z(_10576_));
 MUX2_X1 _36420_ (.A(_10576_),
    .B(\itlb.vtag_cam.mem [196]),
    .S(_10574_),
    .Z(_06930_));
 BUF_X8 _36421_ (.A(_08578_),
    .Z(_10577_));
 MUX2_X1 _36422_ (.A(_10577_),
    .B(\itlb.vtag_cam.mem [197]),
    .S(_10574_),
    .Z(_06931_));
 BUF_X16 _36423_ (.A(_08581_),
    .Z(_10578_));
 MUX2_X1 _36424_ (.A(_10578_),
    .B(\itlb.vtag_cam.mem [198]),
    .S(_10574_),
    .Z(_06932_));
 BUF_X16 _36425_ (.A(_08584_),
    .Z(_10579_));
 MUX2_X1 _36426_ (.A(_10579_),
    .B(\itlb.vtag_cam.mem [199]),
    .S(_10574_),
    .Z(_06933_));
 BUF_X16 _36427_ (.A(_08588_),
    .Z(_10580_));
 MUX2_X1 _36428_ (.A(_10580_),
    .B(\itlb.vtag_cam.mem [200]),
    .S(_10574_),
    .Z(_06936_));
 NOR3_X1 _36429_ (.A1(_10564_),
    .A2(_08591_),
    .A3(_10565_),
    .ZN(_10581_));
 AOI21_X1 _36430_ (.A(_10581_),
    .B1(_10456_),
    .B2(_10568_),
    .ZN(_06937_));
 BUF_X8 _36431_ (.A(_08594_),
    .Z(_10582_));
 MUX2_X1 _36432_ (.A(_10582_),
    .B(\itlb.vtag_cam.mem [202]),
    .S(_10574_),
    .Z(_06938_));
 BUF_X16 _36433_ (.A(_08597_),
    .Z(_10583_));
 MUX2_X1 _36434_ (.A(_10583_),
    .B(\itlb.vtag_cam.mem [203]),
    .S(_10574_),
    .Z(_06939_));
 BUF_X16 _36435_ (.A(_08600_),
    .Z(_10584_));
 MUX2_X1 _36436_ (.A(_10584_),
    .B(\itlb.vtag_cam.mem [204]),
    .S(_10574_),
    .Z(_06940_));
 BUF_X16 _36437_ (.A(_08604_),
    .Z(_10585_));
 MUX2_X1 _36438_ (.A(_10585_),
    .B(\itlb.vtag_cam.mem [205]),
    .S(_10574_),
    .Z(_06941_));
 BUF_X4 _36439_ (.A(_08608_),
    .Z(_10586_));
 MUX2_X1 _36440_ (.A(_10586_),
    .B(\itlb.vtag_cam.mem [206]),
    .S(_10567_),
    .Z(_06942_));
 BUF_X16 _36441_ (.A(_08611_),
    .Z(_10587_));
 MUX2_X1 _36442_ (.A(_10587_),
    .B(\itlb.vtag_cam.mem [207]),
    .S(_10567_),
    .Z(_06943_));
 BUF_X16 _36443_ (.A(_08614_),
    .Z(_10588_));
 MUX2_X1 _36444_ (.A(_10588_),
    .B(\itlb.vtag_cam.mem [208]),
    .S(_10567_),
    .Z(_06944_));
 NOR3_X1 _36445_ (.A1(_10564_),
    .A2(_08617_),
    .A3(_10565_),
    .ZN(_10589_));
 AOI21_X1 _36446_ (.A(_10589_),
    .B1(_10435_),
    .B2(_10568_),
    .ZN(_06945_));
 NOR3_X1 _36447_ (.A1(_10564_),
    .A2(_08620_),
    .A3(_10565_),
    .ZN(_10590_));
 AOI21_X1 _36448_ (.A(_10590_),
    .B1(_10463_),
    .B2(_10568_),
    .ZN(_06947_));
 BUF_X16 _36449_ (.A(_08623_),
    .Z(_10591_));
 MUX2_X1 _36450_ (.A(_10591_),
    .B(\itlb.vtag_cam.mem [211]),
    .S(_10567_),
    .Z(_06948_));
 BUF_X4 _36451_ (.A(_08626_),
    .Z(_10592_));
 MUX2_X1 _36452_ (.A(_10592_),
    .B(\itlb.vtag_cam.mem [212]),
    .S(_10567_),
    .Z(_06949_));
 BUF_X16 _36453_ (.A(_08629_),
    .Z(_10593_));
 MUX2_X1 _36454_ (.A(_10593_),
    .B(\itlb.vtag_cam.mem [213]),
    .S(_10567_),
    .Z(_06950_));
 NOR3_X1 _36455_ (.A1(_10564_),
    .A2(_08632_),
    .A3(_10565_),
    .ZN(_10594_));
 AOI21_X1 _36456_ (.A(_10594_),
    .B1(_10451_),
    .B2(_10568_),
    .ZN(_06951_));
 BUF_X16 _36457_ (.A(_08635_),
    .Z(_10595_));
 MUX2_X1 _36458_ (.A(_10595_),
    .B(\itlb.vtag_cam.mem [215]),
    .S(_10567_),
    .Z(_06952_));
 OR2_X2 _36459_ (.A1(_10564_),
    .A2(_10559_),
    .ZN(_10596_));
 BUF_X4 _36460_ (.A(_10596_),
    .Z(_10597_));
 BUF_X4 _36461_ (.A(_10597_),
    .Z(_10598_));
 MUX2_X1 _36462_ (.A(_10563_),
    .B(\itlb.vtag_cam.mem [135]),
    .S(_10598_),
    .Z(_06863_));
 MUX2_X1 _36463_ (.A(_10569_),
    .B(\itlb.vtag_cam.mem [136]),
    .S(_10598_),
    .Z(_06864_));
 MUX2_X1 _36464_ (.A(_10570_),
    .B(\itlb.vtag_cam.mem [137]),
    .S(_10598_),
    .Z(_06865_));
 MUX2_X1 _36465_ (.A(_10571_),
    .B(\itlb.vtag_cam.mem [138]),
    .S(_10598_),
    .Z(_06866_));
 MUX2_X1 _36466_ (.A(_10572_),
    .B(\itlb.vtag_cam.mem [139]),
    .S(_10598_),
    .Z(_06867_));
 BUF_X16 _36467_ (.A(_08567_),
    .Z(_10599_));
 MUX2_X1 _36468_ (.A(_10599_),
    .B(\itlb.vtag_cam.mem [140]),
    .S(_10598_),
    .Z(_06869_));
 BUF_X16 _36469_ (.A(_08571_),
    .Z(_10600_));
 MUX2_X1 _36470_ (.A(_10600_),
    .B(\itlb.vtag_cam.mem [141]),
    .S(_10598_),
    .Z(_06870_));
 MUX2_X1 _36471_ (.A(_08575_),
    .B(\itlb.vtag_cam.mem [142]),
    .S(_10598_),
    .Z(_06871_));
 MUX2_X1 _36472_ (.A(_10577_),
    .B(\itlb.vtag_cam.mem [143]),
    .S(_10598_),
    .Z(_06872_));
 MUX2_X1 _36473_ (.A(_10578_),
    .B(\itlb.vtag_cam.mem [144]),
    .S(_10598_),
    .Z(_06873_));
 BUF_X4 _36474_ (.A(_10597_),
    .Z(_10601_));
 MUX2_X1 _36475_ (.A(_10579_),
    .B(\itlb.vtag_cam.mem [145]),
    .S(_10601_),
    .Z(_06874_));
 MUX2_X1 _36476_ (.A(_10580_),
    .B(\itlb.vtag_cam.mem [146]),
    .S(_10601_),
    .Z(_06875_));
 BUF_X16 _36477_ (.A(_08591_),
    .Z(_10602_));
 MUX2_X1 _36478_ (.A(_10602_),
    .B(\itlb.vtag_cam.mem [147]),
    .S(_10601_),
    .Z(_06876_));
 MUX2_X1 _36479_ (.A(_10582_),
    .B(\itlb.vtag_cam.mem [148]),
    .S(_10601_),
    .Z(_06877_));
 MUX2_X1 _36480_ (.A(_10583_),
    .B(\itlb.vtag_cam.mem [149]),
    .S(_10601_),
    .Z(_06878_));
 MUX2_X1 _36481_ (.A(_10584_),
    .B(\itlb.vtag_cam.mem [150]),
    .S(_10601_),
    .Z(_06880_));
 MUX2_X1 _36482_ (.A(_10585_),
    .B(\itlb.vtag_cam.mem [151]),
    .S(_10601_),
    .Z(_06881_));
 MUX2_X1 _36483_ (.A(_10586_),
    .B(\itlb.vtag_cam.mem [152]),
    .S(_10601_),
    .Z(_06882_));
 MUX2_X1 _36484_ (.A(_10587_),
    .B(\itlb.vtag_cam.mem [153]),
    .S(_10601_),
    .Z(_06883_));
 MUX2_X1 _36485_ (.A(_10588_),
    .B(\itlb.vtag_cam.mem [154]),
    .S(_10601_),
    .Z(_06884_));
 BUF_X16 _36486_ (.A(_08617_),
    .Z(_10603_));
 MUX2_X1 _36487_ (.A(_10603_),
    .B(\itlb.vtag_cam.mem [155]),
    .S(_10597_),
    .Z(_06885_));
 BUF_X16 _36488_ (.A(_08620_),
    .Z(_10604_));
 MUX2_X1 _36489_ (.A(_10604_),
    .B(\itlb.vtag_cam.mem [156]),
    .S(_10597_),
    .Z(_06886_));
 MUX2_X1 _36490_ (.A(_10591_),
    .B(\itlb.vtag_cam.mem [157]),
    .S(_10597_),
    .Z(_06887_));
 MUX2_X1 _36491_ (.A(_10592_),
    .B(\itlb.vtag_cam.mem [158]),
    .S(_10597_),
    .Z(_06888_));
 MUX2_X1 _36492_ (.A(_10593_),
    .B(\itlb.vtag_cam.mem [159]),
    .S(_10597_),
    .Z(_06889_));
 BUF_X16 _36493_ (.A(_08632_),
    .Z(_10605_));
 MUX2_X1 _36494_ (.A(_10605_),
    .B(\itlb.vtag_cam.mem [160]),
    .S(_10597_),
    .Z(_06891_));
 MUX2_X1 _36495_ (.A(_10595_),
    .B(\itlb.vtag_cam.mem [161]),
    .S(_10597_),
    .Z(_06892_));
 AND4_X1 _36496_ (.A1(_10480_),
    .A2(_10518_),
    .A3(_10520_),
    .A4(_10558_),
    .ZN(_10606_));
 AND2_X1 _36497_ (.A1(_10516_),
    .A2(_10606_),
    .ZN(_10607_));
 BUF_X4 _36498_ (.A(_10607_),
    .Z(_10608_));
 BUF_X4 _36499_ (.A(_10608_),
    .Z(_10609_));
 MUX2_X1 _36500_ (.A(\itlb.vtag_cam.mem [108]),
    .B(_10515_),
    .S(_10609_),
    .Z(_06833_));
 MUX2_X1 _36501_ (.A(\itlb.vtag_cam.mem [109]),
    .B(_10528_),
    .S(_10609_),
    .Z(_06834_));
 MUX2_X1 _36502_ (.A(\itlb.vtag_cam.mem [110]),
    .B(_10529_),
    .S(_10609_),
    .Z(_06836_));
 MUX2_X1 _36503_ (.A(\itlb.vtag_cam.mem [111]),
    .B(_10530_),
    .S(_10609_),
    .Z(_06837_));
 MUX2_X1 _36504_ (.A(\itlb.vtag_cam.mem [112]),
    .B(_10531_),
    .S(_10609_),
    .Z(_06838_));
 MUX2_X1 _36505_ (.A(\itlb.vtag_cam.mem [113]),
    .B(_10532_),
    .S(_10609_),
    .Z(_06839_));
 MUX2_X1 _36506_ (.A(\itlb.vtag_cam.mem [114]),
    .B(_10533_),
    .S(_10609_),
    .Z(_06840_));
 MUX2_X1 _36507_ (.A(\itlb.vtag_cam.mem [115]),
    .B(_10534_),
    .S(_10609_),
    .Z(_06841_));
 MUX2_X1 _36508_ (.A(\itlb.vtag_cam.mem [116]),
    .B(_10535_),
    .S(_10609_),
    .Z(_06842_));
 BUF_X4 _36509_ (.A(_10608_),
    .Z(_10610_));
 MUX2_X1 _36510_ (.A(\itlb.vtag_cam.mem [117]),
    .B(_10536_),
    .S(_10610_),
    .Z(_06843_));
 MUX2_X1 _36511_ (.A(\itlb.vtag_cam.mem [118]),
    .B(_10538_),
    .S(_10610_),
    .Z(_06844_));
 MUX2_X1 _36512_ (.A(\itlb.vtag_cam.mem [119]),
    .B(_10539_),
    .S(_10610_),
    .Z(_06845_));
 MUX2_X1 _36513_ (.A(\itlb.vtag_cam.mem [120]),
    .B(_10540_),
    .S(_10610_),
    .Z(_06847_));
 MUX2_X1 _36514_ (.A(\itlb.vtag_cam.mem [121]),
    .B(_10541_),
    .S(_10610_),
    .Z(_06848_));
 MUX2_X1 _36515_ (.A(\itlb.vtag_cam.mem [122]),
    .B(_10542_),
    .S(_10610_),
    .Z(_06849_));
 MUX2_X1 _36516_ (.A(\itlb.vtag_cam.mem [123]),
    .B(_10543_),
    .S(_10610_),
    .Z(_06850_));
 MUX2_X1 _36517_ (.A(\itlb.vtag_cam.mem [124]),
    .B(_10544_),
    .S(_10610_),
    .Z(_06851_));
 MUX2_X1 _36518_ (.A(\itlb.vtag_cam.mem [125]),
    .B(_10545_),
    .S(_10610_),
    .Z(_06852_));
 MUX2_X1 _36519_ (.A(\itlb.vtag_cam.mem [126]),
    .B(_10546_),
    .S(_10610_),
    .Z(_06853_));
 MUX2_X1 _36520_ (.A(\itlb.vtag_cam.mem [127]),
    .B(_10547_),
    .S(_10608_),
    .Z(_06854_));
 MUX2_X1 _36521_ (.A(\itlb.vtag_cam.mem [128]),
    .B(_10548_),
    .S(_10608_),
    .Z(_06855_));
 MUX2_X1 _36522_ (.A(\itlb.vtag_cam.mem [129]),
    .B(_10549_),
    .S(_10608_),
    .Z(_06856_));
 MUX2_X1 _36523_ (.A(\itlb.vtag_cam.mem [130]),
    .B(_10550_),
    .S(_10608_),
    .Z(_06858_));
 MUX2_X1 _36524_ (.A(\itlb.vtag_cam.mem [131]),
    .B(_10551_),
    .S(_10608_),
    .Z(_06859_));
 MUX2_X1 _36525_ (.A(\itlb.vtag_cam.mem [132]),
    .B(_10552_),
    .S(_10608_),
    .Z(_06860_));
 MUX2_X1 _36526_ (.A(\itlb.vtag_cam.mem [133]),
    .B(_10553_),
    .S(_10608_),
    .Z(_06861_));
 MUX2_X1 _36527_ (.A(\itlb.vtag_cam.mem [134]),
    .B(_10554_),
    .S(_10608_),
    .Z(_06862_));
 AOI221_X4 _36528_ (.A(_00582_),
    .B1(_10522_),
    .B2(_10521_),
    .C1(_10518_),
    .C2(_10520_),
    .ZN(_10611_));
 NAND2_X4 _36529_ (.A1(_10516_),
    .A2(_10611_),
    .ZN(_10612_));
 BUF_X4 _36530_ (.A(_10612_),
    .Z(_10613_));
 MUX2_X1 _36531_ (.A(_10563_),
    .B(\itlb.vtag_cam.mem [81]),
    .S(_10613_),
    .Z(_07019_));
 MUX2_X1 _36532_ (.A(_10569_),
    .B(\itlb.vtag_cam.mem [82]),
    .S(_10613_),
    .Z(_07020_));
 MUX2_X1 _36533_ (.A(_10570_),
    .B(\itlb.vtag_cam.mem [83]),
    .S(_10613_),
    .Z(_07021_));
 MUX2_X1 _36534_ (.A(_10571_),
    .B(\itlb.vtag_cam.mem [84]),
    .S(_10613_),
    .Z(_07022_));
 MUX2_X1 _36535_ (.A(_10572_),
    .B(\itlb.vtag_cam.mem [85]),
    .S(_10613_),
    .Z(_07023_));
 MUX2_X1 _36536_ (.A(_10599_),
    .B(\itlb.vtag_cam.mem [86]),
    .S(_10613_),
    .Z(_07024_));
 MUX2_X1 _36537_ (.A(_10600_),
    .B(\itlb.vtag_cam.mem [87]),
    .S(_10613_),
    .Z(_07025_));
 MUX2_X1 _36538_ (.A(_08575_),
    .B(\itlb.vtag_cam.mem [88]),
    .S(_10613_),
    .Z(_07026_));
 BUF_X32 _36539_ (.A(_08578_),
    .Z(_10614_));
 MUX2_X1 _36540_ (.A(_10614_),
    .B(\itlb.vtag_cam.mem [89]),
    .S(_10613_),
    .Z(_07027_));
 BUF_X4 _36541_ (.A(_10612_),
    .Z(_10615_));
 MUX2_X1 _36542_ (.A(_10578_),
    .B(\itlb.vtag_cam.mem [90]),
    .S(_10615_),
    .Z(_07029_));
 MUX2_X1 _36543_ (.A(_10579_),
    .B(\itlb.vtag_cam.mem [91]),
    .S(_10615_),
    .Z(_07030_));
 MUX2_X1 _36544_ (.A(_10580_),
    .B(\itlb.vtag_cam.mem [92]),
    .S(_10615_),
    .Z(_07031_));
 MUX2_X1 _36545_ (.A(_10602_),
    .B(\itlb.vtag_cam.mem [93]),
    .S(_10615_),
    .Z(_07032_));
 MUX2_X1 _36546_ (.A(_10582_),
    .B(\itlb.vtag_cam.mem [94]),
    .S(_10615_),
    .Z(_07033_));
 MUX2_X1 _36547_ (.A(_10583_),
    .B(\itlb.vtag_cam.mem [95]),
    .S(_10615_),
    .Z(_07034_));
 MUX2_X1 _36548_ (.A(_10584_),
    .B(\itlb.vtag_cam.mem [96]),
    .S(_10615_),
    .Z(_07035_));
 MUX2_X1 _36549_ (.A(_10585_),
    .B(\itlb.vtag_cam.mem [97]),
    .S(_10615_),
    .Z(_07036_));
 BUF_X32 _36550_ (.A(_08608_),
    .Z(_10616_));
 MUX2_X1 _36551_ (.A(_10616_),
    .B(\itlb.vtag_cam.mem [98]),
    .S(_10615_),
    .Z(_07037_));
 MUX2_X1 _36552_ (.A(_10587_),
    .B(\itlb.vtag_cam.mem [99]),
    .S(_10615_),
    .Z(_07038_));
 MUX2_X1 _36553_ (.A(_10588_),
    .B(\itlb.vtag_cam.mem [100]),
    .S(_10612_),
    .Z(_06825_));
 MUX2_X1 _36554_ (.A(_10603_),
    .B(\itlb.vtag_cam.mem [101]),
    .S(_10612_),
    .Z(_06826_));
 MUX2_X1 _36555_ (.A(_10604_),
    .B(\itlb.vtag_cam.mem [102]),
    .S(_10612_),
    .Z(_06827_));
 MUX2_X1 _36556_ (.A(_10591_),
    .B(\itlb.vtag_cam.mem [103]),
    .S(_10612_),
    .Z(_06828_));
 MUX2_X1 _36557_ (.A(_08626_),
    .B(\itlb.vtag_cam.mem [104]),
    .S(_10612_),
    .Z(_06829_));
 MUX2_X1 _36558_ (.A(_10593_),
    .B(\itlb.vtag_cam.mem [105]),
    .S(_10612_),
    .Z(_06830_));
 MUX2_X1 _36559_ (.A(_10605_),
    .B(\itlb.vtag_cam.mem [106]),
    .S(_10612_),
    .Z(_06831_));
 MUX2_X1 _36560_ (.A(_10595_),
    .B(\itlb.vtag_cam.mem [107]),
    .S(_10612_),
    .Z(_06832_));
 AND4_X1 _36561_ (.A1(_10555_),
    .A2(_10518_),
    .A3(_10520_),
    .A4(_10523_),
    .ZN(_10617_));
 AND2_X1 _36562_ (.A1(_10516_),
    .A2(_10617_),
    .ZN(_10618_));
 BUF_X8 _36563_ (.A(_10618_),
    .Z(_10619_));
 BUF_X4 _36564_ (.A(_10619_),
    .Z(_10620_));
 MUX2_X1 _36565_ (.A(\itlb.vtag_cam.mem [54]),
    .B(_10515_),
    .S(_10620_),
    .Z(_06989_));
 MUX2_X1 _36566_ (.A(\itlb.vtag_cam.mem [55]),
    .B(_10528_),
    .S(_10620_),
    .Z(_06990_));
 MUX2_X1 _36567_ (.A(\itlb.vtag_cam.mem [56]),
    .B(_10529_),
    .S(_10620_),
    .Z(_06991_));
 MUX2_X1 _36568_ (.A(\itlb.vtag_cam.mem [57]),
    .B(_10530_),
    .S(_10620_),
    .Z(_06992_));
 MUX2_X1 _36569_ (.A(\itlb.vtag_cam.mem [58]),
    .B(_10531_),
    .S(_10620_),
    .Z(_06993_));
 MUX2_X1 _36570_ (.A(\itlb.vtag_cam.mem [59]),
    .B(_10532_),
    .S(_10620_),
    .Z(_06994_));
 MUX2_X1 _36571_ (.A(\itlb.vtag_cam.mem [60]),
    .B(_10533_),
    .S(_10620_),
    .Z(_06996_));
 MUX2_X1 _36572_ (.A(\itlb.vtag_cam.mem [61]),
    .B(_10534_),
    .S(_10620_),
    .Z(_06997_));
 MUX2_X1 _36573_ (.A(\itlb.vtag_cam.mem [62]),
    .B(_10535_),
    .S(_10620_),
    .Z(_06998_));
 BUF_X4 _36574_ (.A(_10619_),
    .Z(_10621_));
 MUX2_X1 _36575_ (.A(\itlb.vtag_cam.mem [63]),
    .B(_10536_),
    .S(_10621_),
    .Z(_06999_));
 MUX2_X1 _36576_ (.A(\itlb.vtag_cam.mem [64]),
    .B(_10538_),
    .S(_10621_),
    .Z(_07000_));
 MUX2_X1 _36577_ (.A(\itlb.vtag_cam.mem [65]),
    .B(_10539_),
    .S(_10621_),
    .Z(_07001_));
 MUX2_X1 _36578_ (.A(\itlb.vtag_cam.mem [66]),
    .B(_10540_),
    .S(_10621_),
    .Z(_07002_));
 MUX2_X1 _36579_ (.A(\itlb.vtag_cam.mem [67]),
    .B(_10541_),
    .S(_10621_),
    .Z(_07003_));
 MUX2_X1 _36580_ (.A(\itlb.vtag_cam.mem [68]),
    .B(_10542_),
    .S(_10621_),
    .Z(_07004_));
 MUX2_X1 _36581_ (.A(\itlb.vtag_cam.mem [69]),
    .B(_10543_),
    .S(_10621_),
    .Z(_07005_));
 MUX2_X1 _36582_ (.A(\itlb.vtag_cam.mem [70]),
    .B(_10544_),
    .S(_10621_),
    .Z(_07007_));
 MUX2_X1 _36583_ (.A(\itlb.vtag_cam.mem [71]),
    .B(_10545_),
    .S(_10621_),
    .Z(_07008_));
 MUX2_X1 _36584_ (.A(\itlb.vtag_cam.mem [72]),
    .B(_10546_),
    .S(_10621_),
    .Z(_07009_));
 MUX2_X1 _36585_ (.A(\itlb.vtag_cam.mem [73]),
    .B(_10547_),
    .S(_10619_),
    .Z(_07010_));
 MUX2_X1 _36586_ (.A(\itlb.vtag_cam.mem [74]),
    .B(_10548_),
    .S(_10619_),
    .Z(_07011_));
 MUX2_X1 _36587_ (.A(\itlb.vtag_cam.mem [75]),
    .B(_10549_),
    .S(_10619_),
    .Z(_07012_));
 MUX2_X1 _36588_ (.A(\itlb.vtag_cam.mem [76]),
    .B(_10550_),
    .S(_10619_),
    .Z(_07013_));
 MUX2_X1 _36589_ (.A(\itlb.vtag_cam.mem [77]),
    .B(_10551_),
    .S(_10619_),
    .Z(_07014_));
 MUX2_X1 _36590_ (.A(\itlb.vtag_cam.mem [78]),
    .B(_10552_),
    .S(_10619_),
    .Z(_07015_));
 MUX2_X1 _36591_ (.A(\itlb.vtag_cam.mem [79]),
    .B(_10553_),
    .S(_10619_),
    .Z(_07016_));
 MUX2_X1 _36592_ (.A(\itlb.vtag_cam.mem [80]),
    .B(_10554_),
    .S(_10619_),
    .Z(_07018_));
 AND4_X1 _36593_ (.A1(_10555_),
    .A2(_10518_),
    .A3(_10520_),
    .A4(_10558_),
    .ZN(_10622_));
 AND2_X1 _36594_ (.A1(_10516_),
    .A2(_10622_),
    .ZN(_10623_));
 BUF_X8 _36595_ (.A(_10623_),
    .Z(_10624_));
 BUF_X8 _36596_ (.A(_10624_),
    .Z(_10625_));
 MUX2_X1 _36597_ (.A(\itlb.vtag_cam.mem [0]),
    .B(_10515_),
    .S(_10625_),
    .Z(_06824_));
 MUX2_X1 _36598_ (.A(\itlb.vtag_cam.mem [1]),
    .B(_10528_),
    .S(_10625_),
    .Z(_06935_));
 MUX2_X1 _36599_ (.A(\itlb.vtag_cam.mem [2]),
    .B(_10529_),
    .S(_10625_),
    .Z(_06962_));
 MUX2_X1 _36600_ (.A(\itlb.vtag_cam.mem [3]),
    .B(_10530_),
    .S(_10625_),
    .Z(_06973_));
 MUX2_X1 _36601_ (.A(\itlb.vtag_cam.mem [4]),
    .B(_10531_),
    .S(_10625_),
    .Z(_06984_));
 MUX2_X1 _36602_ (.A(\itlb.vtag_cam.mem [5]),
    .B(_10532_),
    .S(_10625_),
    .Z(_06995_));
 MUX2_X1 _36603_ (.A(\itlb.vtag_cam.mem [6]),
    .B(_10533_),
    .S(_10625_),
    .Z(_07006_));
 MUX2_X1 _36604_ (.A(\itlb.vtag_cam.mem [7]),
    .B(_10534_),
    .S(_10625_),
    .Z(_07017_));
 MUX2_X1 _36605_ (.A(\itlb.vtag_cam.mem [8]),
    .B(_10535_),
    .S(_10625_),
    .Z(_07028_));
 BUF_X8 _36606_ (.A(_10624_),
    .Z(_10626_));
 MUX2_X1 _36607_ (.A(\itlb.vtag_cam.mem [9]),
    .B(_10536_),
    .S(_10626_),
    .Z(_07039_));
 MUX2_X1 _36608_ (.A(\itlb.vtag_cam.mem [10]),
    .B(_10538_),
    .S(_10626_),
    .Z(_06835_));
 MUX2_X1 _36609_ (.A(\itlb.vtag_cam.mem [11]),
    .B(_10539_),
    .S(_10626_),
    .Z(_06846_));
 MUX2_X1 _36610_ (.A(\itlb.vtag_cam.mem [12]),
    .B(_10540_),
    .S(_10626_),
    .Z(_06857_));
 MUX2_X1 _36611_ (.A(\itlb.vtag_cam.mem [13]),
    .B(_10541_),
    .S(_10626_),
    .Z(_06868_));
 MUX2_X1 _36612_ (.A(\itlb.vtag_cam.mem [14]),
    .B(_10542_),
    .S(_10626_),
    .Z(_06879_));
 MUX2_X1 _36613_ (.A(\itlb.vtag_cam.mem [15]),
    .B(_10543_),
    .S(_10626_),
    .Z(_06890_));
 MUX2_X1 _36614_ (.A(\itlb.vtag_cam.mem [16]),
    .B(_10544_),
    .S(_10626_),
    .Z(_06901_));
 MUX2_X1 _36615_ (.A(\itlb.vtag_cam.mem [17]),
    .B(_10545_),
    .S(_10626_),
    .Z(_06912_));
 MUX2_X1 _36616_ (.A(\itlb.vtag_cam.mem [18]),
    .B(_10546_),
    .S(_10626_),
    .Z(_06923_));
 MUX2_X1 _36617_ (.A(\itlb.vtag_cam.mem [19]),
    .B(_10547_),
    .S(_10624_),
    .Z(_06934_));
 MUX2_X1 _36618_ (.A(\itlb.vtag_cam.mem [20]),
    .B(_10548_),
    .S(_10624_),
    .Z(_06946_));
 MUX2_X1 _36619_ (.A(\itlb.vtag_cam.mem [21]),
    .B(_10549_),
    .S(_10624_),
    .Z(_06953_));
 MUX2_X1 _36620_ (.A(\itlb.vtag_cam.mem [22]),
    .B(_10550_),
    .S(_10624_),
    .Z(_06954_));
 MUX2_X1 _36621_ (.A(\itlb.vtag_cam.mem [23]),
    .B(_10551_),
    .S(_10624_),
    .Z(_06955_));
 MUX2_X1 _36622_ (.A(\itlb.vtag_cam.mem [24]),
    .B(_10552_),
    .S(_10624_),
    .Z(_06956_));
 MUX2_X1 _36623_ (.A(\itlb.vtag_cam.mem [25]),
    .B(_10553_),
    .S(_10624_),
    .Z(_06957_));
 MUX2_X1 _36624_ (.A(\itlb.vtag_cam.mem [26]),
    .B(_10554_),
    .S(_10624_),
    .Z(_06958_));
 INV_X1 _36625_ (.A(_10625_),
    .ZN(_10627_));
 NAND3_X1 _36626_ (.A1(_10627_),
    .A2(\itlb.vtag_cam.valid [7]),
    .A3(_10206_),
    .ZN(_10628_));
 NAND2_X1 _36627_ (.A1(_10628_),
    .A2(_10627_),
    .ZN(_07047_));
 OAI211_X1 _36628_ (.A(\itlb.vtag_cam.valid [6]),
    .B(_10206_),
    .C1(_10556_),
    .C2(_10559_),
    .ZN(_10629_));
 OAI21_X1 _36629_ (.A(_10629_),
    .B1(_10559_),
    .B2(_10556_),
    .ZN(_07046_));
 INV_X1 _36630_ (.A(_10620_),
    .ZN(_10630_));
 OAI21_X1 _36631_ (.A(_10630_),
    .B1(_10248_),
    .B2(_10071_),
    .ZN(_07045_));
 OAI21_X1 _36632_ (.A(_10613_),
    .B1(_10069_),
    .B2(_10071_),
    .ZN(_07044_));
 INV_X1 _36633_ (.A(_10609_),
    .ZN(_10631_));
 OAI21_X1 _36634_ (.A(_10631_),
    .B1(_10302_),
    .B2(_10071_),
    .ZN(_07043_));
 OAI22_X1 _36635_ (.A1(_10564_),
    .A2(_10559_),
    .B1(_10375_),
    .B2(_10071_),
    .ZN(_07042_));
 OAI22_X1 _36636_ (.A1(_10564_),
    .A2(_10565_),
    .B1(_10440_),
    .B2(_10071_),
    .ZN(_07040_));
 INV_X1 _36637_ (.A(_10527_),
    .ZN(_10632_));
 NAND3_X1 _36638_ (.A1(_10632_),
    .A2(\itlb.vtag_cam.valid [1]),
    .A3(_10206_),
    .ZN(_10633_));
 NAND2_X1 _36639_ (.A1(_10633_),
    .A2(_10632_),
    .ZN(_07041_));
 INV_X4 _36640_ (.A(_08521_),
    .ZN(_10634_));
 NOR3_X1 _36641_ (.A1(_10373_),
    .A2(_10476_),
    .A3(_10634_),
    .ZN(\itlb.miss_v_reg.N3 ));
 OR3_X4 _36642_ (.A1(cfg_addr_i[15]),
    .A2(cfg_addr_i[14]),
    .A3(cfg_addr_i[13]),
    .ZN(_10635_));
 OR4_X4 _36643_ (.A1(cfg_addr_i[12]),
    .A2(_10635_),
    .A3(cfg_addr_i[11]),
    .A4(cfg_addr_i[10]),
    .ZN(_10636_));
 OR3_X4 _36644_ (.A1(_10636_),
    .A2(cfg_addr_i[9]),
    .A3(cfg_addr_i[8]),
    .ZN(_10637_));
 NOR3_X4 _36645_ (.A1(_10637_),
    .A2(cfg_addr_i[7]),
    .A3(cfg_addr_i[6]),
    .ZN(_10638_));
 NAND2_X4 _36646_ (.A1(_10638_),
    .A2(cfg_addr_i[5]),
    .ZN(_10639_));
 NOR4_X2 _36647_ (.A1(_10639_),
    .A2(cfg_addr_i[4]),
    .A3(cfg_addr_i[3]),
    .A4(cfg_addr_i[2]),
    .ZN(_10640_));
 NAND2_X4 _36648_ (.A1(_10640_),
    .A2(cfg_addr_i[1]),
    .ZN(_10641_));
 NOR2_X1 _36649_ (.A1(_10641_),
    .A2(cfg_addr_i[0]),
    .ZN(_10642_));
 AND3_X2 _36650_ (.A1(_10642_),
    .A2(freeze_i),
    .A3(cfg_w_v_i),
    .ZN(_10643_));
 INV_X1 _36651_ (.A(_10643_),
    .ZN(_10644_));
 NAND3_X1 _36652_ (.A1(_10644_),
    .A2(\icache.N7 ),
    .A3(_08723_),
    .ZN(_10645_));
 NAND3_X1 _36653_ (.A1(_10643_),
    .A2(_08723_),
    .A3(cfg_data_i[0]),
    .ZN(_10646_));
 NAND2_X1 _36654_ (.A1(_10645_),
    .A2(_10646_),
    .ZN(_04888_));
 AND2_X1 _36655_ (.A1(_08023_),
    .A2(\icache.lce.lce_req_inst.state_r [0]),
    .ZN(_10647_));
 INV_X2 _36656_ (.A(_10647_),
    .ZN(_10648_));
 NAND2_X2 _36657_ (.A1(_08023_),
    .A2(_00002_),
    .ZN(_10649_));
 NAND2_X4 _36658_ (.A1(_10648_),
    .A2(_10649_),
    .ZN(lce_resp_o[40]));
 INV_X2 _36659_ (.A(_07979_),
    .ZN(_10650_));
 BUF_X16 _36660_ (.A(_10650_),
    .Z(_10651_));
 NOR2_X1 _36661_ (.A1(_07884_),
    .A2(_00584_),
    .ZN(_10652_));
 NOR2_X1 _36662_ (.A1(_07886_),
    .A2(_00583_),
    .ZN(_10653_));
 NOR2_X4 _36663_ (.A1(_10652_),
    .A2(_10653_),
    .ZN(_10654_));
 NOR3_X1 _36664_ (.A1(_10651_),
    .A2(_07892_),
    .A3(_10654_),
    .ZN(_10655_));
 INV_X8 _36665_ (.A(lce_resp_o[40]),
    .ZN(_10656_));
 BUF_X16 _36666_ (.A(_10656_),
    .Z(_10657_));
 MUX2_X2 _36667_ (.A(\icache.lce.lce_data_cmd.miss_addr_i [0]),
    .B(_10655_),
    .S(_10657_),
    .Z(lce_resp_o[0]));
 BUF_X8 _36668_ (.A(_07891_),
    .Z(_10658_));
 NOR2_X1 _36669_ (.A1(_07884_),
    .A2(_00586_),
    .ZN(_10659_));
 NOR2_X1 _36670_ (.A1(_07886_),
    .A2(_00585_),
    .ZN(_10660_));
 NOR2_X4 _36671_ (.A1(_10659_),
    .A2(_10660_),
    .ZN(_10661_));
 NOR3_X1 _36672_ (.A1(_10651_),
    .A2(_10658_),
    .A3(_10661_),
    .ZN(_10662_));
 MUX2_X2 _36673_ (.A(\icache.lce.lce_data_cmd.miss_addr_i [1]),
    .B(_10662_),
    .S(_10657_),
    .Z(lce_resp_o[1]));
 NOR2_X1 _36674_ (.A1(_07884_),
    .A2(_00588_),
    .ZN(_10663_));
 NOR2_X1 _36675_ (.A1(_07886_),
    .A2(_00587_),
    .ZN(_10664_));
 NOR2_X4 _36676_ (.A1(_10663_),
    .A2(_10664_),
    .ZN(_10665_));
 NOR3_X1 _36677_ (.A1(_10651_),
    .A2(_10658_),
    .A3(_10665_),
    .ZN(_10666_));
 MUX2_X2 _36678_ (.A(\icache.lce.lce_data_cmd.miss_addr_i [2]),
    .B(_10666_),
    .S(_10657_),
    .Z(lce_resp_o[2]));
 NOR2_X1 _36679_ (.A1(_07884_),
    .A2(_00590_),
    .ZN(_10667_));
 NOR2_X1 _36680_ (.A1(_07886_),
    .A2(_00589_),
    .ZN(_10668_));
 NOR2_X4 _36681_ (.A1(_10667_),
    .A2(_10668_),
    .ZN(_10669_));
 NOR3_X1 _36682_ (.A1(_10651_),
    .A2(_10658_),
    .A3(_10669_),
    .ZN(_10670_));
 MUX2_X2 _36683_ (.A(lce_req_o[10]),
    .B(_10670_),
    .S(_10657_),
    .Z(lce_resp_o[3]));
 BUF_X4 _36684_ (.A(_07979_),
    .Z(_10671_));
 NAND2_X1 _36685_ (.A1(_07884_),
    .A2(_00591_),
    .ZN(_10672_));
 NAND2_X2 _36686_ (.A1(_07973_),
    .A2(_00592_),
    .ZN(_10673_));
 AND4_X2 _36687_ (.A1(_07971_),
    .A2(_10671_),
    .A3(_10672_),
    .A4(_10673_),
    .ZN(_10674_));
 MUX2_X2 _36688_ (.A(lce_req_o[11]),
    .B(_10674_),
    .S(_10657_),
    .Z(lce_resp_o[4]));
 NAND2_X2 _36689_ (.A1(_07884_),
    .A2(_00593_),
    .ZN(_10675_));
 NAND2_X2 _36690_ (.A1(_07973_),
    .A2(_00594_),
    .ZN(_10676_));
 AND4_X4 _36691_ (.A1(_07971_),
    .A2(_10671_),
    .A3(_10675_),
    .A4(_10676_),
    .ZN(_10677_));
 MUX2_X2 _36692_ (.A(lce_req_o[12]),
    .B(_10677_),
    .S(_10657_),
    .Z(lce_resp_o[5]));
 BUF_X4 _36693_ (.A(_07978_),
    .Z(_10678_));
 BUF_X4 _36694_ (.A(_07889_),
    .Z(_10679_));
 AND4_X1 _36695_ (.A1(_07626_),
    .A2(_07976_),
    .A3(_10678_),
    .A4(_10679_),
    .ZN(_10680_));
 MUX2_X2 _36696_ (.A(_10680_),
    .B(lce_req_o[13]),
    .S(lce_resp_o[40]),
    .Z(lce_resp_o[6]));
 AND4_X1 _36697_ (.A1(_10678_),
    .A2(_07976_),
    .A3(_07632_),
    .A4(_10679_),
    .ZN(_10681_));
 MUX2_X2 _36698_ (.A(_10681_),
    .B(lce_req_o[14]),
    .S(lce_resp_o[40]),
    .Z(lce_resp_o[7]));
 AND4_X1 _36699_ (.A1(_10678_),
    .A2(_07976_),
    .A3(_07637_),
    .A4(_10679_),
    .ZN(_10682_));
 MUX2_X2 _36700_ (.A(_10682_),
    .B(lce_req_o[15]),
    .S(lce_resp_o[40]),
    .Z(lce_resp_o[8]));
 AND4_X4 _36701_ (.A1(_10678_),
    .A2(_07976_),
    .A3(_07642_),
    .A4(_10679_),
    .ZN(_10683_));
 MUX2_X2 _36702_ (.A(_10683_),
    .B(lce_req_o[16]),
    .S(lce_resp_o[40]),
    .Z(lce_resp_o[9]));
 AND4_X1 _36703_ (.A1(_10678_),
    .A2(_07976_),
    .A3(_07647_),
    .A4(_10679_),
    .ZN(_10684_));
 MUX2_X2 _36704_ (.A(_10684_),
    .B(lce_req_o[17]),
    .S(lce_resp_o[40]),
    .Z(lce_resp_o[10]));
 AND4_X2 _36705_ (.A1(_10678_),
    .A2(_07976_),
    .A3(_07652_),
    .A4(_07889_),
    .ZN(_10685_));
 MUX2_X2 _36706_ (.A(_10685_),
    .B(lce_req_o[18]),
    .S(lce_resp_o[40]),
    .Z(lce_resp_o[11]));
 NOR3_X4 _36707_ (.A1(_10651_),
    .A2(_07888_),
    .A3(_07891_),
    .ZN(_10686_));
 MUX2_X2 _36708_ (.A(lce_req_o[19]),
    .B(_10686_),
    .S(_10657_),
    .Z(lce_resp_o[12]));
 AND4_X1 _36709_ (.A1(_07971_),
    .A2(_10671_),
    .A3(_07901_),
    .A4(_07902_),
    .ZN(_10687_));
 MUX2_X2 _36710_ (.A(lce_req_o[20]),
    .B(_10687_),
    .S(_10657_),
    .Z(lce_resp_o[13]));
 NOR3_X4 _36711_ (.A1(_10651_),
    .A2(_10658_),
    .A3(_07905_),
    .ZN(_10688_));
 MUX2_X2 _36712_ (.A(lce_req_o[21]),
    .B(_10688_),
    .S(_10657_),
    .Z(lce_resp_o[14]));
 AND4_X1 _36713_ (.A1(_07971_),
    .A2(_10671_),
    .A3(_07907_),
    .A4(_07908_),
    .ZN(_10689_));
 BUF_X8 _36714_ (.A(_10656_),
    .Z(_10690_));
 MUX2_X2 _36715_ (.A(lce_req_o[22]),
    .B(_10689_),
    .S(_10690_),
    .Z(lce_resp_o[15]));
 AND4_X4 _36716_ (.A1(_07971_),
    .A2(_10671_),
    .A3(_07909_),
    .A4(_07910_),
    .ZN(_10691_));
 MUX2_X2 _36717_ (.A(lce_req_o[23]),
    .B(_10691_),
    .S(_10690_),
    .Z(lce_resp_o[16]));
 AND4_X2 _36718_ (.A1(_07971_),
    .A2(_10671_),
    .A3(_07911_),
    .A4(_07912_),
    .ZN(_10692_));
 MUX2_X2 _36719_ (.A(lce_req_o[24]),
    .B(_10692_),
    .S(_10690_),
    .Z(lce_resp_o[17]));
 NOR3_X4 _36720_ (.A1(_10651_),
    .A2(_10658_),
    .A3(_07916_),
    .ZN(_10693_));
 MUX2_X2 _36721_ (.A(lce_req_o[25]),
    .B(_10693_),
    .S(_10690_),
    .Z(lce_resp_o[18]));
 NOR3_X4 _36722_ (.A1(_10651_),
    .A2(_10658_),
    .A3(_07919_),
    .ZN(_10694_));
 MUX2_X2 _36723_ (.A(lce_req_o[26]),
    .B(_10694_),
    .S(_10690_),
    .Z(lce_resp_o[19]));
 AND4_X1 _36724_ (.A1(_07971_),
    .A2(_10671_),
    .A3(_07920_),
    .A4(_07921_),
    .ZN(_10695_));
 MUX2_X2 _36725_ (.A(lce_req_o[27]),
    .B(_10695_),
    .S(_10690_),
    .Z(lce_resp_o[20]));
 AND4_X1 _36726_ (.A1(_07971_),
    .A2(_10671_),
    .A3(_07922_),
    .A4(_07923_),
    .ZN(_10696_));
 MUX2_X2 _36727_ (.A(lce_req_o[28]),
    .B(_10696_),
    .S(_10690_),
    .Z(lce_resp_o[21]));
 NOR3_X1 _36728_ (.A1(_10651_),
    .A2(_10658_),
    .A3(_07926_),
    .ZN(_10697_));
 MUX2_X2 _36729_ (.A(lce_req_o[29]),
    .B(_10697_),
    .S(_10690_),
    .Z(lce_resp_o[22]));
 AND4_X1 _36730_ (.A1(_07971_),
    .A2(_10671_),
    .A3(_07927_),
    .A4(_07928_),
    .ZN(_10698_));
 MUX2_X2 _36731_ (.A(lce_req_o[30]),
    .B(_10698_),
    .S(_10690_),
    .Z(lce_resp_o[23]));
 AND4_X1 _36732_ (.A1(_10679_),
    .A2(_10671_),
    .A3(_07929_),
    .A4(_07930_),
    .ZN(_10699_));
 MUX2_X2 _36733_ (.A(lce_req_o[31]),
    .B(_10699_),
    .S(_10690_),
    .Z(lce_resp_o[24]));
 NOR3_X1 _36734_ (.A1(_10651_),
    .A2(_10658_),
    .A3(_07933_),
    .ZN(_10700_));
 BUF_X8 _36735_ (.A(_10656_),
    .Z(_10701_));
 MUX2_X2 _36736_ (.A(lce_req_o[32]),
    .B(_10700_),
    .S(_10701_),
    .Z(lce_resp_o[25]));
 BUF_X8 _36737_ (.A(_10650_),
    .Z(_10702_));
 NOR3_X1 _36738_ (.A1(_10702_),
    .A2(_10658_),
    .A3(_07936_),
    .ZN(_10703_));
 MUX2_X2 _36739_ (.A(lce_req_o[33]),
    .B(_10703_),
    .S(_10701_),
    .Z(lce_resp_o[26]));
 AND4_X1 _36740_ (.A1(_10679_),
    .A2(_07979_),
    .A3(_07937_),
    .A4(_07938_),
    .ZN(_10704_));
 MUX2_X2 _36741_ (.A(lce_req_o[34]),
    .B(_10704_),
    .S(_10701_),
    .Z(lce_resp_o[27]));
 AND4_X2 _36742_ (.A1(_10679_),
    .A2(_07979_),
    .A3(_07940_),
    .A4(_07941_),
    .ZN(_10705_));
 MUX2_X2 _36743_ (.A(lce_req_o[35]),
    .B(_10705_),
    .S(_10701_),
    .Z(lce_resp_o[28]));
 NOR3_X4 _36744_ (.A1(_10702_),
    .A2(_10658_),
    .A3(_07944_),
    .ZN(_10706_));
 MUX2_X2 _36745_ (.A(lce_req_o[36]),
    .B(_10706_),
    .S(_10701_),
    .Z(lce_resp_o[29]));
 AND4_X1 _36746_ (.A1(_10679_),
    .A2(_07979_),
    .A3(_07945_),
    .A4(_07946_),
    .ZN(_10707_));
 MUX2_X2 _36747_ (.A(lce_req_o[37]),
    .B(_10707_),
    .S(_10701_),
    .Z(lce_resp_o[30]));
 NOR3_X4 _36748_ (.A1(_10702_),
    .A2(_07891_),
    .A3(_07949_),
    .ZN(_10708_));
 MUX2_X2 _36749_ (.A(lce_req_o[38]),
    .B(_10708_),
    .S(_10701_),
    .Z(lce_resp_o[31]));
 NOR3_X4 _36750_ (.A1(_10702_),
    .A2(_07891_),
    .A3(_07952_),
    .ZN(_10709_));
 MUX2_X2 _36751_ (.A(lce_req_o[39]),
    .B(_10709_),
    .S(_10701_),
    .Z(lce_resp_o[32]));
 NOR3_X1 _36752_ (.A1(_10702_),
    .A2(_07891_),
    .A3(_07955_),
    .ZN(_10710_));
 MUX2_X2 _36753_ (.A(lce_req_o[40]),
    .B(_10710_),
    .S(_10701_),
    .Z(lce_resp_o[33]));
 NOR3_X1 _36754_ (.A1(_10702_),
    .A2(_07891_),
    .A3(_07958_),
    .ZN(_10711_));
 MUX2_X2 _36755_ (.A(lce_req_o[41]),
    .B(_10711_),
    .S(_10701_),
    .Z(lce_resp_o[34]));
 NOR3_X4 _36756_ (.A1(_10702_),
    .A2(_07891_),
    .A3(_07961_),
    .ZN(_10712_));
 MUX2_X2 _36757_ (.A(lce_req_o[42]),
    .B(_10712_),
    .S(_10656_),
    .Z(lce_resp_o[35]));
 AND4_X1 _36758_ (.A1(_10679_),
    .A2(_07979_),
    .A3(_07962_),
    .A4(_07963_),
    .ZN(_10713_));
 MUX2_X2 _36759_ (.A(lce_req_o[43]),
    .B(_10713_),
    .S(_10656_),
    .Z(lce_resp_o[36]));
 NOR3_X1 _36760_ (.A1(_10702_),
    .A2(_07891_),
    .A3(_07966_),
    .ZN(_10714_));
 MUX2_X2 _36761_ (.A(lce_req_o[44]),
    .B(_10714_),
    .S(_10656_),
    .Z(lce_resp_o[37]));
 NOR3_X4 _36762_ (.A1(_10702_),
    .A2(_07891_),
    .A3(_07969_),
    .ZN(_10715_));
 MUX2_X2 _36763_ (.A(lce_req_o[45]),
    .B(_10715_),
    .S(_10656_),
    .Z(lce_resp_o[38]));
 NAND3_X4 _36764_ (.A1(_08023_),
    .A2(\icache.lce.lce_req_inst.state_r [0]),
    .A3(_08018_),
    .ZN(_10716_));
 INV_X4 _36765_ (.A(_07981_),
    .ZN(_10717_));
 OAI21_X4 _36766_ (.A(_10716_),
    .B1(_10717_),
    .B2(lce_resp_o[40]),
    .ZN(lce_resp_o[39]));
 NOR2_X1 _36767_ (.A1(_07884_),
    .A2(_00596_),
    .ZN(_10718_));
 NOR2_X1 _36768_ (.A1(_07973_),
    .A2(_00595_),
    .ZN(_10719_));
 NOR2_X4 _36769_ (.A1(_10718_),
    .A2(_10719_),
    .ZN(_10720_));
 NAND3_X2 _36770_ (.A1(_07618_),
    .A2(_08009_),
    .A3(_10678_),
    .ZN(_10721_));
 AOI211_X2 _36771_ (.A(lce_resp_o[40]),
    .B(_10720_),
    .C1(_10717_),
    .C2(_10721_),
    .ZN(lce_resp_o[42]));
 INV_X2 _36772_ (.A(_07656_),
    .ZN(_10722_));
 INV_X1 _36773_ (.A(\icache.lce.lce_cmd_inst.N0 ),
    .ZN(_10723_));
 AOI21_X1 _36774_ (.A(_07898_),
    .B1(_07979_),
    .B2(_10723_),
    .ZN(_10724_));
 INV_X1 _36775_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.empty_r ),
    .ZN(_10725_));
 AND3_X1 _36776_ (.A1(_07604_),
    .A2(_10725_),
    .A3(_07605_),
    .ZN(_10726_));
 INV_X1 _36777_ (.A(_10726_),
    .ZN(_10727_));
 OAI21_X2 _36778_ (.A(_10722_),
    .B1(_10724_),
    .B2(_10727_),
    .ZN(_10728_));
 INV_X2 _36779_ (.A(_10728_),
    .ZN(_10729_));
 NOR2_X4 _36780_ (.A1(_08037_),
    .A2(_10729_),
    .ZN(\icache.lce.lce_cmd_inst.tag_mem_pkt_yumi_i ));
 NAND4_X4 _36781_ (.A1(_07618_),
    .A2(_00001_),
    .A3(_08009_),
    .A4(_07978_),
    .ZN(_10730_));
 AOI21_X2 _36782_ (.A(\icache.lce.lce_cmd_inst.N0 ),
    .B1(_08480_),
    .B2(_10728_),
    .ZN(_10731_));
 OAI21_X1 _36783_ (.A(_10730_),
    .B1(_10731_),
    .B2(_10717_),
    .ZN(_10732_));
 AND3_X1 _36784_ (.A1(_10648_),
    .A2(lce_resp_ready_i),
    .A3(_10649_),
    .ZN(_10733_));
 AND2_X1 _36785_ (.A1(_10732_),
    .A2(_10733_),
    .ZN(_10734_));
 NOR3_X1 _36786_ (.A1(_10734_),
    .A2(_10702_),
    .A3(_10731_),
    .ZN(_10735_));
 AOI21_X1 _36787_ (.A(_00597_),
    .B1(_07976_),
    .B2(_10678_),
    .ZN(_10736_));
 NAND2_X1 _36788_ (.A1(_07605_),
    .A2(_00598_),
    .ZN(_10737_));
 NOR3_X1 _36789_ (.A1(_10735_),
    .A2(_10736_),
    .A3(_10737_),
    .ZN(_10738_));
 AOI211_X1 _36790_ (.A(_08957_),
    .B(_10738_),
    .C1(_10723_),
    .C2(_10737_),
    .ZN(_05402_));
 BUF_X8 _36791_ (.A(_08722_),
    .Z(_10739_));
 AND2_X2 _36792_ (.A1(_08747_),
    .A2(_08748_),
    .ZN(_10740_));
 BUF_X4 _36793_ (.A(fe_cmd_i[33]),
    .Z(_10741_));
 AND3_X1 _36794_ (.A1(_08324_),
    .A2(fe_cmd_v_i),
    .A3(_10741_),
    .ZN(_10742_));
 NOR2_X1 _36795_ (.A1(_08323_),
    .A2(fe_cmd_i[74]),
    .ZN(_10743_));
 AND2_X4 _36796_ (.A1(_10742_),
    .A2(_10743_),
    .ZN(_10744_));
 OR3_X4 _36797_ (.A1(_10740_),
    .A2(_08743_),
    .A3(_10744_),
    .ZN(_10745_));
 INV_X8 _36798_ (.A(_10744_),
    .ZN(_10746_));
 OR2_X2 _36799_ (.A1(_10746_),
    .A2(fe_cmd_i[15]),
    .ZN(_10747_));
 AND2_X1 _36800_ (.A1(_10745_),
    .A2(_10747_),
    .ZN(_10748_));
 NAND3_X4 _36801_ (.A1(_08475_),
    .A2(_08478_),
    .A3(_10746_),
    .ZN(_10749_));
 OR2_X2 _36802_ (.A1(_10746_),
    .A2(fe_cmd_i[16]),
    .ZN(_10750_));
 AND3_X4 _36803_ (.A1(_10748_),
    .A2(_10749_),
    .A3(_10750_),
    .ZN(_10751_));
 NAND2_X1 _36804_ (.A1(_08755_),
    .A2(_10746_),
    .ZN(_10752_));
 AND2_X1 _36805_ (.A1(_08510_),
    .A2(fe_cmd_i[20]),
    .ZN(_10753_));
 OR3_X4 _36806_ (.A1(_10746_),
    .A2(_10753_),
    .A3(fe_cmd_i[17]),
    .ZN(_10754_));
 NAND2_X4 _36807_ (.A1(_10752_),
    .A2(_10754_),
    .ZN(_10755_));
 AND2_X4 _36808_ (.A1(_10751_),
    .A2(_10755_),
    .ZN(_10756_));
 BUF_X32 _36809_ (.A(net112),
    .Z(_10757_));
 NAND2_X2 _36810_ (.A1(_08757_),
    .A2(_10746_),
    .ZN(_10758_));
 AND2_X1 _36811_ (.A1(_08510_),
    .A2(fe_cmd_i[21]),
    .ZN(_10759_));
 OR3_X4 _36812_ (.A1(_10746_),
    .A2(_10759_),
    .A3(fe_cmd_i[18]),
    .ZN(_10760_));
 NAND2_X4 _36813_ (.A1(_10758_),
    .A2(_10760_),
    .ZN(_10761_));
 BUF_X32 _36814_ (.A(_10744_),
    .Z(_10762_));
 OR3_X4 _36815_ (.A1(_08351_),
    .A2(_08358_),
    .A3(_10762_),
    .ZN(_10763_));
 AND2_X1 _36816_ (.A1(_08510_),
    .A2(fe_cmd_i[22]),
    .ZN(_10764_));
 OR3_X4 _36817_ (.A1(_10746_),
    .A2(_10764_),
    .A3(fe_cmd_i[19]),
    .ZN(_10765_));
 NAND2_X4 _36818_ (.A1(_10763_),
    .A2(_10765_),
    .ZN(_10766_));
 OR2_X4 _36819_ (.A1(_10761_),
    .A2(_10766_),
    .ZN(_10767_));
 OR3_X2 _36820_ (.A1(_08365_),
    .A2(_08368_),
    .A3(_10762_),
    .ZN(_10768_));
 AOI21_X4 _36821_ (.A(fe_cmd_i[20]),
    .B1(_08510_),
    .B2(fe_cmd_i[23]),
    .ZN(_10769_));
 NAND2_X1 _36822_ (.A1(_10769_),
    .A2(_10762_),
    .ZN(_10770_));
 NAND2_X4 _36823_ (.A1(_10768_),
    .A2(_10770_),
    .ZN(_10771_));
 NOR2_X4 _36824_ (.A1(_10767_),
    .A2(_10771_),
    .ZN(_10772_));
 AND2_X4 _36825_ (.A1(_10757_),
    .A2(net107),
    .ZN(_10773_));
 INV_X8 _36826_ (.A(_10773_),
    .ZN(_10774_));
 BUF_X8 _36827_ (.A(_10746_),
    .Z(_10775_));
 BUF_X4 _36828_ (.A(_10775_),
    .Z(_10776_));
 OAI211_X1 _36829_ (.A(\bp_fe_pc_gen_1.btb.v_r [59]),
    .B(_10739_),
    .C1(_10774_),
    .C2(_10776_),
    .ZN(_10777_));
 BUF_X32 _36830_ (.A(net113),
    .Z(_10778_));
 BUF_X32 _36831_ (.A(_10778_),
    .Z(_10779_));
 BUF_X32 _36832_ (.A(_10779_),
    .Z(_10780_));
 BUF_X32 _36833_ (.A(_10780_),
    .Z(_10781_));
 BUF_X8 _36834_ (.A(_10781_),
    .Z(_10782_));
 BUF_X8 _36835_ (.A(_08722_),
    .Z(_10783_));
 BUF_X32 _36836_ (.A(_10762_),
    .Z(_10784_));
 BUF_X16 _36837_ (.A(_10784_),
    .Z(_10785_));
 BUF_X8 _36838_ (.A(_10785_),
    .Z(_10786_));
 BUF_X16 _36839_ (.A(net105),
    .Z(_10787_));
 BUF_X16 _36840_ (.A(_10787_),
    .Z(_10788_));
 BUF_X16 _36841_ (.A(_10788_),
    .Z(_10789_));
 BUF_X16 _36842_ (.A(_10789_),
    .Z(_10790_));
 BUF_X8 _36843_ (.A(_10790_),
    .Z(_10791_));
 BUF_X8 _36844_ (.A(_10791_),
    .Z(_10792_));
 NAND4_X1 _36845_ (.A1(_10782_),
    .A2(_10783_),
    .A3(_10786_),
    .A4(_10792_),
    .ZN(_10793_));
 NAND2_X1 _36846_ (.A1(_10777_),
    .A2(_10793_),
    .ZN(_00812_));
 INV_X1 _36847_ (.A(_10755_),
    .ZN(_10794_));
 BUF_X8 _36848_ (.A(_10794_),
    .Z(_10795_));
 AND2_X4 _36849_ (.A1(_10751_),
    .A2(_10795_),
    .ZN(_10796_));
 BUF_X32 _36850_ (.A(net88),
    .Z(_10797_));
 BUF_X32 _36851_ (.A(_10797_),
    .Z(_10798_));
 AND2_X4 _36852_ (.A1(_10798_),
    .A2(_10787_),
    .ZN(_10799_));
 BUF_X16 _36853_ (.A(_10799_),
    .Z(_10800_));
 INV_X8 _36854_ (.A(_10800_),
    .ZN(_10801_));
 OAI211_X1 _36855_ (.A(\bp_fe_pc_gen_1.btb.v_r [63]),
    .B(_10739_),
    .C1(_10801_),
    .C2(_10776_),
    .ZN(_10802_));
 BUF_X32 _36856_ (.A(_10798_),
    .Z(_10803_));
 BUF_X32 _36857_ (.A(_10803_),
    .Z(_10804_));
 BUF_X32 _36858_ (.A(_10804_),
    .Z(_10805_));
 BUF_X8 _36859_ (.A(_10805_),
    .Z(_10806_));
 NAND4_X2 _36860_ (.A1(_10806_),
    .A2(_10783_),
    .A3(_10786_),
    .A4(_10792_),
    .ZN(_10807_));
 NAND2_X1 _36861_ (.A1(_10802_),
    .A2(_10807_),
    .ZN(_00817_));
 NAND2_X4 _36862_ (.A1(_10749_),
    .A2(_10750_),
    .ZN(_10808_));
 AOI21_X4 _36863_ (.A(_10808_),
    .B1(_10745_),
    .B2(_10747_),
    .ZN(_10809_));
 AND2_X4 _36864_ (.A1(_10809_),
    .A2(_10794_),
    .ZN(_10810_));
 BUF_X32 _36865_ (.A(net86),
    .Z(_10811_));
 AND2_X4 _36866_ (.A1(_10811_),
    .A2(_10787_),
    .ZN(_10812_));
 BUF_X16 _36867_ (.A(_10812_),
    .Z(_10813_));
 INV_X1 _36868_ (.A(_10813_),
    .ZN(_10814_));
 OAI211_X1 _36869_ (.A(\bp_fe_pc_gen_1.btb.v_r [62]),
    .B(_10739_),
    .C1(_10814_),
    .C2(_10776_),
    .ZN(_10815_));
 BUF_X32 _36870_ (.A(net84),
    .Z(_10816_));
 BUF_X32 _36871_ (.A(_10816_),
    .Z(_10817_));
 BUF_X32 _36872_ (.A(_10817_),
    .Z(_10818_));
 BUF_X32 _36873_ (.A(_10818_),
    .Z(_10819_));
 BUF_X8 _36874_ (.A(_10819_),
    .Z(_10820_));
 NAND4_X1 _36875_ (.A1(_10820_),
    .A2(_10783_),
    .A3(_10786_),
    .A4(_10792_),
    .ZN(_10821_));
 NAND2_X1 _36876_ (.A1(_10815_),
    .A2(_10821_),
    .ZN(_00816_));
 NAND3_X4 _36877_ (.A1(_10808_),
    .A2(_10745_),
    .A3(_10747_),
    .ZN(_10822_));
 NOR2_X4 _36878_ (.A1(_10822_),
    .A2(_10755_),
    .ZN(_10823_));
 BUF_X32 _36879_ (.A(net79),
    .Z(_10824_));
 BUF_X16 _36880_ (.A(net104),
    .Z(_10825_));
 AND2_X4 _36881_ (.A1(_10824_),
    .A2(_10825_),
    .ZN(_10826_));
 INV_X1 _36882_ (.A(_10826_),
    .ZN(_10827_));
 OAI211_X1 _36883_ (.A(\bp_fe_pc_gen_1.btb.v_r [61]),
    .B(_10739_),
    .C1(_10827_),
    .C2(_10776_),
    .ZN(_10828_));
 BUF_X32 _36884_ (.A(_10824_),
    .Z(_10829_));
 BUF_X32 _36885_ (.A(_10829_),
    .Z(_10830_));
 BUF_X32 _36886_ (.A(_10830_),
    .Z(_10831_));
 BUF_X16 _36887_ (.A(_10831_),
    .Z(_10832_));
 BUF_X8 _36888_ (.A(_10832_),
    .Z(_10833_));
 NAND4_X1 _36889_ (.A1(_10833_),
    .A2(_10783_),
    .A3(_10786_),
    .A4(_10792_),
    .ZN(_10834_));
 NAND2_X1 _36890_ (.A1(_10828_),
    .A2(_10834_),
    .ZN(_00815_));
 INV_X1 _36891_ (.A(_10748_),
    .ZN(_10835_));
 NAND2_X2 _36892_ (.A1(_10835_),
    .A2(_10808_),
    .ZN(_10836_));
 NOR2_X4 _36893_ (.A1(_10836_),
    .A2(_10755_),
    .ZN(_10837_));
 AND2_X4 _36894_ (.A1(net69),
    .A2(net109),
    .ZN(_10838_));
 BUF_X16 _36895_ (.A(_10838_),
    .Z(_10839_));
 INV_X8 _36896_ (.A(_10839_),
    .ZN(_10840_));
 OAI211_X1 _36897_ (.A(\bp_fe_pc_gen_1.btb.v_r [60]),
    .B(_10739_),
    .C1(_10840_),
    .C2(_10776_),
    .ZN(_10841_));
 BUF_X32 _36898_ (.A(net72),
    .Z(_10842_));
 BUF_X32 _36899_ (.A(_10842_),
    .Z(_10843_));
 BUF_X16 _36900_ (.A(_10843_),
    .Z(_10844_));
 BUF_X32 _36901_ (.A(_10844_),
    .Z(_10845_));
 BUF_X8 _36902_ (.A(_10845_),
    .Z(_10846_));
 BUF_X4 _36903_ (.A(_08722_),
    .Z(_10847_));
 NAND4_X1 _36904_ (.A1(_10846_),
    .A2(_10847_),
    .A3(_10786_),
    .A4(_10792_),
    .ZN(_10848_));
 NAND2_X1 _36905_ (.A1(_10841_),
    .A2(_10848_),
    .ZN(_00814_));
 AND2_X4 _36906_ (.A1(_10809_),
    .A2(_10755_),
    .ZN(_10849_));
 AND2_X1 _36907_ (.A1(_10849_),
    .A2(net104),
    .ZN(_10850_));
 BUF_X8 _36908_ (.A(_10850_),
    .Z(_10851_));
 INV_X16 _36909_ (.A(_10851_),
    .ZN(_10852_));
 OAI211_X1 _36910_ (.A(\bp_fe_pc_gen_1.btb.v_r [58]),
    .B(_10739_),
    .C1(_10852_),
    .C2(_10776_),
    .ZN(_10853_));
 BUF_X32 _36911_ (.A(_10849_),
    .Z(_10854_));
 BUF_X32 _36912_ (.A(_10854_),
    .Z(_10855_));
 BUF_X32 _36913_ (.A(_10855_),
    .Z(_10856_));
 BUF_X32 _36914_ (.A(_10856_),
    .Z(_10857_));
 BUF_X16 _36915_ (.A(_10857_),
    .Z(_10858_));
 BUF_X16 _36916_ (.A(_10858_),
    .Z(_10859_));
 BUF_X8 _36917_ (.A(_10859_),
    .Z(_10860_));
 NAND4_X2 _36918_ (.A1(_10860_),
    .A2(_10847_),
    .A3(_10786_),
    .A4(_10792_),
    .ZN(_10861_));
 NAND2_X1 _36919_ (.A1(_10853_),
    .A2(_10861_),
    .ZN(_00811_));
 NOR2_X4 _36920_ (.A1(_10822_),
    .A2(_10795_),
    .ZN(_10862_));
 AND2_X4 _36921_ (.A1(net66),
    .A2(net108),
    .ZN(_10863_));
 INV_X8 _36922_ (.A(_10863_),
    .ZN(_10864_));
 OAI211_X1 _36923_ (.A(\bp_fe_pc_gen_1.btb.v_r [57]),
    .B(_10739_),
    .C1(_10864_),
    .C2(_10776_),
    .ZN(_10865_));
 BUF_X32 _36924_ (.A(net63),
    .Z(_10866_));
 BUF_X32 _36925_ (.A(_10866_),
    .Z(_10867_));
 BUF_X32 _36926_ (.A(_10867_),
    .Z(_10868_));
 BUF_X32 _36927_ (.A(_10868_),
    .Z(_10869_));
 BUF_X8 _36928_ (.A(_10869_),
    .Z(_10870_));
 NAND4_X1 _36929_ (.A1(_10870_),
    .A2(_10847_),
    .A3(_10786_),
    .A4(_10792_),
    .ZN(_10871_));
 NAND2_X1 _36930_ (.A1(_10865_),
    .A2(_10871_),
    .ZN(_00810_));
 NOR2_X4 _36931_ (.A1(_10836_),
    .A2(_10795_),
    .ZN(_10872_));
 BUF_X32 _36932_ (.A(net60),
    .Z(_10873_));
 AND2_X4 _36933_ (.A1(_10873_),
    .A2(net109),
    .ZN(_10874_));
 INV_X8 _36934_ (.A(_10874_),
    .ZN(_10875_));
 OAI211_X1 _36935_ (.A(\bp_fe_pc_gen_1.btb.v_r [56]),
    .B(_10739_),
    .C1(_10875_),
    .C2(_10776_),
    .ZN(_10876_));
 BUF_X32 _36936_ (.A(net60),
    .Z(_10877_));
 BUF_X32 _36937_ (.A(_10877_),
    .Z(_10878_));
 BUF_X32 _36938_ (.A(_10878_),
    .Z(_10879_));
 BUF_X32 _36939_ (.A(_10879_),
    .Z(_10880_));
 BUF_X8 _36940_ (.A(_10880_),
    .Z(_10881_));
 NAND4_X1 _36941_ (.A1(_10881_),
    .A2(_10847_),
    .A3(_10786_),
    .A4(_10792_),
    .ZN(_10882_));
 NAND2_X1 _36942_ (.A1(_10876_),
    .A2(_10882_),
    .ZN(_00809_));
 BUF_X4 _36943_ (.A(_08674_),
    .Z(_10883_));
 NAND3_X4 _36944_ (.A1(_10761_),
    .A2(_10765_),
    .A3(_10763_),
    .ZN(_10884_));
 NOR2_X4 _36945_ (.A1(_10884_),
    .A2(_10771_),
    .ZN(_10885_));
 BUF_X8 _36946_ (.A(_10885_),
    .Z(_10886_));
 AND2_X4 _36947_ (.A1(net92),
    .A2(_10886_),
    .ZN(_10887_));
 INV_X8 _36948_ (.A(_10887_),
    .ZN(_10888_));
 OAI211_X1 _36949_ (.A(\bp_fe_pc_gen_1.btb.v_r [55]),
    .B(_10883_),
    .C1(_10888_),
    .C2(_10776_),
    .ZN(_10889_));
 BUF_X8 _36950_ (.A(_10885_),
    .Z(_10890_));
 BUF_X8 _36951_ (.A(_10890_),
    .Z(_10891_));
 BUF_X8 _36952_ (.A(_10891_),
    .Z(_10892_));
 BUF_X16 _36953_ (.A(_10892_),
    .Z(_10893_));
 BUF_X8 _36954_ (.A(_10893_),
    .Z(_10894_));
 NAND4_X1 _36955_ (.A1(_10806_),
    .A2(_10847_),
    .A3(_10786_),
    .A4(_10894_),
    .ZN(_10895_));
 NAND2_X1 _36956_ (.A1(_10889_),
    .A2(_10895_),
    .ZN(_00808_));
 AND2_X4 _36957_ (.A1(net83),
    .A2(_10885_),
    .ZN(_10896_));
 INV_X16 _36958_ (.A(_10896_),
    .ZN(_10897_));
 OAI211_X1 _36959_ (.A(\bp_fe_pc_gen_1.btb.v_r [54]),
    .B(_10883_),
    .C1(_10897_),
    .C2(_10776_),
    .ZN(_10898_));
 BUF_X4 _36960_ (.A(_10785_),
    .Z(_10899_));
 NAND4_X1 _36961_ (.A1(_10820_),
    .A2(_10847_),
    .A3(_10899_),
    .A4(_10894_),
    .ZN(_10900_));
 NAND2_X1 _36962_ (.A1(_10898_),
    .A2(_10900_),
    .ZN(_00807_));
 BUF_X32 _36963_ (.A(net78),
    .Z(_10901_));
 AND2_X4 _36964_ (.A1(_10901_),
    .A2(_10886_),
    .ZN(_10902_));
 INV_X8 _36965_ (.A(_10902_),
    .ZN(_10903_));
 BUF_X4 _36966_ (.A(_10775_),
    .Z(_10904_));
 OAI211_X1 _36967_ (.A(\bp_fe_pc_gen_1.btb.v_r [53]),
    .B(_10883_),
    .C1(_10903_),
    .C2(_10904_),
    .ZN(_10905_));
 NAND4_X1 _36968_ (.A1(_10833_),
    .A2(_10847_),
    .A3(_10899_),
    .A4(_10894_),
    .ZN(_10906_));
 NAND2_X1 _36969_ (.A1(_10905_),
    .A2(_10906_),
    .ZN(_00806_));
 AND2_X4 _36970_ (.A1(net70),
    .A2(_10885_),
    .ZN(_10907_));
 INV_X16 _36971_ (.A(_10907_),
    .ZN(_10908_));
 OAI211_X1 _36972_ (.A(\bp_fe_pc_gen_1.btb.v_r [52]),
    .B(_10883_),
    .C1(_10908_),
    .C2(_10904_),
    .ZN(_10909_));
 NAND4_X1 _36973_ (.A1(_10846_),
    .A2(_10847_),
    .A3(_10899_),
    .A4(_10894_),
    .ZN(_10910_));
 NAND2_X1 _36974_ (.A1(_10909_),
    .A2(_10910_),
    .ZN(_00805_));
 AND2_X4 _36975_ (.A1(net110),
    .A2(_10885_),
    .ZN(_10911_));
 BUF_X16 _36976_ (.A(_10911_),
    .Z(_10912_));
 INV_X8 _36977_ (.A(_10912_),
    .ZN(_10913_));
 OAI211_X1 _36978_ (.A(\bp_fe_pc_gen_1.btb.v_r [51]),
    .B(_10883_),
    .C1(_10913_),
    .C2(_10904_),
    .ZN(_10914_));
 NAND4_X1 _36979_ (.A1(_10782_),
    .A2(_10847_),
    .A3(_10899_),
    .A4(_10894_),
    .ZN(_10915_));
 NAND2_X1 _36980_ (.A1(_10914_),
    .A2(_10915_),
    .ZN(_00804_));
 AND2_X4 _36981_ (.A1(_10854_),
    .A2(_10885_),
    .ZN(_10916_));
 INV_X8 _36982_ (.A(_10916_),
    .ZN(_10917_));
 OAI211_X1 _36983_ (.A(\bp_fe_pc_gen_1.btb.v_r [50]),
    .B(_10883_),
    .C1(_10917_),
    .C2(_10904_),
    .ZN(_10918_));
 NAND4_X1 _36984_ (.A1(_10860_),
    .A2(_10847_),
    .A3(_10899_),
    .A4(_10894_),
    .ZN(_10919_));
 NAND2_X1 _36985_ (.A1(_10918_),
    .A2(_10919_),
    .ZN(_00803_));
 BUF_X32 _36986_ (.A(net65),
    .Z(_10920_));
 AND2_X4 _36987_ (.A1(_10920_),
    .A2(_10890_),
    .ZN(_10921_));
 BUF_X16 _36988_ (.A(_10921_),
    .Z(_10922_));
 INV_X8 _36989_ (.A(_10922_),
    .ZN(_10923_));
 OAI211_X1 _36990_ (.A(\bp_fe_pc_gen_1.btb.v_r [49]),
    .B(_10883_),
    .C1(_10923_),
    .C2(_10904_),
    .ZN(_10924_));
 BUF_X4 _36991_ (.A(_08722_),
    .Z(_10925_));
 NAND4_X2 _36992_ (.A1(_10870_),
    .A2(_10925_),
    .A3(_10899_),
    .A4(_10894_),
    .ZN(_10926_));
 NAND2_X1 _36993_ (.A1(_10924_),
    .A2(_10926_),
    .ZN(_00801_));
 AND2_X2 _36994_ (.A1(net61),
    .A2(_10885_),
    .ZN(_10927_));
 BUF_X16 _36995_ (.A(_10927_),
    .Z(_10928_));
 BUF_X16 _36996_ (.A(_10928_),
    .Z(_10929_));
 INV_X8 _36997_ (.A(_10929_),
    .ZN(_10930_));
 OAI211_X1 _36998_ (.A(\bp_fe_pc_gen_1.btb.v_r [48]),
    .B(_10883_),
    .C1(_10930_),
    .C2(_10904_),
    .ZN(_10931_));
 NAND4_X1 _36999_ (.A1(_10881_),
    .A2(_10925_),
    .A3(_10899_),
    .A4(_10894_),
    .ZN(_10932_));
 NAND2_X1 _37000_ (.A1(_10931_),
    .A2(_10932_),
    .ZN(_00800_));
 NAND3_X4 _37001_ (.A1(_10766_),
    .A2(_10760_),
    .A3(_10758_),
    .ZN(_10933_));
 NOR2_X4 _37002_ (.A1(_10933_),
    .A2(_10771_),
    .ZN(_10934_));
 BUF_X16 _37003_ (.A(_10934_),
    .Z(_10935_));
 AND2_X4 _37004_ (.A1(_10797_),
    .A2(_10935_),
    .ZN(_10936_));
 INV_X16 _37005_ (.A(_10936_),
    .ZN(_10937_));
 OAI211_X1 _37006_ (.A(\bp_fe_pc_gen_1.btb.v_r [47]),
    .B(_10883_),
    .C1(_10937_),
    .C2(_10904_),
    .ZN(_10938_));
 BUF_X8 _37007_ (.A(_10935_),
    .Z(_10939_));
 BUF_X8 _37008_ (.A(_10939_),
    .Z(_10940_));
 BUF_X8 _37009_ (.A(_10940_),
    .Z(_10941_));
 BUF_X8 _37010_ (.A(_10941_),
    .Z(_10942_));
 BUF_X8 _37011_ (.A(_10942_),
    .Z(_10943_));
 NAND4_X2 _37012_ (.A1(_10806_),
    .A2(_10925_),
    .A3(_10899_),
    .A4(_10943_),
    .ZN(_10944_));
 NAND2_X1 _37013_ (.A1(_10938_),
    .A2(_10944_),
    .ZN(_00799_));
 AND2_X4 _37014_ (.A1(net83),
    .A2(_10934_),
    .ZN(_10945_));
 INV_X16 _37015_ (.A(_10945_),
    .ZN(_10946_));
 OAI211_X1 _37016_ (.A(\bp_fe_pc_gen_1.btb.v_r [46]),
    .B(_10883_),
    .C1(_10946_),
    .C2(_10904_),
    .ZN(_10947_));
 NAND4_X1 _37017_ (.A1(_10820_),
    .A2(_10925_),
    .A3(_10899_),
    .A4(_10943_),
    .ZN(_10948_));
 NAND2_X1 _37018_ (.A1(_10947_),
    .A2(_10948_),
    .ZN(_00798_));
 BUF_X4 _37019_ (.A(_08674_),
    .Z(_10949_));
 AND2_X4 _37020_ (.A1(net82),
    .A2(_10934_),
    .ZN(_10950_));
 INV_X8 _37021_ (.A(_10950_),
    .ZN(_10951_));
 OAI211_X1 _37022_ (.A(\bp_fe_pc_gen_1.btb.v_r [45]),
    .B(_10949_),
    .C1(_10951_),
    .C2(_10904_),
    .ZN(_10952_));
 NAND4_X1 _37023_ (.A1(_10833_),
    .A2(_10925_),
    .A3(_10899_),
    .A4(_10943_),
    .ZN(_10953_));
 NAND2_X1 _37024_ (.A1(_10952_),
    .A2(_10953_),
    .ZN(_00797_));
 AND2_X2 _37025_ (.A1(net69),
    .A2(_10935_),
    .ZN(_10954_));
 BUF_X16 _37026_ (.A(_10954_),
    .Z(_10955_));
 BUF_X16 _37027_ (.A(_10955_),
    .Z(_10956_));
 INV_X16 _37028_ (.A(_10956_),
    .ZN(_10957_));
 OAI211_X1 _37029_ (.A(\bp_fe_pc_gen_1.btb.v_r [44]),
    .B(_10949_),
    .C1(_10957_),
    .C2(_10904_),
    .ZN(_10958_));
 BUF_X2 _37030_ (.A(_10785_),
    .Z(_10959_));
 NAND4_X1 _37031_ (.A1(_10846_),
    .A2(_10925_),
    .A3(_10959_),
    .A4(_10943_),
    .ZN(_10960_));
 NAND2_X1 _37032_ (.A1(_10958_),
    .A2(_10960_),
    .ZN(_00796_));
 AND2_X4 _37033_ (.A1(_10757_),
    .A2(_10935_),
    .ZN(_10961_));
 BUF_X16 _37034_ (.A(_10961_),
    .Z(_10962_));
 INV_X16 _37035_ (.A(_10962_),
    .ZN(_10963_));
 BUF_X4 _37036_ (.A(_10775_),
    .Z(_10964_));
 OAI211_X1 _37037_ (.A(\bp_fe_pc_gen_1.btb.v_r [43]),
    .B(_10949_),
    .C1(_10963_),
    .C2(_10964_),
    .ZN(_10965_));
 NAND4_X1 _37038_ (.A1(_10782_),
    .A2(_10925_),
    .A3(_10959_),
    .A4(_10943_),
    .ZN(_10966_));
 NAND2_X1 _37039_ (.A1(_10965_),
    .A2(_10966_),
    .ZN(_00795_));
 AND2_X2 _37040_ (.A1(_10854_),
    .A2(_10934_),
    .ZN(_10967_));
 BUF_X16 _37041_ (.A(_10967_),
    .Z(_10968_));
 INV_X16 _37042_ (.A(_10968_),
    .ZN(_10969_));
 OAI211_X1 _37043_ (.A(\bp_fe_pc_gen_1.btb.v_r [42]),
    .B(_10949_),
    .C1(_10969_),
    .C2(_10964_),
    .ZN(_10970_));
 NAND4_X1 _37044_ (.A1(_10860_),
    .A2(_10925_),
    .A3(_10959_),
    .A4(_10943_),
    .ZN(_10971_));
 NAND2_X1 _37045_ (.A1(_10970_),
    .A2(_10971_),
    .ZN(_00794_));
 AND2_X4 _37046_ (.A1(net67),
    .A2(_10934_),
    .ZN(_10972_));
 INV_X16 _37047_ (.A(_10972_),
    .ZN(_10973_));
 OAI211_X1 _37048_ (.A(\bp_fe_pc_gen_1.btb.v_r [41]),
    .B(_10949_),
    .C1(_10973_),
    .C2(_10964_),
    .ZN(_10974_));
 NAND4_X1 _37049_ (.A1(_10870_),
    .A2(_10925_),
    .A3(_10959_),
    .A4(_10943_),
    .ZN(_10975_));
 NAND2_X1 _37050_ (.A1(_10974_),
    .A2(_10975_),
    .ZN(_00793_));
 AND2_X4 _37051_ (.A1(_10873_),
    .A2(_10935_),
    .ZN(_10976_));
 INV_X8 _37052_ (.A(_10976_),
    .ZN(_10977_));
 OAI211_X1 _37053_ (.A(\bp_fe_pc_gen_1.btb.v_r [40]),
    .B(_10949_),
    .C1(_10977_),
    .C2(_10964_),
    .ZN(_10978_));
 NAND4_X1 _37054_ (.A1(_10881_),
    .A2(_10925_),
    .A3(_10959_),
    .A4(_10943_),
    .ZN(_10979_));
 NAND2_X1 _37055_ (.A1(_10978_),
    .A2(_10979_),
    .ZN(_00792_));
 NAND2_X4 _37056_ (.A1(_10761_),
    .A2(_10766_),
    .ZN(_10980_));
 NOR2_X4 _37057_ (.A1(_10980_),
    .A2(_10771_),
    .ZN(_10981_));
 BUF_X8 _37058_ (.A(_10981_),
    .Z(_10982_));
 AND2_X4 _37059_ (.A1(net93),
    .A2(_10982_),
    .ZN(_10983_));
 INV_X16 _37060_ (.A(_10983_),
    .ZN(_10984_));
 OAI211_X1 _37061_ (.A(\bp_fe_pc_gen_1.btb.v_r [39]),
    .B(_10949_),
    .C1(_10984_),
    .C2(_10964_),
    .ZN(_10985_));
 BUF_X2 _37062_ (.A(_08722_),
    .Z(_10986_));
 BUF_X16 _37063_ (.A(_10981_),
    .Z(_10987_));
 BUF_X8 _37064_ (.A(_10987_),
    .Z(_10988_));
 BUF_X8 _37065_ (.A(_10988_),
    .Z(_10989_));
 BUF_X16 _37066_ (.A(_10989_),
    .Z(_10990_));
 BUF_X16 _37067_ (.A(_10990_),
    .Z(_10991_));
 NAND4_X1 _37068_ (.A1(_10806_),
    .A2(_10986_),
    .A3(_10959_),
    .A4(_10991_),
    .ZN(_10992_));
 NAND2_X1 _37069_ (.A1(_10985_),
    .A2(_10992_),
    .ZN(_00790_));
 AND2_X4 _37070_ (.A1(net83),
    .A2(_10981_),
    .ZN(_10993_));
 INV_X16 _37071_ (.A(_10993_),
    .ZN(_10994_));
 OAI211_X1 _37072_ (.A(\bp_fe_pc_gen_1.btb.v_r [38]),
    .B(_10949_),
    .C1(_10994_),
    .C2(_10964_),
    .ZN(_10995_));
 NAND4_X1 _37073_ (.A1(_10820_),
    .A2(_10986_),
    .A3(_10959_),
    .A4(_10991_),
    .ZN(_10996_));
 NAND2_X1 _37074_ (.A1(_10995_),
    .A2(_10996_),
    .ZN(_00789_));
 AND2_X4 _37075_ (.A1(net81),
    .A2(_10982_),
    .ZN(_10997_));
 INV_X16 _37076_ (.A(_10997_),
    .ZN(_10998_));
 OAI211_X1 _37077_ (.A(\bp_fe_pc_gen_1.btb.v_r [37]),
    .B(_10949_),
    .C1(_10998_),
    .C2(_10964_),
    .ZN(_10999_));
 NAND4_X1 _37078_ (.A1(_10833_),
    .A2(_10986_),
    .A3(_10959_),
    .A4(_10991_),
    .ZN(_11000_));
 NAND2_X1 _37079_ (.A1(_10999_),
    .A2(_11000_),
    .ZN(_00788_));
 AND2_X2 _37080_ (.A1(net71),
    .A2(_10982_),
    .ZN(_11001_));
 BUF_X16 _37081_ (.A(_11001_),
    .Z(_11002_));
 BUF_X16 _37082_ (.A(_11002_),
    .Z(_11003_));
 INV_X16 _37083_ (.A(_11003_),
    .ZN(_11004_));
 OAI211_X1 _37084_ (.A(\bp_fe_pc_gen_1.btb.v_r [36]),
    .B(_10949_),
    .C1(_11004_),
    .C2(_10964_),
    .ZN(_11005_));
 NAND4_X1 _37085_ (.A1(_10846_),
    .A2(_10986_),
    .A3(_10959_),
    .A4(_10991_),
    .ZN(_11006_));
 NAND2_X1 _37086_ (.A1(_11005_),
    .A2(_11006_),
    .ZN(_00787_));
 BUF_X4 _37087_ (.A(_08674_),
    .Z(_11007_));
 AND2_X4 _37088_ (.A1(_10757_),
    .A2(_10982_),
    .ZN(_11008_));
 INV_X16 _37089_ (.A(_11008_),
    .ZN(_11009_));
 OAI211_X1 _37090_ (.A(\bp_fe_pc_gen_1.btb.v_r [35]),
    .B(_11007_),
    .C1(_11009_),
    .C2(_10964_),
    .ZN(_11010_));
 NAND4_X1 _37091_ (.A1(_10782_),
    .A2(_10986_),
    .A3(_10959_),
    .A4(_10991_),
    .ZN(_11011_));
 NAND2_X1 _37092_ (.A1(_11010_),
    .A2(_11011_),
    .ZN(_00786_));
 AND2_X4 _37093_ (.A1(_10855_),
    .A2(_10987_),
    .ZN(_11012_));
 INV_X16 _37094_ (.A(_11012_),
    .ZN(_11013_));
 OAI211_X1 _37095_ (.A(\bp_fe_pc_gen_1.btb.v_r [34]),
    .B(_11007_),
    .C1(_11013_),
    .C2(_10964_),
    .ZN(_11014_));
 BUF_X32 _37096_ (.A(_10784_),
    .Z(_11015_));
 BUF_X2 _37097_ (.A(_11015_),
    .Z(_11016_));
 NAND4_X1 _37098_ (.A1(_10860_),
    .A2(_10986_),
    .A3(_11016_),
    .A4(_10991_),
    .ZN(_11017_));
 NAND2_X1 _37099_ (.A1(_11014_),
    .A2(_11017_),
    .ZN(_00785_));
 AND2_X2 _37100_ (.A1(net66),
    .A2(_10982_),
    .ZN(_11018_));
 BUF_X16 _37101_ (.A(_11018_),
    .Z(_11019_));
 INV_X16 _37102_ (.A(_11019_),
    .ZN(_11020_));
 BUF_X4 _37103_ (.A(_10775_),
    .Z(_11021_));
 OAI211_X1 _37104_ (.A(\bp_fe_pc_gen_1.btb.v_r [33]),
    .B(_11007_),
    .C1(_11020_),
    .C2(_11021_),
    .ZN(_11022_));
 NAND4_X1 _37105_ (.A1(_10870_),
    .A2(_10986_),
    .A3(_11016_),
    .A4(_10991_),
    .ZN(_11023_));
 NAND2_X1 _37106_ (.A1(_11022_),
    .A2(_11023_),
    .ZN(_00784_));
 AND2_X2 _37107_ (.A1(_10873_),
    .A2(_10982_),
    .ZN(_11024_));
 BUF_X16 _37108_ (.A(_11024_),
    .Z(_11025_));
 INV_X16 _37109_ (.A(_11025_),
    .ZN(_11026_));
 OAI211_X1 _37110_ (.A(\bp_fe_pc_gen_1.btb.v_r [32]),
    .B(_11007_),
    .C1(_11026_),
    .C2(_11021_),
    .ZN(_11027_));
 NAND4_X1 _37111_ (.A1(_10881_),
    .A2(_10986_),
    .A3(_11016_),
    .A4(_10991_),
    .ZN(_11028_));
 NAND2_X1 _37112_ (.A1(_11027_),
    .A2(_11028_),
    .ZN(_00783_));
 INV_X4 _37113_ (.A(_10771_),
    .ZN(_11029_));
 NOR2_X4 _37114_ (.A1(_10767_),
    .A2(_11029_),
    .ZN(_11030_));
 AND2_X4 _37115_ (.A1(net89),
    .A2(net101),
    .ZN(_11031_));
 INV_X32 _37116_ (.A(_11031_),
    .ZN(_11032_));
 OAI211_X1 _37117_ (.A(\bp_fe_pc_gen_1.btb.v_r [31]),
    .B(_11007_),
    .C1(_11032_),
    .C2(_11021_),
    .ZN(_11033_));
 BUF_X8 _37118_ (.A(net97),
    .Z(_11034_));
 BUF_X8 _37119_ (.A(_11034_),
    .Z(_11035_));
 BUF_X16 _37120_ (.A(_11035_),
    .Z(_11036_));
 BUF_X8 _37121_ (.A(_11036_),
    .Z(_11037_));
 BUF_X8 _37122_ (.A(_11037_),
    .Z(_11038_));
 BUF_X16 _37123_ (.A(_11038_),
    .Z(_11039_));
 NAND4_X1 _37124_ (.A1(_10806_),
    .A2(_10986_),
    .A3(_11016_),
    .A4(_11039_),
    .ZN(_11040_));
 NAND2_X1 _37125_ (.A1(_11033_),
    .A2(_11040_),
    .ZN(_00782_));
 AND2_X4 _37126_ (.A1(_10811_),
    .A2(net103),
    .ZN(_11041_));
 INV_X16 _37127_ (.A(_11041_),
    .ZN(_11042_));
 OAI211_X1 _37128_ (.A(\bp_fe_pc_gen_1.btb.v_r [30]),
    .B(_11007_),
    .C1(_11042_),
    .C2(_11021_),
    .ZN(_11043_));
 NAND4_X1 _37129_ (.A1(_10820_),
    .A2(_10986_),
    .A3(_11016_),
    .A4(_11039_),
    .ZN(_11044_));
 NAND2_X1 _37130_ (.A1(_11043_),
    .A2(_11044_),
    .ZN(_00781_));
 AND2_X4 _37131_ (.A1(_10901_),
    .A2(net98),
    .ZN(_11045_));
 INV_X16 _37132_ (.A(_11045_),
    .ZN(_11046_));
 OAI211_X1 _37133_ (.A(\bp_fe_pc_gen_1.btb.v_r [29]),
    .B(_11007_),
    .C1(_11046_),
    .C2(_11021_),
    .ZN(_11047_));
 BUF_X4 _37134_ (.A(_08722_),
    .Z(_11048_));
 NAND4_X1 _37135_ (.A1(_10833_),
    .A2(_11048_),
    .A3(_11016_),
    .A4(_11039_),
    .ZN(_11049_));
 NAND2_X1 _37136_ (.A1(_11047_),
    .A2(_11049_),
    .ZN(_00779_));
 AND2_X4 _37137_ (.A1(net76),
    .A2(net102),
    .ZN(_11050_));
 INV_X16 _37138_ (.A(_11050_),
    .ZN(_11051_));
 OAI211_X1 _37139_ (.A(\bp_fe_pc_gen_1.btb.v_r [28]),
    .B(_11007_),
    .C1(_11051_),
    .C2(_11021_),
    .ZN(_11052_));
 NAND4_X1 _37140_ (.A1(_10846_),
    .A2(_11048_),
    .A3(_11016_),
    .A4(_11039_),
    .ZN(_11053_));
 NAND2_X1 _37141_ (.A1(_11052_),
    .A2(_11053_),
    .ZN(_00778_));
 AND2_X4 _37142_ (.A1(_10757_),
    .A2(_11034_),
    .ZN(_11054_));
 INV_X16 _37143_ (.A(_11054_),
    .ZN(_11055_));
 OAI211_X1 _37144_ (.A(\bp_fe_pc_gen_1.btb.v_r [27]),
    .B(_11007_),
    .C1(_11055_),
    .C2(_11021_),
    .ZN(_11056_));
 NAND4_X1 _37145_ (.A1(_10782_),
    .A2(_11048_),
    .A3(_11016_),
    .A4(_11039_),
    .ZN(_11057_));
 NAND2_X1 _37146_ (.A1(_11056_),
    .A2(_11057_),
    .ZN(_00777_));
 AND2_X1 _37147_ (.A1(_10854_),
    .A2(net97),
    .ZN(_11058_));
 BUF_X8 _37148_ (.A(_11058_),
    .Z(_11059_));
 BUF_X16 _37149_ (.A(_11059_),
    .Z(_11060_));
 INV_X16 _37150_ (.A(_11060_),
    .ZN(_11061_));
 OAI211_X1 _37151_ (.A(\bp_fe_pc_gen_1.btb.v_r [26]),
    .B(_11007_),
    .C1(_11061_),
    .C2(_11021_),
    .ZN(_11062_));
 NAND4_X1 _37152_ (.A1(_10860_),
    .A2(_11048_),
    .A3(_11016_),
    .A4(_11039_),
    .ZN(_11063_));
 NAND2_X1 _37153_ (.A1(_11062_),
    .A2(_11063_),
    .ZN(_00776_));
 BUF_X4 _37154_ (.A(_08674_),
    .Z(_11064_));
 AND2_X4 _37155_ (.A1(net68),
    .A2(net100),
    .ZN(_11065_));
 INV_X16 _37156_ (.A(_11065_),
    .ZN(_11066_));
 OAI211_X1 _37157_ (.A(\bp_fe_pc_gen_1.btb.v_r [25]),
    .B(_11064_),
    .C1(_11066_),
    .C2(_11021_),
    .ZN(_11067_));
 NAND4_X1 _37158_ (.A1(_10870_),
    .A2(_11048_),
    .A3(_11016_),
    .A4(_11039_),
    .ZN(_11068_));
 NAND2_X1 _37159_ (.A1(_11067_),
    .A2(_11068_),
    .ZN(_00775_));
 AND2_X4 _37160_ (.A1(net62),
    .A2(net99),
    .ZN(_11069_));
 INV_X16 _37161_ (.A(_11069_),
    .ZN(_11070_));
 OAI211_X1 _37162_ (.A(\bp_fe_pc_gen_1.btb.v_r [24]),
    .B(_11064_),
    .C1(_11070_),
    .C2(_11021_),
    .ZN(_11071_));
 BUF_X4 _37163_ (.A(_11015_),
    .Z(_11072_));
 NAND4_X1 _37164_ (.A1(_10881_),
    .A2(_11048_),
    .A3(_11072_),
    .A4(_11039_),
    .ZN(_11073_));
 NAND2_X1 _37165_ (.A1(_11071_),
    .A2(_11073_),
    .ZN(_00774_));
 NOR2_X4 _37166_ (.A1(_10884_),
    .A2(_11029_),
    .ZN(_11074_));
 AND2_X4 _37167_ (.A1(net90),
    .A2(net96),
    .ZN(_11075_));
 INV_X16 _37168_ (.A(_11075_),
    .ZN(_11076_));
 BUF_X4 _37169_ (.A(_10775_),
    .Z(_11077_));
 OAI211_X1 _37170_ (.A(\bp_fe_pc_gen_1.btb.v_r [23]),
    .B(_11064_),
    .C1(_11076_),
    .C2(_11077_),
    .ZN(_11078_));
 BUF_X16 _37171_ (.A(net94),
    .Z(_11079_));
 BUF_X8 _37172_ (.A(_11079_),
    .Z(_11080_));
 BUF_X8 _37173_ (.A(_11080_),
    .Z(_11081_));
 BUF_X8 _37174_ (.A(_11081_),
    .Z(_11082_));
 BUF_X16 _37175_ (.A(_11082_),
    .Z(_11083_));
 NAND4_X1 _37176_ (.A1(_10806_),
    .A2(_11048_),
    .A3(_11072_),
    .A4(_11083_),
    .ZN(_11084_));
 NAND2_X1 _37177_ (.A1(_11078_),
    .A2(_11084_),
    .ZN(_00773_));
 AND2_X4 _37178_ (.A1(net87),
    .A2(net95),
    .ZN(_11085_));
 INV_X16 _37179_ (.A(_11085_),
    .ZN(_11086_));
 OAI211_X1 _37180_ (.A(\bp_fe_pc_gen_1.btb.v_r [22]),
    .B(_11064_),
    .C1(_11086_),
    .C2(_11077_),
    .ZN(_11087_));
 NAND4_X1 _37181_ (.A1(_10820_),
    .A2(_11048_),
    .A3(_11072_),
    .A4(_11083_),
    .ZN(_11088_));
 NAND2_X1 _37182_ (.A1(_11087_),
    .A2(_11088_),
    .ZN(_00772_));
 BUF_X8 _37183_ (.A(net94),
    .Z(_11089_));
 AND2_X4 _37184_ (.A1(_10901_),
    .A2(_11089_),
    .ZN(_11090_));
 INV_X16 _37185_ (.A(_11090_),
    .ZN(_11091_));
 OAI211_X1 _37186_ (.A(\bp_fe_pc_gen_1.btb.v_r [21]),
    .B(_11064_),
    .C1(_11091_),
    .C2(_11077_),
    .ZN(_11092_));
 NAND4_X1 _37187_ (.A1(_10833_),
    .A2(_11048_),
    .A3(_11072_),
    .A4(_11083_),
    .ZN(_11093_));
 NAND2_X1 _37188_ (.A1(_11092_),
    .A2(_11093_),
    .ZN(_00771_));
 AND2_X4 _37189_ (.A1(net74),
    .A2(_11089_),
    .ZN(_11094_));
 INV_X2 _37190_ (.A(_11094_),
    .ZN(_11095_));
 BUF_X16 _37191_ (.A(_11095_),
    .Z(_11096_));
 OAI211_X1 _37192_ (.A(\bp_fe_pc_gen_1.btb.v_r [20]),
    .B(_11064_),
    .C1(_11096_),
    .C2(_11077_),
    .ZN(_11097_));
 NAND4_X1 _37193_ (.A1(_10846_),
    .A2(_11048_),
    .A3(_11072_),
    .A4(_11083_),
    .ZN(_11098_));
 NAND2_X1 _37194_ (.A1(_11097_),
    .A2(_11098_),
    .ZN(_00770_));
 AND2_X4 _37195_ (.A1(net111),
    .A2(_11089_),
    .ZN(_11099_));
 BUF_X16 _37196_ (.A(_11099_),
    .Z(_11100_));
 INV_X16 _37197_ (.A(_11100_),
    .ZN(_11101_));
 OAI211_X1 _37198_ (.A(\bp_fe_pc_gen_1.btb.v_r [19]),
    .B(_11064_),
    .C1(_11101_),
    .C2(_11077_),
    .ZN(_11102_));
 BUF_X4 _37199_ (.A(_08722_),
    .Z(_11103_));
 NAND4_X1 _37200_ (.A1(_10782_),
    .A2(_11103_),
    .A3(_11072_),
    .A4(_11083_),
    .ZN(_11104_));
 NAND2_X1 _37201_ (.A1(_11102_),
    .A2(_11104_),
    .ZN(_00768_));
 AND2_X4 _37202_ (.A1(_10854_),
    .A2(net94),
    .ZN(_11105_));
 BUF_X8 _37203_ (.A(_11105_),
    .Z(_11106_));
 INV_X16 _37204_ (.A(_11106_),
    .ZN(_11107_));
 OAI211_X1 _37205_ (.A(\bp_fe_pc_gen_1.btb.v_r [18]),
    .B(_11064_),
    .C1(_11107_),
    .C2(_11077_),
    .ZN(_11108_));
 NAND4_X1 _37206_ (.A1(_10860_),
    .A2(_11103_),
    .A3(_11072_),
    .A4(_11083_),
    .ZN(_11109_));
 NAND2_X1 _37207_ (.A1(_11108_),
    .A2(_11109_),
    .ZN(_00767_));
 AND2_X4 _37208_ (.A1(_10920_),
    .A2(_11079_),
    .ZN(_11110_));
 INV_X16 _37209_ (.A(_11110_),
    .ZN(_11111_));
 OAI211_X1 _37210_ (.A(\bp_fe_pc_gen_1.btb.v_r [17]),
    .B(_11064_),
    .C1(_11111_),
    .C2(_11077_),
    .ZN(_11112_));
 NAND4_X1 _37211_ (.A1(_10870_),
    .A2(_11103_),
    .A3(_11072_),
    .A4(_11083_),
    .ZN(_11113_));
 NAND2_X1 _37212_ (.A1(_11112_),
    .A2(_11113_),
    .ZN(_00766_));
 AND2_X4 _37213_ (.A1(_10873_),
    .A2(_11089_),
    .ZN(_11114_));
 INV_X16 _37214_ (.A(_11114_),
    .ZN(_11115_));
 OAI211_X1 _37215_ (.A(\bp_fe_pc_gen_1.btb.v_r [16]),
    .B(_11064_),
    .C1(_11115_),
    .C2(_11077_),
    .ZN(_11116_));
 NAND4_X1 _37216_ (.A1(_10881_),
    .A2(_11103_),
    .A3(_11072_),
    .A4(_11083_),
    .ZN(_11117_));
 NAND2_X1 _37217_ (.A1(_11116_),
    .A2(_11117_),
    .ZN(_00765_));
 BUF_X4 _37218_ (.A(_08722_),
    .Z(_11118_));
 NOR2_X4 _37219_ (.A1(_10933_),
    .A2(_11029_),
    .ZN(_11119_));
 AND2_X4 _37220_ (.A1(net89),
    .A2(_11119_),
    .ZN(_11120_));
 INV_X16 _37221_ (.A(_11120_),
    .ZN(_11121_));
 OAI211_X1 _37222_ (.A(\bp_fe_pc_gen_1.btb.v_r [15]),
    .B(_11118_),
    .C1(_11121_),
    .C2(_11077_),
    .ZN(_11122_));
 BUF_X8 _37223_ (.A(_11119_),
    .Z(_11123_));
 BUF_X16 _37224_ (.A(_11123_),
    .Z(_11124_));
 BUF_X16 _37225_ (.A(_11124_),
    .Z(_11125_));
 BUF_X16 _37226_ (.A(_11125_),
    .Z(_11126_));
 BUF_X16 _37227_ (.A(_11126_),
    .Z(_11127_));
 BUF_X16 _37228_ (.A(_11127_),
    .Z(_11128_));
 NAND4_X1 _37229_ (.A1(_10806_),
    .A2(_11103_),
    .A3(_11072_),
    .A4(_11128_),
    .ZN(_11129_));
 NAND2_X1 _37230_ (.A1(_11122_),
    .A2(_11129_),
    .ZN(_00764_));
 AND2_X2 _37231_ (.A1(net87),
    .A2(_11119_),
    .ZN(_11130_));
 BUF_X16 _37232_ (.A(_11130_),
    .Z(_11131_));
 INV_X16 _37233_ (.A(_11131_),
    .ZN(_11132_));
 OAI211_X1 _37234_ (.A(\bp_fe_pc_gen_1.btb.v_r [14]),
    .B(_11118_),
    .C1(_11132_),
    .C2(_11077_),
    .ZN(_11133_));
 BUF_X2 _37235_ (.A(_11015_),
    .Z(_11134_));
 NAND4_X1 _37236_ (.A1(_10820_),
    .A2(_11103_),
    .A3(_11134_),
    .A4(_11128_),
    .ZN(_11135_));
 NAND2_X1 _37237_ (.A1(_11133_),
    .A2(_11135_),
    .ZN(_00763_));
 AND2_X4 _37238_ (.A1(net80),
    .A2(_11123_),
    .ZN(_11136_));
 INV_X16 _37239_ (.A(_11136_),
    .ZN(_11137_));
 BUF_X4 _37240_ (.A(_10775_),
    .Z(_11138_));
 OAI211_X1 _37241_ (.A(\bp_fe_pc_gen_1.btb.v_r [13]),
    .B(_11118_),
    .C1(_11137_),
    .C2(_11138_),
    .ZN(_11139_));
 NAND4_X1 _37242_ (.A1(_10833_),
    .A2(_11103_),
    .A3(_11134_),
    .A4(_11128_),
    .ZN(_11140_));
 NAND2_X1 _37243_ (.A1(_11139_),
    .A2(_11140_),
    .ZN(_00762_));
 AND2_X4 _37244_ (.A1(net75),
    .A2(_11123_),
    .ZN(_11141_));
 INV_X16 _37245_ (.A(_11141_),
    .ZN(_11142_));
 OAI211_X1 _37246_ (.A(\bp_fe_pc_gen_1.btb.v_r [12]),
    .B(_11118_),
    .C1(_11142_),
    .C2(_11138_),
    .ZN(_11143_));
 NAND4_X1 _37247_ (.A1(_10846_),
    .A2(_11103_),
    .A3(_11134_),
    .A4(_11128_),
    .ZN(_11144_));
 NAND2_X1 _37248_ (.A1(_11143_),
    .A2(_11144_),
    .ZN(_00761_));
 BUF_X8 _37249_ (.A(_11119_),
    .Z(_11145_));
 AND2_X4 _37250_ (.A1(_10778_),
    .A2(_11145_),
    .ZN(_11146_));
 BUF_X16 _37251_ (.A(_11146_),
    .Z(_11147_));
 INV_X8 _37252_ (.A(_11147_),
    .ZN(_11148_));
 OAI211_X1 _37253_ (.A(\bp_fe_pc_gen_1.btb.v_r [11]),
    .B(_11118_),
    .C1(_11148_),
    .C2(_11138_),
    .ZN(_11149_));
 NAND4_X1 _37254_ (.A1(_10782_),
    .A2(_11103_),
    .A3(_11134_),
    .A4(_11128_),
    .ZN(_11150_));
 NAND2_X1 _37255_ (.A1(_11149_),
    .A2(_11150_),
    .ZN(_00760_));
 AND2_X4 _37256_ (.A1(_10854_),
    .A2(_11123_),
    .ZN(_11151_));
 BUF_X16 _37257_ (.A(_11151_),
    .Z(_11152_));
 BUF_X16 _37258_ (.A(_11152_),
    .Z(_11153_));
 INV_X16 _37259_ (.A(_11153_),
    .ZN(_11154_));
 OAI211_X1 _37260_ (.A(\bp_fe_pc_gen_1.btb.v_r [10]),
    .B(_11118_),
    .C1(_11154_),
    .C2(_11138_),
    .ZN(_11155_));
 NAND4_X1 _37261_ (.A1(_10860_),
    .A2(_11103_),
    .A3(_11134_),
    .A4(_11128_),
    .ZN(_11156_));
 NAND2_X1 _37262_ (.A1(_11155_),
    .A2(_11156_),
    .ZN(_00759_));
 AND2_X2 _37263_ (.A1(_10920_),
    .A2(_11123_),
    .ZN(_11157_));
 BUF_X16 _37264_ (.A(_11157_),
    .Z(_11158_));
 BUF_X32 _37265_ (.A(_11158_),
    .Z(_11159_));
 INV_X1 _37266_ (.A(_11159_),
    .ZN(_11160_));
 OAI211_X1 _37267_ (.A(\bp_fe_pc_gen_1.btb.v_r [9]),
    .B(_11118_),
    .C1(_11160_),
    .C2(_11138_),
    .ZN(_11161_));
 BUF_X2 _37268_ (.A(_08722_),
    .Z(_11162_));
 NAND4_X1 _37269_ (.A1(_10870_),
    .A2(_11162_),
    .A3(_11134_),
    .A4(_11128_),
    .ZN(_11163_));
 NAND2_X1 _37270_ (.A1(_11161_),
    .A2(_11163_),
    .ZN(_00821_));
 AND2_X4 _37271_ (.A1(_10873_),
    .A2(_11123_),
    .ZN(_11164_));
 INV_X16 _37272_ (.A(_11164_),
    .ZN(_11165_));
 OAI211_X1 _37273_ (.A(\bp_fe_pc_gen_1.btb.v_r [8]),
    .B(_11118_),
    .C1(_11165_),
    .C2(_11138_),
    .ZN(_11166_));
 NAND4_X1 _37274_ (.A1(_10881_),
    .A2(_11162_),
    .A3(_11134_),
    .A4(_11128_),
    .ZN(_11167_));
 NAND2_X1 _37275_ (.A1(_11166_),
    .A2(_11167_),
    .ZN(_00820_));
 NOR2_X4 _37276_ (.A1(_10980_),
    .A2(_11029_),
    .ZN(_11168_));
 AND2_X2 _37277_ (.A1(net88),
    .A2(_11168_),
    .ZN(_11169_));
 BUF_X16 _37278_ (.A(_11169_),
    .Z(_11170_));
 INV_X8 _37279_ (.A(_11170_),
    .ZN(_11171_));
 OAI211_X1 _37280_ (.A(\bp_fe_pc_gen_1.btb.v_r [7]),
    .B(_11118_),
    .C1(_11171_),
    .C2(_11138_),
    .ZN(_11172_));
 BUF_X8 _37281_ (.A(_11168_),
    .Z(_11173_));
 BUF_X16 _37282_ (.A(_11173_),
    .Z(_11174_));
 BUF_X16 _37283_ (.A(_11174_),
    .Z(_11175_));
 BUF_X8 _37284_ (.A(_11175_),
    .Z(_11176_));
 BUF_X4 _37285_ (.A(_11176_),
    .Z(_11177_));
 BUF_X8 _37286_ (.A(_11177_),
    .Z(_11178_));
 NAND4_X1 _37287_ (.A1(_10806_),
    .A2(_11162_),
    .A3(_11134_),
    .A4(_11178_),
    .ZN(_11179_));
 NAND2_X1 _37288_ (.A1(_11172_),
    .A2(_11179_),
    .ZN(_00819_));
 AND2_X1 _37289_ (.A1(net85),
    .A2(_11168_),
    .ZN(_11180_));
 BUF_X8 _37290_ (.A(_11180_),
    .Z(_11181_));
 INV_X8 _37291_ (.A(_11181_),
    .ZN(_11182_));
 OAI211_X1 _37292_ (.A(\bp_fe_pc_gen_1.btb.v_r [6]),
    .B(_11118_),
    .C1(_11182_),
    .C2(_11138_),
    .ZN(_11183_));
 NAND4_X1 _37293_ (.A1(_10820_),
    .A2(_11162_),
    .A3(_11134_),
    .A4(_11178_),
    .ZN(_11184_));
 NAND2_X1 _37294_ (.A1(_11183_),
    .A2(_11184_),
    .ZN(_00818_));
 BUF_X8 _37295_ (.A(_11168_),
    .Z(_11185_));
 AND2_X4 _37296_ (.A1(_10901_),
    .A2(_11185_),
    .ZN(_11186_));
 INV_X16 _37297_ (.A(_11186_),
    .ZN(_11187_));
 OAI211_X1 _37298_ (.A(\bp_fe_pc_gen_1.btb.v_r [5]),
    .B(_10783_),
    .C1(_11187_),
    .C2(_11138_),
    .ZN(_11188_));
 NAND4_X1 _37299_ (.A1(_10833_),
    .A2(_11162_),
    .A3(_11134_),
    .A4(_11178_),
    .ZN(_11189_));
 NAND2_X1 _37300_ (.A1(_11188_),
    .A2(_11189_),
    .ZN(_00813_));
 AND2_X4 _37301_ (.A1(_10842_),
    .A2(_11173_),
    .ZN(_11190_));
 INV_X8 _37302_ (.A(_11190_),
    .ZN(_11191_));
 OAI211_X1 _37303_ (.A(\bp_fe_pc_gen_1.btb.v_r [4]),
    .B(_10783_),
    .C1(_11191_),
    .C2(_11138_),
    .ZN(_11192_));
 BUF_X8 _37304_ (.A(_11015_),
    .Z(_11193_));
 NAND4_X2 _37305_ (.A1(_10846_),
    .A2(_11162_),
    .A3(_11193_),
    .A4(_11178_),
    .ZN(_11194_));
 NAND2_X1 _37306_ (.A1(_11192_),
    .A2(_11194_),
    .ZN(_00802_));
 AND2_X4 _37307_ (.A1(_10757_),
    .A2(_11173_),
    .ZN(_11195_));
 BUF_X16 _37308_ (.A(_11195_),
    .Z(_11196_));
 INV_X8 _37309_ (.A(_11196_),
    .ZN(_11197_));
 OAI211_X1 _37310_ (.A(\bp_fe_pc_gen_1.btb.v_r [3]),
    .B(_10783_),
    .C1(_11197_),
    .C2(_10775_),
    .ZN(_11198_));
 NAND4_X1 _37311_ (.A1(_10782_),
    .A2(_11162_),
    .A3(_11193_),
    .A4(_11178_),
    .ZN(_11199_));
 NAND2_X1 _37312_ (.A1(_11198_),
    .A2(_11199_),
    .ZN(_00791_));
 AND2_X4 _37313_ (.A1(_10854_),
    .A2(_11185_),
    .ZN(_11200_));
 INV_X16 _37314_ (.A(_11200_),
    .ZN(_11201_));
 OAI211_X1 _37315_ (.A(\bp_fe_pc_gen_1.btb.v_r [2]),
    .B(_10783_),
    .C1(_11201_),
    .C2(_10775_),
    .ZN(_11202_));
 NAND4_X1 _37316_ (.A1(_10860_),
    .A2(_11162_),
    .A3(_11193_),
    .A4(_11178_),
    .ZN(_11203_));
 NAND2_X1 _37317_ (.A1(_11202_),
    .A2(_11203_),
    .ZN(_00780_));
 AND2_X1 _37318_ (.A1(net62),
    .A2(_11185_),
    .ZN(_11204_));
 BUF_X8 _37319_ (.A(_11204_),
    .Z(_11205_));
 BUF_X16 _37320_ (.A(_11205_),
    .Z(_11206_));
 INV_X8 _37321_ (.A(_11206_),
    .ZN(_11207_));
 OAI211_X1 _37322_ (.A(\bp_fe_pc_gen_1.btb.v_r [0]),
    .B(_10783_),
    .C1(_11207_),
    .C2(_10775_),
    .ZN(_11208_));
 NAND4_X1 _37323_ (.A1(_10881_),
    .A2(_11162_),
    .A3(_11193_),
    .A4(_11178_),
    .ZN(_11209_));
 NAND2_X1 _37324_ (.A1(_11208_),
    .A2(_11209_),
    .ZN(_00758_));
 AND2_X2 _37325_ (.A1(net64),
    .A2(_11185_),
    .ZN(_11210_));
 BUF_X16 _37326_ (.A(_11210_),
    .Z(_11211_));
 INV_X8 _37327_ (.A(_11211_),
    .ZN(_11212_));
 OAI211_X1 _37328_ (.A(\bp_fe_pc_gen_1.btb.v_r [1]),
    .B(_10783_),
    .C1(_11212_),
    .C2(_10775_),
    .ZN(_11213_));
 NAND4_X2 _37329_ (.A1(_10870_),
    .A2(_11162_),
    .A3(_11193_),
    .A4(_11178_),
    .ZN(_11214_));
 NAND2_X1 _37330_ (.A1(_11213_),
    .A2(_11214_),
    .ZN(_00769_));
 NOR2_X4 _37331_ (.A1(_10740_),
    .A2(_08743_),
    .ZN(_11215_));
 NOR2_X1 _37332_ (.A1(_11215_),
    .A2(_08999_),
    .ZN(\bp_fe_pc_gen_1.btb.N160 ));
 AOI21_X2 _37333_ (.A(_09000_),
    .B1(_08475_),
    .B2(_08478_),
    .ZN(\bp_fe_pc_gen_1.btb.N161 ));
 NOR2_X1 _37334_ (.A1(_08755_),
    .A2(_08999_),
    .ZN(\bp_fe_pc_gen_1.btb.N162 ));
 NOR2_X1 _37335_ (.A1(_08757_),
    .A2(_08999_),
    .ZN(\bp_fe_pc_gen_1.btb.N163 ));
 NOR2_X1 _37336_ (.A1(_08759_),
    .A2(_08999_),
    .ZN(\bp_fe_pc_gen_1.btb.N164 ));
 NOR2_X2 _37337_ (.A1(_08762_),
    .A2(_08999_),
    .ZN(\bp_fe_pc_gen_1.btb.N165 ));
 NOR2_X1 _37338_ (.A1(_08764_),
    .A2(_08999_),
    .ZN(\bp_fe_pc_gen_1.btb.N150 ));
 NOR2_X2 _37339_ (.A1(_08384_),
    .A2(_08388_),
    .ZN(_11216_));
 NOR2_X1 _37340_ (.A1(_11216_),
    .A2(_08999_),
    .ZN(\bp_fe_pc_gen_1.btb.N151 ));
 NOR2_X1 _37341_ (.A1(_08767_),
    .A2(_08999_),
    .ZN(\bp_fe_pc_gen_1.btb.N152 ));
 NOR2_X1 _37342_ (.A1(_08769_),
    .A2(_09000_),
    .ZN(\bp_fe_pc_gen_1.btb.N153 ));
 NOR2_X1 _37343_ (.A1(_08784_),
    .A2(_09000_),
    .ZN(\bp_fe_pc_gen_1.btb.N154 ));
 NOR2_X1 _37344_ (.A1(_10077_),
    .A2(_09000_),
    .ZN(\bp_fe_pc_gen_1.btb.N155 ));
 AOI21_X1 _37345_ (.A(_08651_),
    .B1(net212),
    .B2(_08803_),
    .ZN(\bp_fe_pc_gen_1.btb.N156 ));
 NOR2_X1 _37346_ (.A1(_10033_),
    .A2(_09000_),
    .ZN(\bp_fe_pc_gen_1.btb.N157 ));
 NOR2_X1 _37347_ (.A1(_08822_),
    .A2(_09000_),
    .ZN(\bp_fe_pc_gen_1.btb.N158 ));
 NOR2_X1 _37348_ (.A1(_10100_),
    .A2(_09000_),
    .ZN(\bp_fe_pc_gen_1.btb.N159 ));
 NOR4_X1 _37349_ (.A1(_08026_),
    .A2(_08651_),
    .A3(_08035_),
    .A4(_10786_),
    .ZN(\bp_fe_pc_gen_1.btb.N149 ));
 BUF_X4 _37350_ (.A(_08648_),
    .Z(_11217_));
 BUF_X4 _37351_ (.A(_08649_),
    .Z(_11218_));
 AOI211_X1 _37352_ (.A(_08957_),
    .B(_09005_),
    .C1(_11217_),
    .C2(_11218_),
    .ZN(_00731_));
 AOI211_X1 _37353_ (.A(_08957_),
    .B(_09010_),
    .C1(_11217_),
    .C2(_11218_),
    .ZN(_00742_));
 AOI211_X1 _37354_ (.A(_08957_),
    .B(_09011_),
    .C1(_11217_),
    .C2(_11218_),
    .ZN(_00750_));
 AOI211_X1 _37355_ (.A(_08957_),
    .B(_09012_),
    .C1(_11217_),
    .C2(_11218_),
    .ZN(_00751_));
 BUF_X4 _37356_ (.A(_08650_),
    .Z(_11219_));
 AOI211_X1 _37357_ (.A(_11219_),
    .B(_09013_),
    .C1(_11217_),
    .C2(_11218_),
    .ZN(_00752_));
 AOI211_X1 _37358_ (.A(_11219_),
    .B(_09014_),
    .C1(_11217_),
    .C2(_11218_),
    .ZN(_00753_));
 AOI211_X1 _37359_ (.A(_11219_),
    .B(_09015_),
    .C1(_11217_),
    .C2(_11218_),
    .ZN(_00754_));
 AOI211_X1 _37360_ (.A(_11219_),
    .B(_09016_),
    .C1(_11217_),
    .C2(_11218_),
    .ZN(_00755_));
 AOI211_X1 _37361_ (.A(_11219_),
    .B(_09017_),
    .C1(_11217_),
    .C2(_11218_),
    .ZN(_00756_));
 AOI211_X1 _37362_ (.A(_11219_),
    .B(_09018_),
    .C1(_11217_),
    .C2(_11218_),
    .ZN(_00757_));
 AOI211_X1 _37363_ (.A(_11219_),
    .B(_09019_),
    .C1(_08648_),
    .C2(_08649_),
    .ZN(_00732_));
 OR2_X4 _37364_ (.A1(fe_queue_v_o),
    .A2(_08516_),
    .ZN(_11220_));
 BUF_X4 _37365_ (.A(_11220_),
    .Z(_11221_));
 INV_X1 _37366_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [11]),
    .ZN(_11222_));
 NAND2_X4 _37367_ (.A1(fe_queue_v_o),
    .A2(_08674_),
    .ZN(_11223_));
 OAI22_X1 _37368_ (.A1(_11221_),
    .A2(_09022_),
    .B1(_11222_),
    .B2(_11223_),
    .ZN(_00733_));
 INV_X1 _37369_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [12]),
    .ZN(_11224_));
 OAI22_X1 _37370_ (.A1(_11221_),
    .A2(_09023_),
    .B1(_11224_),
    .B2(_11223_),
    .ZN(_00734_));
 INV_X1 _37371_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [13]),
    .ZN(_11225_));
 OAI22_X1 _37372_ (.A1(_11221_),
    .A2(_09024_),
    .B1(_11225_),
    .B2(_11223_),
    .ZN(_00735_));
 INV_X1 _37373_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [14]),
    .ZN(_11226_));
 OAI22_X1 _37374_ (.A1(_11221_),
    .A2(_09025_),
    .B1(_11226_),
    .B2(_11223_),
    .ZN(_00736_));
 INV_X1 _37375_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [15]),
    .ZN(_11227_));
 OAI22_X1 _37376_ (.A1(_11220_),
    .A2(_09026_),
    .B1(_11227_),
    .B2(_11223_),
    .ZN(_00737_));
 INV_X1 _37377_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [16]),
    .ZN(_11228_));
 OAI22_X1 _37378_ (.A1(_11220_),
    .A2(_09027_),
    .B1(_11228_),
    .B2(_11223_),
    .ZN(_00738_));
 INV_X1 _37379_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [17]),
    .ZN(_11229_));
 OAI22_X1 _37380_ (.A1(_11220_),
    .A2(_09028_),
    .B1(_11229_),
    .B2(_11223_),
    .ZN(_00739_));
 INV_X1 _37381_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [18]),
    .ZN(_11230_));
 OAI22_X1 _37382_ (.A1(_11220_),
    .A2(_09029_),
    .B1(_11230_),
    .B2(_11223_),
    .ZN(_00740_));
 INV_X1 _37383_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [19]),
    .ZN(_11231_));
 OAI22_X1 _37384_ (.A1(_11220_),
    .A2(_09030_),
    .B1(_11231_),
    .B2(_11223_),
    .ZN(_00741_));
 INV_X1 _37385_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [20]),
    .ZN(_11232_));
 OAI22_X1 _37386_ (.A1(_11220_),
    .A2(_09031_),
    .B1(_11232_),
    .B2(_11223_),
    .ZN(_00743_));
 NAND4_X1 _37387_ (.A1(_08648_),
    .A2(_08649_),
    .A3(_08727_),
    .A4(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [21]),
    .ZN(_11233_));
 OAI21_X1 _37388_ (.A(_11233_),
    .B1(_11221_),
    .B2(_09032_),
    .ZN(_00744_));
 NAND4_X1 _37389_ (.A1(_08648_),
    .A2(_08649_),
    .A3(_08727_),
    .A4(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [22]),
    .ZN(_11234_));
 OAI21_X1 _37390_ (.A(_11234_),
    .B1(_11221_),
    .B2(_09033_),
    .ZN(_00745_));
 NAND4_X1 _37391_ (.A1(_08648_),
    .A2(_08649_),
    .A3(_08727_),
    .A4(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [23]),
    .ZN(_11235_));
 OAI21_X1 _37392_ (.A(_11235_),
    .B1(_11221_),
    .B2(_09034_),
    .ZN(_00746_));
 NAND4_X1 _37393_ (.A1(_08648_),
    .A2(_08649_),
    .A3(_08727_),
    .A4(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [24]),
    .ZN(_11236_));
 OAI21_X1 _37394_ (.A(_11236_),
    .B1(_11221_),
    .B2(_09035_),
    .ZN(_00747_));
 NAND4_X1 _37395_ (.A1(_08648_),
    .A2(_08649_),
    .A3(_08727_),
    .A4(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [25]),
    .ZN(_11237_));
 OAI21_X1 _37396_ (.A(_11237_),
    .B1(_11221_),
    .B2(_09036_),
    .ZN(_00748_));
 NAND4_X1 _37397_ (.A1(_08648_),
    .A2(_08649_),
    .A3(_08727_),
    .A4(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [26]),
    .ZN(_11238_));
 OAI21_X1 _37398_ (.A(_11238_),
    .B1(_11221_),
    .B2(_09037_),
    .ZN(_00749_));
 BUF_X32 _37399_ (.A(_08447_),
    .Z(_11239_));
 BUF_X8 _37400_ (.A(_11239_),
    .Z(_11240_));
 BUF_X16 _37401_ (.A(_08427_),
    .Z(_11241_));
 BUF_X16 _37402_ (.A(_11241_),
    .Z(_11242_));
 MUX2_X1 _37403_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [6]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [524]),
    .S(_11242_),
    .Z(_11243_));
 BUF_X16 _37404_ (.A(_08426_),
    .Z(_11244_));
 BUF_X16 _37405_ (.A(_11244_),
    .Z(_11245_));
 AND2_X4 _37406_ (.A1(_11243_),
    .A2(_11245_),
    .ZN(_11246_));
 NAND2_X1 _37407_ (.A1(_08491_),
    .A2(_11246_),
    .ZN(_11247_));
 BUF_X16 _37408_ (.A(_08428_),
    .Z(_11248_));
 MUX2_X1 _37409_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [70]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [588]),
    .S(_11248_),
    .Z(_11249_));
 AND2_X4 _37410_ (.A1(_11249_),
    .A2(_08501_),
    .ZN(_11250_));
 BUF_X32 _37411_ (.A(_08483_),
    .Z(_11251_));
 BUF_X4 _37412_ (.A(_11251_),
    .Z(_11252_));
 BUF_X32 _37413_ (.A(_08487_),
    .Z(_11253_));
 BUF_X4 _37414_ (.A(_11253_),
    .Z(_11254_));
 OAI21_X1 _37415_ (.A(_11250_),
    .B1(_11252_),
    .B2(_11254_),
    .ZN(_11255_));
 AOI21_X1 _37416_ (.A(_11240_),
    .B1(_11247_),
    .B2(_11255_),
    .ZN(_11256_));
 BUF_X16 _37417_ (.A(_08446_),
    .Z(_11257_));
 BUF_X8 _37418_ (.A(_11257_),
    .Z(_11258_));
 BUF_X4 _37419_ (.A(_08490_),
    .Z(_11259_));
 MUX2_X1 _37420_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [134]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [652]),
    .S(_11248_),
    .Z(_11260_));
 AND2_X4 _37421_ (.A1(_11260_),
    .A2(_08501_),
    .ZN(_11261_));
 NAND2_X1 _37422_ (.A1(_11259_),
    .A2(_11261_),
    .ZN(_11262_));
 BUF_X32 _37423_ (.A(_08427_),
    .Z(_11263_));
 BUF_X16 _37424_ (.A(_11263_),
    .Z(_11264_));
 MUX2_X1 _37425_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [198]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [716]),
    .S(_11264_),
    .Z(_11265_));
 BUF_X16 _37426_ (.A(_08426_),
    .Z(_11266_));
 BUF_X4 _37427_ (.A(_11266_),
    .Z(_11267_));
 AND2_X1 _37428_ (.A1(_11265_),
    .A2(_11267_),
    .ZN(_11268_));
 BUF_X16 _37429_ (.A(_08483_),
    .Z(_11269_));
 BUF_X4 _37430_ (.A(_11269_),
    .Z(_11270_));
 BUF_X16 _37431_ (.A(_08487_),
    .Z(_11271_));
 BUF_X4 _37432_ (.A(_11271_),
    .Z(_11272_));
 OAI21_X1 _37433_ (.A(_11268_),
    .B1(_11270_),
    .B2(_11272_),
    .ZN(_11273_));
 AOI21_X1 _37434_ (.A(_11258_),
    .B1(_11262_),
    .B2(_11273_),
    .ZN(_11274_));
 OR2_X1 _37435_ (.A1(_11256_),
    .A2(_11274_),
    .ZN(_11275_));
 BUF_X16 _37436_ (.A(_11263_),
    .Z(_11276_));
 MUX2_X2 _37437_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [262]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [780]),
    .S(_11276_),
    .Z(_11277_));
 AND2_X1 _37438_ (.A1(_11277_),
    .A2(_11267_),
    .ZN(_11278_));
 NAND2_X1 _37439_ (.A1(_11259_),
    .A2(_11278_),
    .ZN(_11279_));
 MUX2_X2 _37440_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [326]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [844]),
    .S(_11276_),
    .Z(_11280_));
 AND2_X1 _37441_ (.A1(_11280_),
    .A2(_11267_),
    .ZN(_11281_));
 OAI21_X1 _37442_ (.A(_11281_),
    .B1(_11270_),
    .B2(_11272_),
    .ZN(_11282_));
 AOI21_X1 _37443_ (.A(_08448_),
    .B1(_11279_),
    .B2(_11282_),
    .ZN(_11283_));
 MUX2_X2 _37444_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [390]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [908]),
    .S(_11276_),
    .Z(_11284_));
 AND2_X1 _37445_ (.A1(_11284_),
    .A2(_11267_),
    .ZN(_11285_));
 NAND2_X1 _37446_ (.A1(_08491_),
    .A2(_11285_),
    .ZN(_11286_));
 MUX2_X1 _37447_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [454]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [972]),
    .S(_11248_),
    .Z(_11287_));
 AND2_X4 _37448_ (.A1(_11287_),
    .A2(_08501_),
    .ZN(_11288_));
 OAI21_X1 _37449_ (.A(_11288_),
    .B1(_11252_),
    .B2(_11254_),
    .ZN(_11289_));
 AOI21_X1 _37450_ (.A(_08494_),
    .B1(_11286_),
    .B2(_11289_),
    .ZN(_11290_));
 OR2_X1 _37451_ (.A1(_11283_),
    .A2(_11290_),
    .ZN(_11291_));
 MUX2_X2 _37452_ (.A(_11275_),
    .B(_11291_),
    .S(_08434_),
    .Z(\icache.data_mem_data_li [0]));
 MUX2_X1 _37453_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [263]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [781]),
    .S(_11248_),
    .Z(_11292_));
 BUF_X16 _37454_ (.A(_08426_),
    .Z(_11293_));
 BUF_X4 _37455_ (.A(_11293_),
    .Z(_11294_));
 AND2_X1 _37456_ (.A1(_11292_),
    .A2(_11294_),
    .ZN(_11295_));
 NAND2_X1 _37457_ (.A1(_08491_),
    .A2(_11295_),
    .ZN(_11296_));
 MUX2_X1 _37458_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [327]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [845]),
    .S(_11248_),
    .Z(_11297_));
 AND2_X1 _37459_ (.A1(_11297_),
    .A2(_11294_),
    .ZN(_11298_));
 OAI21_X1 _37460_ (.A(_11298_),
    .B1(_11252_),
    .B2(_11254_),
    .ZN(_11299_));
 AOI21_X1 _37461_ (.A(_11240_),
    .B1(_11296_),
    .B2(_11299_),
    .ZN(_11300_));
 BUF_X32 _37462_ (.A(_08489_),
    .Z(_11301_));
 BUF_X4 _37463_ (.A(_11301_),
    .Z(_11302_));
 MUX2_X2 _37464_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [391]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [909]),
    .S(_11264_),
    .Z(_11303_));
 AND2_X1 _37465_ (.A1(_11303_),
    .A2(_11267_),
    .ZN(_11304_));
 NAND2_X1 _37466_ (.A1(_11302_),
    .A2(_11304_),
    .ZN(_11305_));
 MUX2_X2 _37467_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [455]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [973]),
    .S(_11264_),
    .Z(_11306_));
 AND2_X1 _37468_ (.A1(_11306_),
    .A2(_11267_),
    .ZN(_11307_));
 OAI21_X1 _37469_ (.A(_11307_),
    .B1(_11270_),
    .B2(_11272_),
    .ZN(_11308_));
 AOI21_X1 _37470_ (.A(_11258_),
    .B1(_11305_),
    .B2(_11308_),
    .ZN(_11309_));
 OR2_X1 _37471_ (.A1(_11300_),
    .A2(_11309_),
    .ZN(_11310_));
 BUF_X16 _37472_ (.A(_08427_),
    .Z(_11311_));
 MUX2_X1 _37473_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [7]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [525]),
    .S(_11311_),
    .Z(_11312_));
 BUF_X16 _37474_ (.A(_11244_),
    .Z(_11313_));
 AND2_X4 _37475_ (.A1(_11312_),
    .A2(_11313_),
    .ZN(_11314_));
 NAND2_X1 _37476_ (.A1(_11302_),
    .A2(_11314_),
    .ZN(_11315_));
 MUX2_X2 _37477_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [71]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [589]),
    .S(_11264_),
    .Z(_11316_));
 AND2_X1 _37478_ (.A1(_11316_),
    .A2(_11267_),
    .ZN(_11317_));
 OAI21_X1 _37479_ (.A(_11317_),
    .B1(_11270_),
    .B2(_11272_),
    .ZN(_11318_));
 AOI21_X1 _37480_ (.A(_08448_),
    .B1(_11315_),
    .B2(_11318_),
    .ZN(_11319_));
 MUX2_X1 _37481_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [135]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [653]),
    .S(_11248_),
    .Z(_11320_));
 AND2_X1 _37482_ (.A1(_11320_),
    .A2(_11294_),
    .ZN(_11321_));
 NAND2_X1 _37483_ (.A1(_08491_),
    .A2(_11321_),
    .ZN(_11322_));
 MUX2_X1 _37484_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [199]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [717]),
    .S(_11248_),
    .Z(_11323_));
 AND2_X1 _37485_ (.A1(_11323_),
    .A2(_11294_),
    .ZN(_11324_));
 OAI21_X1 _37486_ (.A(_11324_),
    .B1(_11252_),
    .B2(_11254_),
    .ZN(_11325_));
 AOI21_X1 _37487_ (.A(_08494_),
    .B1(_11322_),
    .B2(_11325_),
    .ZN(_11326_));
 OR2_X1 _37488_ (.A1(_11319_),
    .A2(_11326_),
    .ZN(_11327_));
 MUX2_X2 _37489_ (.A(_11310_),
    .B(_11327_),
    .S(_08496_),
    .Z(\icache.data_mem_data_li [1]));
 BUF_X8 _37490_ (.A(_11239_),
    .Z(_11328_));
 MUX2_X2 _37491_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [264]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [782]),
    .S(_11264_),
    .Z(_11329_));
 BUF_X4 _37492_ (.A(_11266_),
    .Z(_11330_));
 AND2_X1 _37493_ (.A1(_11329_),
    .A2(_11330_),
    .ZN(_11331_));
 NAND2_X1 _37494_ (.A1(_11302_),
    .A2(_11331_),
    .ZN(_11332_));
 MUX2_X2 _37495_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [328]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [846]),
    .S(_11264_),
    .Z(_11333_));
 AND2_X1 _37496_ (.A1(_11333_),
    .A2(_11330_),
    .ZN(_11334_));
 BUF_X4 _37497_ (.A(_11269_),
    .Z(_11335_));
 BUF_X4 _37498_ (.A(_11271_),
    .Z(_11336_));
 OAI21_X1 _37499_ (.A(_11334_),
    .B1(_11335_),
    .B2(_11336_),
    .ZN(_11337_));
 AOI21_X1 _37500_ (.A(_11328_),
    .B1(_11332_),
    .B2(_11337_),
    .ZN(_11338_));
 MUX2_X2 _37501_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [392]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [910]),
    .S(_11264_),
    .Z(_11339_));
 AND2_X1 _37502_ (.A1(_11339_),
    .A2(_11330_),
    .ZN(_11340_));
 NAND2_X1 _37503_ (.A1(_11302_),
    .A2(_11340_),
    .ZN(_11341_));
 MUX2_X2 _37504_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [456]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [974]),
    .S(_11264_),
    .Z(_11342_));
 AND2_X1 _37505_ (.A1(_11342_),
    .A2(_11330_),
    .ZN(_11343_));
 OAI21_X1 _37506_ (.A(_11343_),
    .B1(_11335_),
    .B2(_11336_),
    .ZN(_11344_));
 AOI21_X1 _37507_ (.A(_11258_),
    .B1(_11341_),
    .B2(_11344_),
    .ZN(_11345_));
 OR2_X1 _37508_ (.A1(_11338_),
    .A2(_11345_),
    .ZN(_11346_));
 BUF_X16 _37509_ (.A(_11241_),
    .Z(_11347_));
 MUX2_X2 _37510_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [8]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [526]),
    .S(_11347_),
    .Z(_11348_));
 AND2_X4 _37511_ (.A1(_11348_),
    .A2(_11245_),
    .ZN(_11349_));
 NAND2_X1 _37512_ (.A1(_08491_),
    .A2(_11349_),
    .ZN(_11350_));
 MUX2_X2 _37513_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [72]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [590]),
    .S(_11248_),
    .Z(_11351_));
 AND2_X1 _37514_ (.A1(_11351_),
    .A2(_11294_),
    .ZN(_11352_));
 OAI21_X1 _37515_ (.A(_11352_),
    .B1(_11252_),
    .B2(_11254_),
    .ZN(_11353_));
 AOI21_X1 _37516_ (.A(_08448_),
    .B1(_11350_),
    .B2(_11353_),
    .ZN(_11354_));
 MUX2_X1 _37517_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [136]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [654]),
    .S(_11248_),
    .Z(_11355_));
 AND2_X1 _37518_ (.A1(_11355_),
    .A2(_11294_),
    .ZN(_11356_));
 NAND2_X1 _37519_ (.A1(_08491_),
    .A2(_11356_),
    .ZN(_11357_));
 BUF_X16 _37520_ (.A(_08428_),
    .Z(_11358_));
 MUX2_X1 _37521_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [200]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [718]),
    .S(_11358_),
    .Z(_11359_));
 AND2_X2 _37522_ (.A1(_11359_),
    .A2(_11294_),
    .ZN(_11360_));
 OAI21_X1 _37523_ (.A(_11360_),
    .B1(_11252_),
    .B2(_11254_),
    .ZN(_11361_));
 AOI21_X1 _37524_ (.A(_08494_),
    .B1(_11357_),
    .B2(_11361_),
    .ZN(_11362_));
 OR2_X1 _37525_ (.A1(_11354_),
    .A2(_11362_),
    .ZN(_11363_));
 MUX2_X2 _37526_ (.A(_11346_),
    .B(_11363_),
    .S(_08496_),
    .Z(\icache.data_mem_data_li [2]));
 MUX2_X1 _37527_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [265]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [783]),
    .S(_11264_),
    .Z(_11364_));
 AND2_X1 _37528_ (.A1(_11364_),
    .A2(_11330_),
    .ZN(_11365_));
 NAND2_X1 _37529_ (.A1(_11302_),
    .A2(_11365_),
    .ZN(_11366_));
 MUX2_X1 _37530_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [329]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [847]),
    .S(_11264_),
    .Z(_11367_));
 AND2_X1 _37531_ (.A1(_11367_),
    .A2(_11330_),
    .ZN(_11368_));
 OAI21_X1 _37532_ (.A(_11368_),
    .B1(_11335_),
    .B2(_11336_),
    .ZN(_11369_));
 AOI21_X1 _37533_ (.A(_11328_),
    .B1(_11366_),
    .B2(_11369_),
    .ZN(_11370_));
 BUF_X8 _37534_ (.A(_11257_),
    .Z(_11371_));
 BUF_X16 _37535_ (.A(_11263_),
    .Z(_11372_));
 MUX2_X2 _37536_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [393]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [911]),
    .S(_11372_),
    .Z(_11373_));
 AND2_X1 _37537_ (.A1(_11373_),
    .A2(_11330_),
    .ZN(_11374_));
 NAND2_X1 _37538_ (.A1(_11302_),
    .A2(_11374_),
    .ZN(_11375_));
 MUX2_X2 _37539_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [457]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [975]),
    .S(_11372_),
    .Z(_11376_));
 AND2_X1 _37540_ (.A1(_11376_),
    .A2(_11330_),
    .ZN(_11377_));
 OAI21_X1 _37541_ (.A(_11377_),
    .B1(_11335_),
    .B2(_11336_),
    .ZN(_11378_));
 AOI21_X1 _37542_ (.A(_11371_),
    .B1(_11375_),
    .B2(_11378_),
    .ZN(_11379_));
 OR2_X1 _37543_ (.A1(_11370_),
    .A2(_11379_),
    .ZN(_11380_));
 MUX2_X2 _37544_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [9]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [527]),
    .S(_11347_),
    .Z(_11381_));
 AND2_X4 _37545_ (.A1(_11381_),
    .A2(_11245_),
    .ZN(_11382_));
 NAND2_X1 _37546_ (.A1(_08491_),
    .A2(_11382_),
    .ZN(_11383_));
 MUX2_X1 _37547_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [73]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [591]),
    .S(_11358_),
    .Z(_11384_));
 AND2_X1 _37548_ (.A1(_11384_),
    .A2(_11294_),
    .ZN(_11385_));
 OAI21_X1 _37549_ (.A(_11385_),
    .B1(_11252_),
    .B2(_11254_),
    .ZN(_11386_));
 AOI21_X1 _37550_ (.A(_08448_),
    .B1(_11383_),
    .B2(_11386_),
    .ZN(_11387_));
 MUX2_X1 _37551_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [137]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [655]),
    .S(_11358_),
    .Z(_11388_));
 AND2_X2 _37552_ (.A1(_11388_),
    .A2(_11294_),
    .ZN(_11389_));
 NAND2_X1 _37553_ (.A1(_08491_),
    .A2(_11389_),
    .ZN(_11390_));
 MUX2_X2 _37554_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [201]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [719]),
    .S(_11358_),
    .Z(_11391_));
 AND2_X1 _37555_ (.A1(_11391_),
    .A2(_11294_),
    .ZN(_11392_));
 OAI21_X1 _37556_ (.A(_11392_),
    .B1(_11252_),
    .B2(_11254_),
    .ZN(_11393_));
 AOI21_X1 _37557_ (.A(_08494_),
    .B1(_11390_),
    .B2(_11393_),
    .ZN(_11394_));
 OR2_X1 _37558_ (.A1(_11387_),
    .A2(_11394_),
    .ZN(_11395_));
 MUX2_X2 _37559_ (.A(_11380_),
    .B(_11395_),
    .S(_08496_),
    .Z(\icache.data_mem_data_li [3]));
 MUX2_X1 _37560_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [266]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [784]),
    .S(_11372_),
    .Z(_11396_));
 AND2_X1 _37561_ (.A1(_11396_),
    .A2(_11330_),
    .ZN(_11397_));
 NAND2_X1 _37562_ (.A1(_11302_),
    .A2(_11397_),
    .ZN(_11398_));
 MUX2_X2 _37563_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [330]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [848]),
    .S(_11372_),
    .Z(_11399_));
 BUF_X4 _37564_ (.A(_11266_),
    .Z(_11400_));
 AND2_X1 _37565_ (.A1(_11399_),
    .A2(_11400_),
    .ZN(_11401_));
 OAI21_X1 _37566_ (.A(_11401_),
    .B1(_11335_),
    .B2(_11336_),
    .ZN(_11402_));
 AOI21_X1 _37567_ (.A(_11328_),
    .B1(_11398_),
    .B2(_11402_),
    .ZN(_11403_));
 MUX2_X1 _37568_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [394]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [912]),
    .S(_11358_),
    .Z(_11404_));
 BUF_X4 _37569_ (.A(_11293_),
    .Z(_11405_));
 AND2_X1 _37570_ (.A1(_11404_),
    .A2(_11405_),
    .ZN(_11406_));
 NAND2_X1 _37571_ (.A1(_11302_),
    .A2(_11406_),
    .ZN(_11407_));
 MUX2_X2 _37572_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [458]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [976]),
    .S(_11372_),
    .Z(_11408_));
 AND2_X2 _37573_ (.A1(_11408_),
    .A2(_11400_),
    .ZN(_11409_));
 OAI21_X1 _37574_ (.A(_11409_),
    .B1(_11335_),
    .B2(_11336_),
    .ZN(_11410_));
 AOI21_X1 _37575_ (.A(_11371_),
    .B1(_11407_),
    .B2(_11410_),
    .ZN(_11411_));
 OR2_X1 _37576_ (.A1(_11403_),
    .A2(_11411_),
    .ZN(_11412_));
 BUF_X16 _37577_ (.A(_08489_),
    .Z(_11413_));
 BUF_X4 _37578_ (.A(_11413_),
    .Z(_11414_));
 MUX2_X2 _37579_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [10]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [528]),
    .S(_11347_),
    .Z(_11415_));
 AND2_X4 _37580_ (.A1(_11415_),
    .A2(_11245_),
    .ZN(_11416_));
 NAND2_X1 _37581_ (.A1(_11414_),
    .A2(_11416_),
    .ZN(_11417_));
 MUX2_X1 _37582_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [74]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [592]),
    .S(_11358_),
    .Z(_11418_));
 AND2_X2 _37583_ (.A1(_11418_),
    .A2(_11405_),
    .ZN(_11419_));
 OAI21_X1 _37584_ (.A(_11419_),
    .B1(_11252_),
    .B2(_11254_),
    .ZN(_11420_));
 AOI21_X1 _37585_ (.A(_08448_),
    .B1(_11417_),
    .B2(_11420_),
    .ZN(_11421_));
 MUX2_X2 _37586_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [138]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [656]),
    .S(_11372_),
    .Z(_11422_));
 AND2_X1 _37587_ (.A1(_11422_),
    .A2(_11330_),
    .ZN(_11423_));
 NAND2_X1 _37588_ (.A1(_11414_),
    .A2(_11423_),
    .ZN(_11424_));
 MUX2_X2 _37589_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [202]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [720]),
    .S(_11358_),
    .Z(_11425_));
 AND2_X1 _37590_ (.A1(_11425_),
    .A2(_11405_),
    .ZN(_11426_));
 OAI21_X1 _37591_ (.A(_11426_),
    .B1(_11252_),
    .B2(_11254_),
    .ZN(_11427_));
 AOI21_X1 _37592_ (.A(_08494_),
    .B1(_11424_),
    .B2(_11427_),
    .ZN(_11428_));
 OR2_X1 _37593_ (.A1(_11421_),
    .A2(_11428_),
    .ZN(_11429_));
 MUX2_X2 _37594_ (.A(_11412_),
    .B(_11429_),
    .S(_08496_),
    .Z(\icache.data_mem_data_li [4]));
 MUX2_X2 _37595_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [267]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [785]),
    .S(_11358_),
    .Z(_11430_));
 AND2_X1 _37596_ (.A1(_11430_),
    .A2(_11405_),
    .ZN(_11431_));
 NAND2_X1 _37597_ (.A1(_11414_),
    .A2(_11431_),
    .ZN(_11432_));
 BUF_X16 _37598_ (.A(_08428_),
    .Z(_11433_));
 MUX2_X2 _37599_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [331]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [849]),
    .S(_11433_),
    .Z(_11434_));
 AND2_X1 _37600_ (.A1(_11434_),
    .A2(_11405_),
    .ZN(_11435_));
 BUF_X4 _37601_ (.A(_11251_),
    .Z(_11436_));
 BUF_X4 _37602_ (.A(_11253_),
    .Z(_11437_));
 OAI21_X1 _37603_ (.A(_11435_),
    .B1(_11436_),
    .B2(_11437_),
    .ZN(_11438_));
 AOI21_X1 _37604_ (.A(_11328_),
    .B1(_11432_),
    .B2(_11438_),
    .ZN(_11439_));
 MUX2_X2 _37605_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [395]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [913]),
    .S(_11372_),
    .Z(_11440_));
 AND2_X1 _37606_ (.A1(_11440_),
    .A2(_11400_),
    .ZN(_11441_));
 NAND2_X1 _37607_ (.A1(_11302_),
    .A2(_11441_),
    .ZN(_11442_));
 MUX2_X1 _37608_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [459]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [977]),
    .S(_11372_),
    .Z(_11443_));
 AND2_X1 _37609_ (.A1(_11443_),
    .A2(_11400_),
    .ZN(_11444_));
 OAI21_X1 _37610_ (.A(_11444_),
    .B1(_11335_),
    .B2(_11336_),
    .ZN(_11445_));
 AOI21_X1 _37611_ (.A(_11371_),
    .B1(_11442_),
    .B2(_11445_),
    .ZN(_11446_));
 OR2_X1 _37612_ (.A1(_11439_),
    .A2(_11446_),
    .ZN(_11447_));
 BUF_X16 _37613_ (.A(_08427_),
    .Z(_11448_));
 MUX2_X2 _37614_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [11]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [529]),
    .S(_11448_),
    .Z(_11449_));
 AND2_X4 _37615_ (.A1(_11449_),
    .A2(_11313_),
    .ZN(_11450_));
 NAND2_X1 _37616_ (.A1(_11302_),
    .A2(_11450_),
    .ZN(_11451_));
 MUX2_X2 _37617_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [75]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [593]),
    .S(_11372_),
    .Z(_11452_));
 AND2_X1 _37618_ (.A1(_11452_),
    .A2(_11400_),
    .ZN(_11453_));
 OAI21_X1 _37619_ (.A(_11453_),
    .B1(_11335_),
    .B2(_11336_),
    .ZN(_11454_));
 AOI21_X1 _37620_ (.A(_08448_),
    .B1(_11451_),
    .B2(_11454_),
    .ZN(_11455_));
 MUX2_X2 _37621_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [139]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [657]),
    .S(_11358_),
    .Z(_11456_));
 AND2_X1 _37622_ (.A1(_11456_),
    .A2(_11405_),
    .ZN(_11457_));
 NAND2_X1 _37623_ (.A1(_11414_),
    .A2(_11457_),
    .ZN(_11458_));
 MUX2_X2 _37624_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [203]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [721]),
    .S(_11358_),
    .Z(_11459_));
 AND2_X1 _37625_ (.A1(_11459_),
    .A2(_11405_),
    .ZN(_11460_));
 OAI21_X1 _37626_ (.A(_11460_),
    .B1(_11436_),
    .B2(_11437_),
    .ZN(_11461_));
 AOI21_X1 _37627_ (.A(_08494_),
    .B1(_11458_),
    .B2(_11461_),
    .ZN(_11462_));
 OR2_X1 _37628_ (.A1(_11455_),
    .A2(_11462_),
    .ZN(_11463_));
 MUX2_X2 _37629_ (.A(_11447_),
    .B(_11463_),
    .S(_08496_),
    .Z(\icache.data_mem_data_li [5]));
 MUX2_X2 _37630_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [268]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [786]),
    .S(_11433_),
    .Z(_11464_));
 AND2_X1 _37631_ (.A1(_11464_),
    .A2(_11405_),
    .ZN(_11465_));
 NAND2_X1 _37632_ (.A1(_11414_),
    .A2(_11465_),
    .ZN(_11466_));
 MUX2_X2 _37633_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [332]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [850]),
    .S(_11433_),
    .Z(_11467_));
 BUF_X4 _37634_ (.A(_11293_),
    .Z(_11468_));
 AND2_X1 _37635_ (.A1(_11467_),
    .A2(_11468_),
    .ZN(_11469_));
 OAI21_X1 _37636_ (.A(_11469_),
    .B1(_11436_),
    .B2(_11437_),
    .ZN(_11470_));
 AOI21_X1 _37637_ (.A(_11328_),
    .B1(_11466_),
    .B2(_11470_),
    .ZN(_11471_));
 BUF_X4 _37638_ (.A(_11301_),
    .Z(_11472_));
 BUF_X16 _37639_ (.A(_11263_),
    .Z(_11473_));
 MUX2_X2 _37640_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [396]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [914]),
    .S(_11473_),
    .Z(_11474_));
 AND2_X1 _37641_ (.A1(_11474_),
    .A2(_11400_),
    .ZN(_11475_));
 NAND2_X1 _37642_ (.A1(_11472_),
    .A2(_11475_),
    .ZN(_11476_));
 MUX2_X2 _37643_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [460]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [978]),
    .S(_11473_),
    .Z(_11477_));
 AND2_X1 _37644_ (.A1(_11477_),
    .A2(_11400_),
    .ZN(_11478_));
 OAI21_X1 _37645_ (.A(_11478_),
    .B1(_11335_),
    .B2(_11336_),
    .ZN(_11479_));
 AOI21_X1 _37646_ (.A(_11371_),
    .B1(_11476_),
    .B2(_11479_),
    .ZN(_11480_));
 OR2_X1 _37647_ (.A1(_11471_),
    .A2(_11480_),
    .ZN(_11481_));
 MUX2_X1 _37648_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [12]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [530]),
    .S(_11448_),
    .Z(_11482_));
 AND2_X4 _37649_ (.A1(_11482_),
    .A2(_11313_),
    .ZN(_11483_));
 NAND2_X1 _37650_ (.A1(_11472_),
    .A2(_11483_),
    .ZN(_11484_));
 MUX2_X2 _37651_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [76]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [594]),
    .S(_11372_),
    .Z(_11485_));
 AND2_X1 _37652_ (.A1(_11485_),
    .A2(_11400_),
    .ZN(_11486_));
 OAI21_X1 _37653_ (.A(_11486_),
    .B1(_11335_),
    .B2(_11336_),
    .ZN(_11487_));
 AOI21_X1 _37654_ (.A(_08448_),
    .B1(_11484_),
    .B2(_11487_),
    .ZN(_11488_));
 MUX2_X1 _37655_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [140]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [658]),
    .S(_11433_),
    .Z(_11489_));
 AND2_X1 _37656_ (.A1(_11489_),
    .A2(_11405_),
    .ZN(_11490_));
 NAND2_X1 _37657_ (.A1(_11414_),
    .A2(_11490_),
    .ZN(_11491_));
 MUX2_X1 _37658_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [204]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [722]),
    .S(_11433_),
    .Z(_11492_));
 AND2_X1 _37659_ (.A1(_11492_),
    .A2(_11405_),
    .ZN(_11493_));
 OAI21_X1 _37660_ (.A(_11493_),
    .B1(_11436_),
    .B2(_11437_),
    .ZN(_11494_));
 AOI21_X1 _37661_ (.A(_08494_),
    .B1(_11491_),
    .B2(_11494_),
    .ZN(_11495_));
 OR2_X1 _37662_ (.A1(_11488_),
    .A2(_11495_),
    .ZN(_11496_));
 MUX2_X2 _37663_ (.A(_11481_),
    .B(_11496_),
    .S(_08496_),
    .Z(\icache.data_mem_data_li [6]));
 MUX2_X2 _37664_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [13]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [531]),
    .S(_11347_),
    .Z(_11497_));
 AND2_X4 _37665_ (.A1(_11497_),
    .A2(_11245_),
    .ZN(_11498_));
 NAND2_X1 _37666_ (.A1(_11414_),
    .A2(_11498_),
    .ZN(_11499_));
 MUX2_X1 _37667_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [77]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [595]),
    .S(_11433_),
    .Z(_11500_));
 AND2_X1 _37668_ (.A1(_11500_),
    .A2(_11468_),
    .ZN(_11501_));
 OAI21_X1 _37669_ (.A(_11501_),
    .B1(_11436_),
    .B2(_11437_),
    .ZN(_11502_));
 AOI21_X1 _37670_ (.A(_11328_),
    .B1(_11499_),
    .B2(_11502_),
    .ZN(_11503_));
 MUX2_X1 _37671_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [141]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [659]),
    .S(_11433_),
    .Z(_11504_));
 AND2_X1 _37672_ (.A1(_11504_),
    .A2(_11468_),
    .ZN(_11505_));
 NAND2_X1 _37673_ (.A1(_11472_),
    .A2(_11505_),
    .ZN(_11506_));
 MUX2_X2 _37674_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [205]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [723]),
    .S(_11473_),
    .Z(_11507_));
 BUF_X4 _37675_ (.A(_11266_),
    .Z(_11508_));
 AND2_X1 _37676_ (.A1(_11507_),
    .A2(_11508_),
    .ZN(_11509_));
 BUF_X4 _37677_ (.A(_11269_),
    .Z(_11510_));
 BUF_X4 _37678_ (.A(_11271_),
    .Z(_11511_));
 OAI21_X1 _37679_ (.A(_11509_),
    .B1(_11510_),
    .B2(_11511_),
    .ZN(_11512_));
 AOI21_X1 _37680_ (.A(_11371_),
    .B1(_11506_),
    .B2(_11512_),
    .ZN(_11513_));
 OR2_X1 _37681_ (.A1(_11503_),
    .A2(_11513_),
    .ZN(_11514_));
 MUX2_X2 _37682_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [269]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [787]),
    .S(_11473_),
    .Z(_11515_));
 AND2_X1 _37683_ (.A1(_11515_),
    .A2(_11400_),
    .ZN(_11516_));
 NAND2_X1 _37684_ (.A1(_11472_),
    .A2(_11516_),
    .ZN(_11517_));
 MUX2_X1 _37685_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [333]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [851]),
    .S(_11473_),
    .Z(_11518_));
 AND2_X1 _37686_ (.A1(_11518_),
    .A2(_11400_),
    .ZN(_11519_));
 OAI21_X1 _37687_ (.A(_11519_),
    .B1(_11510_),
    .B2(_11511_),
    .ZN(_11520_));
 AOI21_X1 _37688_ (.A(_08448_),
    .B1(_11517_),
    .B2(_11520_),
    .ZN(_11521_));
 MUX2_X2 _37689_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [397]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [915]),
    .S(_11473_),
    .Z(_11522_));
 AND2_X1 _37690_ (.A1(_11522_),
    .A2(_11508_),
    .ZN(_11523_));
 NAND2_X1 _37691_ (.A1(_11414_),
    .A2(_11523_),
    .ZN(_11524_));
 MUX2_X2 _37692_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [461]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [979]),
    .S(_11433_),
    .Z(_11525_));
 AND2_X1 _37693_ (.A1(_11525_),
    .A2(_11468_),
    .ZN(_11526_));
 OAI21_X1 _37694_ (.A(_11526_),
    .B1(_11436_),
    .B2(_11437_),
    .ZN(_11527_));
 AOI21_X1 _37695_ (.A(_08494_),
    .B1(_11524_),
    .B2(_11527_),
    .ZN(_11528_));
 OR2_X1 _37696_ (.A1(_11521_),
    .A2(_11528_),
    .ZN(_11529_));
 MUX2_X2 _37697_ (.A(_11514_),
    .B(_11529_),
    .S(_08434_),
    .Z(\icache.data_mem_data_li [7]));
 MUX2_X1 _37698_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [270]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [788]),
    .S(_11433_),
    .Z(_11530_));
 AND2_X2 _37699_ (.A1(_11530_),
    .A2(_11468_),
    .ZN(_11531_));
 NAND2_X1 _37700_ (.A1(_11414_),
    .A2(_11531_),
    .ZN(_11532_));
 BUF_X8 _37701_ (.A(_08428_),
    .Z(_11533_));
 MUX2_X2 _37702_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [334]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [852]),
    .S(_11533_),
    .Z(_11534_));
 AND2_X1 _37703_ (.A1(_11534_),
    .A2(_11468_),
    .ZN(_11535_));
 OAI21_X1 _37704_ (.A(_11535_),
    .B1(_11436_),
    .B2(_11437_),
    .ZN(_11536_));
 AOI21_X1 _37705_ (.A(_11328_),
    .B1(_11532_),
    .B2(_11536_),
    .ZN(_11537_));
 MUX2_X2 _37706_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [398]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [916]),
    .S(_11533_),
    .Z(_11538_));
 AND2_X1 _37707_ (.A1(_11538_),
    .A2(_11468_),
    .ZN(_11539_));
 NAND2_X1 _37708_ (.A1(_11472_),
    .A2(_11539_),
    .ZN(_11540_));
 MUX2_X1 _37709_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [462]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [980]),
    .S(_11473_),
    .Z(_11541_));
 AND2_X1 _37710_ (.A1(_11541_),
    .A2(_11508_),
    .ZN(_11542_));
 OAI21_X1 _37711_ (.A(_11542_),
    .B1(_11510_),
    .B2(_11511_),
    .ZN(_11543_));
 AOI21_X1 _37712_ (.A(_11371_),
    .B1(_11540_),
    .B2(_11543_),
    .ZN(_11544_));
 OR2_X1 _37713_ (.A1(_11537_),
    .A2(_11544_),
    .ZN(_11545_));
 BUF_X16 _37714_ (.A(_08447_),
    .Z(_11546_));
 BUF_X8 _37715_ (.A(_11546_),
    .Z(_11547_));
 MUX2_X2 _37716_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [14]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [532]),
    .S(_11448_),
    .Z(_11548_));
 AND2_X4 _37717_ (.A1(_11548_),
    .A2(_11313_),
    .ZN(_11549_));
 NAND2_X1 _37718_ (.A1(_11472_),
    .A2(_11549_),
    .ZN(_11550_));
 MUX2_X2 _37719_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [78]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [596]),
    .S(_11473_),
    .Z(_11551_));
 AND2_X1 _37720_ (.A1(_11551_),
    .A2(_11508_),
    .ZN(_11552_));
 OAI21_X1 _37721_ (.A(_11552_),
    .B1(_11510_),
    .B2(_11511_),
    .ZN(_11553_));
 AOI21_X1 _37722_ (.A(_11547_),
    .B1(_11550_),
    .B2(_11553_),
    .ZN(_11554_));
 MUX2_X1 _37723_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [142]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [660]),
    .S(_11473_),
    .Z(_11555_));
 AND2_X1 _37724_ (.A1(_11555_),
    .A2(_11508_),
    .ZN(_11556_));
 NAND2_X1 _37725_ (.A1(_11414_),
    .A2(_11556_),
    .ZN(_11557_));
 MUX2_X2 _37726_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [206]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [724]),
    .S(_11433_),
    .Z(_11558_));
 AND2_X1 _37727_ (.A1(_11558_),
    .A2(_11468_),
    .ZN(_11559_));
 OAI21_X1 _37728_ (.A(_11559_),
    .B1(_11436_),
    .B2(_11437_),
    .ZN(_11560_));
 AOI21_X1 _37729_ (.A(_08494_),
    .B1(_11557_),
    .B2(_11560_),
    .ZN(_11561_));
 OR2_X1 _37730_ (.A1(_11554_),
    .A2(_11561_),
    .ZN(_11562_));
 MUX2_X2 _37731_ (.A(_11545_),
    .B(_11562_),
    .S(_08496_),
    .Z(\icache.data_mem_data_li [8]));
 BUF_X4 _37732_ (.A(_11413_),
    .Z(_11563_));
 MUX2_X2 _37733_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [15]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [533]),
    .S(_11347_),
    .Z(_11564_));
 BUF_X16 _37734_ (.A(_11244_),
    .Z(_11565_));
 AND2_X4 _37735_ (.A1(_11564_),
    .A2(_11565_),
    .ZN(_11566_));
 NAND2_X1 _37736_ (.A1(_11563_),
    .A2(_11566_),
    .ZN(_11567_));
 MUX2_X1 _37737_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [79]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [597]),
    .S(_11533_),
    .Z(_11568_));
 AND2_X1 _37738_ (.A1(_11568_),
    .A2(_11468_),
    .ZN(_11569_));
 OAI21_X1 _37739_ (.A(_11569_),
    .B1(_11436_),
    .B2(_11437_),
    .ZN(_11570_));
 AOI21_X1 _37740_ (.A(_11328_),
    .B1(_11567_),
    .B2(_11570_),
    .ZN(_11571_));
 MUX2_X1 _37741_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [143]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [661]),
    .S(_11533_),
    .Z(_11572_));
 BUF_X4 _37742_ (.A(_11293_),
    .Z(_11573_));
 AND2_X2 _37743_ (.A1(_11572_),
    .A2(_11573_),
    .ZN(_11574_));
 NAND2_X1 _37744_ (.A1(_11472_),
    .A2(_11574_),
    .ZN(_11575_));
 BUF_X8 _37745_ (.A(_11263_),
    .Z(_11576_));
 MUX2_X1 _37746_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [207]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [725]),
    .S(_11576_),
    .Z(_11577_));
 AND2_X1 _37747_ (.A1(_11577_),
    .A2(_11508_),
    .ZN(_11578_));
 OAI21_X1 _37748_ (.A(_11578_),
    .B1(_11510_),
    .B2(_11511_),
    .ZN(_11579_));
 AOI21_X1 _37749_ (.A(_11371_),
    .B1(_11575_),
    .B2(_11579_),
    .ZN(_11580_));
 OR2_X2 _37750_ (.A1(_11571_),
    .A2(_11580_),
    .ZN(_11581_));
 MUX2_X2 _37751_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [271]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [789]),
    .S(_11473_),
    .Z(_11582_));
 AND2_X1 _37752_ (.A1(_11582_),
    .A2(_11508_),
    .ZN(_11583_));
 NAND2_X1 _37753_ (.A1(_11472_),
    .A2(_11583_),
    .ZN(_11584_));
 MUX2_X1 _37754_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [335]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [853]),
    .S(_11576_),
    .Z(_11585_));
 AND2_X1 _37755_ (.A1(_11585_),
    .A2(_11508_),
    .ZN(_11586_));
 OAI21_X1 _37756_ (.A(_11586_),
    .B1(_11510_),
    .B2(_11511_),
    .ZN(_11587_));
 AOI21_X1 _37757_ (.A(_11547_),
    .B1(_11584_),
    .B2(_11587_),
    .ZN(_11588_));
 BUF_X8 _37758_ (.A(_08493_),
    .Z(_11589_));
 MUX2_X2 _37759_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [399]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [917]),
    .S(_11576_),
    .Z(_11590_));
 AND2_X1 _37760_ (.A1(_11590_),
    .A2(_11508_),
    .ZN(_11591_));
 NAND2_X1 _37761_ (.A1(_11563_),
    .A2(_11591_),
    .ZN(_11592_));
 MUX2_X1 _37762_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [463]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [981]),
    .S(_11533_),
    .Z(_11593_));
 AND2_X2 _37763_ (.A1(_11593_),
    .A2(_11468_),
    .ZN(_11594_));
 OAI21_X2 _37764_ (.A(_11594_),
    .B1(_11436_),
    .B2(_11437_),
    .ZN(_11595_));
 AOI21_X1 _37765_ (.A(_11589_),
    .B1(_11592_),
    .B2(_11595_),
    .ZN(_11596_));
 OR2_X2 _37766_ (.A1(_11588_),
    .A2(_11596_),
    .ZN(_11597_));
 MUX2_X2 _37767_ (.A(_11581_),
    .B(_11597_),
    .S(_08434_),
    .Z(\icache.data_mem_data_li [9]));
 MUX2_X2 _37768_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [16]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [534]),
    .S(_11347_),
    .Z(_11598_));
 AND2_X4 _37769_ (.A1(_11598_),
    .A2(_11565_),
    .ZN(_11599_));
 NAND2_X1 _37770_ (.A1(_11472_),
    .A2(_11599_),
    .ZN(_11600_));
 MUX2_X1 _37771_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [80]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [598]),
    .S(_11576_),
    .Z(_11601_));
 BUF_X4 _37772_ (.A(_11266_),
    .Z(_11602_));
 AND2_X1 _37773_ (.A1(_11601_),
    .A2(_11602_),
    .ZN(_11603_));
 OAI21_X1 _37774_ (.A(_11603_),
    .B1(_11510_),
    .B2(_11511_),
    .ZN(_11604_));
 AOI21_X1 _37775_ (.A(_11328_),
    .B1(_11600_),
    .B2(_11604_),
    .ZN(_11605_));
 MUX2_X2 _37776_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [144]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [662]),
    .S(_11533_),
    .Z(_11606_));
 AND2_X2 _37777_ (.A1(_11606_),
    .A2(_11573_),
    .ZN(_11607_));
 NAND2_X1 _37778_ (.A1(_11472_),
    .A2(_11607_),
    .ZN(_11608_));
 MUX2_X1 _37779_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [208]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [726]),
    .S(_11576_),
    .Z(_11609_));
 AND2_X1 _37780_ (.A1(_11609_),
    .A2(_11602_),
    .ZN(_11610_));
 OAI21_X1 _37781_ (.A(_11610_),
    .B1(_11510_),
    .B2(_11511_),
    .ZN(_11611_));
 AOI21_X1 _37782_ (.A(_11371_),
    .B1(_11608_),
    .B2(_11611_),
    .ZN(_11612_));
 OR2_X1 _37783_ (.A1(_11605_),
    .A2(_11612_),
    .ZN(_11613_));
 MUX2_X1 _37784_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [272]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [790]),
    .S(_11576_),
    .Z(_11614_));
 AND2_X1 _37785_ (.A1(_11614_),
    .A2(_11508_),
    .ZN(_11615_));
 NAND2_X1 _37786_ (.A1(_11563_),
    .A2(_11615_),
    .ZN(_11616_));
 MUX2_X2 _37787_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [336]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [854]),
    .S(_11533_),
    .Z(_11617_));
 AND2_X1 _37788_ (.A1(_11617_),
    .A2(_11573_),
    .ZN(_11618_));
 BUF_X4 _37789_ (.A(_11251_),
    .Z(_11619_));
 BUF_X4 _37790_ (.A(_11253_),
    .Z(_11620_));
 OAI21_X1 _37791_ (.A(_11618_),
    .B1(_11619_),
    .B2(_11620_),
    .ZN(_11621_));
 AOI21_X1 _37792_ (.A(_11547_),
    .B1(_11616_),
    .B2(_11621_),
    .ZN(_11622_));
 MUX2_X1 _37793_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [400]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [918]),
    .S(_11576_),
    .Z(_11623_));
 AND2_X2 _37794_ (.A1(_11623_),
    .A2(_11602_),
    .ZN(_11624_));
 NAND2_X1 _37795_ (.A1(_11563_),
    .A2(_11624_),
    .ZN(_11625_));
 MUX2_X2 _37796_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [464]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [982]),
    .S(_11533_),
    .Z(_11626_));
 AND2_X1 _37797_ (.A1(_11626_),
    .A2(_11573_),
    .ZN(_11627_));
 OAI21_X1 _37798_ (.A(_11627_),
    .B1(_11619_),
    .B2(_11620_),
    .ZN(_11628_));
 AOI21_X1 _37799_ (.A(_11589_),
    .B1(_11625_),
    .B2(_11628_),
    .ZN(_11629_));
 OR2_X1 _37800_ (.A1(_11622_),
    .A2(_11629_),
    .ZN(_11630_));
 MUX2_X2 _37801_ (.A(_11613_),
    .B(_11630_),
    .S(_08434_),
    .Z(\icache.data_mem_data_li [10]));
 MUX2_X1 _37802_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [17]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [535]),
    .S(_11347_),
    .Z(_11631_));
 AND2_X4 _37803_ (.A1(_11631_),
    .A2(_11565_),
    .ZN(_11632_));
 NAND2_X1 _37804_ (.A1(_11563_),
    .A2(_11632_),
    .ZN(_11633_));
 MUX2_X1 _37805_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [81]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [599]),
    .S(_11533_),
    .Z(_11634_));
 AND2_X1 _37806_ (.A1(_11634_),
    .A2(_11573_),
    .ZN(_11635_));
 OAI21_X1 _37807_ (.A(_11635_),
    .B1(_11619_),
    .B2(_11620_),
    .ZN(_11636_));
 AOI21_X1 _37808_ (.A(_11328_),
    .B1(_11633_),
    .B2(_11636_),
    .ZN(_11637_));
 BUF_X4 _37809_ (.A(_11301_),
    .Z(_11638_));
 BUF_X8 _37810_ (.A(_08428_),
    .Z(_11639_));
 MUX2_X1 _37811_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [145]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [663]),
    .S(_11639_),
    .Z(_11640_));
 AND2_X1 _37812_ (.A1(_11640_),
    .A2(_11573_),
    .ZN(_11641_));
 NAND2_X1 _37813_ (.A1(_11638_),
    .A2(_11641_),
    .ZN(_11642_));
 BUF_X16 _37814_ (.A(_08427_),
    .Z(_11643_));
 BUF_X8 _37815_ (.A(_11643_),
    .Z(_11644_));
 MUX2_X1 _37816_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [209]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [727]),
    .S(_11644_),
    .Z(_11645_));
 AND2_X2 _37817_ (.A1(_11645_),
    .A2(_11602_),
    .ZN(_11646_));
 OAI21_X1 _37818_ (.A(_11646_),
    .B1(_11510_),
    .B2(_11511_),
    .ZN(_11647_));
 AOI21_X1 _37819_ (.A(_11371_),
    .B1(_11642_),
    .B2(_11647_),
    .ZN(_11648_));
 OR2_X1 _37820_ (.A1(_11637_),
    .A2(_11648_),
    .ZN(_11649_));
 MUX2_X1 _37821_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [273]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [791]),
    .S(_11576_),
    .Z(_11650_));
 AND2_X1 _37822_ (.A1(_11650_),
    .A2(_11602_),
    .ZN(_11651_));
 NAND2_X1 _37823_ (.A1(_11638_),
    .A2(_11651_),
    .ZN(_11652_));
 MUX2_X2 _37824_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [337]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [855]),
    .S(_11576_),
    .Z(_11653_));
 AND2_X1 _37825_ (.A1(_11653_),
    .A2(_11602_),
    .ZN(_11654_));
 OAI21_X1 _37826_ (.A(_11654_),
    .B1(_11510_),
    .B2(_11511_),
    .ZN(_11655_));
 AOI21_X1 _37827_ (.A(_11547_),
    .B1(_11652_),
    .B2(_11655_),
    .ZN(_11656_));
 MUX2_X1 _37828_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [401]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [919]),
    .S(_11576_),
    .Z(_11657_));
 AND2_X1 _37829_ (.A1(_11657_),
    .A2(_11602_),
    .ZN(_11658_));
 NAND2_X1 _37830_ (.A1(_11563_),
    .A2(_11658_),
    .ZN(_11659_));
 MUX2_X1 _37831_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [465]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [983]),
    .S(_11533_),
    .Z(_11660_));
 AND2_X1 _37832_ (.A1(_11660_),
    .A2(_11573_),
    .ZN(_11661_));
 OAI21_X1 _37833_ (.A(_11661_),
    .B1(_11619_),
    .B2(_11620_),
    .ZN(_11662_));
 AOI21_X1 _37834_ (.A(_11589_),
    .B1(_11659_),
    .B2(_11662_),
    .ZN(_11663_));
 OR2_X1 _37835_ (.A1(_11656_),
    .A2(_11663_),
    .ZN(_11664_));
 MUX2_X2 _37836_ (.A(_11649_),
    .B(_11664_),
    .S(_08434_),
    .Z(\icache.data_mem_data_li [11]));
 BUF_X32 _37837_ (.A(_08447_),
    .Z(_11665_));
 BUF_X8 _37838_ (.A(_11665_),
    .Z(_11666_));
 MUX2_X1 _37839_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [274]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [792]),
    .S(_11639_),
    .Z(_11667_));
 AND2_X1 _37840_ (.A1(_11667_),
    .A2(_11573_),
    .ZN(_11668_));
 NAND2_X1 _37841_ (.A1(_11563_),
    .A2(_11668_),
    .ZN(_11669_));
 MUX2_X1 _37842_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [338]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [856]),
    .S(_11639_),
    .Z(_11670_));
 BUF_X4 _37843_ (.A(_11293_),
    .Z(_11671_));
 AND2_X2 _37844_ (.A1(_11670_),
    .A2(_11671_),
    .ZN(_11672_));
 OAI21_X1 _37845_ (.A(_11672_),
    .B1(_11619_),
    .B2(_11620_),
    .ZN(_11673_));
 AOI21_X1 _37846_ (.A(_11666_),
    .B1(_11669_),
    .B2(_11673_),
    .ZN(_11674_));
 MUX2_X2 _37847_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [402]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [920]),
    .S(_11644_),
    .Z(_11675_));
 AND2_X1 _37848_ (.A1(_11675_),
    .A2(_11602_),
    .ZN(_11676_));
 NAND2_X1 _37849_ (.A1(_11638_),
    .A2(_11676_),
    .ZN(_11677_));
 MUX2_X1 _37850_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [466]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [984]),
    .S(_11644_),
    .Z(_11678_));
 AND2_X1 _37851_ (.A1(_11678_),
    .A2(_11602_),
    .ZN(_11679_));
 BUF_X16 _37852_ (.A(_08483_),
    .Z(_11680_));
 BUF_X4 _37853_ (.A(_11680_),
    .Z(_11681_));
 BUF_X16 _37854_ (.A(_08487_),
    .Z(_11682_));
 BUF_X4 _37855_ (.A(_11682_),
    .Z(_11683_));
 OAI21_X1 _37856_ (.A(_11679_),
    .B1(_11681_),
    .B2(_11683_),
    .ZN(_11684_));
 AOI21_X1 _37857_ (.A(_11371_),
    .B1(_11677_),
    .B2(_11684_),
    .ZN(_11685_));
 OR2_X1 _37858_ (.A1(_11674_),
    .A2(_11685_),
    .ZN(_11686_));
 MUX2_X2 _37859_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [18]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [536]),
    .S(_11448_),
    .Z(_11687_));
 AND2_X4 _37860_ (.A1(_11687_),
    .A2(_11313_),
    .ZN(_11688_));
 NAND2_X1 _37861_ (.A1(_11638_),
    .A2(_11688_),
    .ZN(_11689_));
 MUX2_X2 _37862_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [82]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [600]),
    .S(_11644_),
    .Z(_11690_));
 AND2_X1 _37863_ (.A1(_11690_),
    .A2(_11602_),
    .ZN(_11691_));
 OAI21_X2 _37864_ (.A(_11691_),
    .B1(_11681_),
    .B2(_11683_),
    .ZN(_11692_));
 AOI21_X1 _37865_ (.A(_11547_),
    .B1(_11689_),
    .B2(_11692_),
    .ZN(_11693_));
 MUX2_X2 _37866_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [146]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [664]),
    .S(_11639_),
    .Z(_11694_));
 AND2_X1 _37867_ (.A1(_11694_),
    .A2(_11573_),
    .ZN(_11695_));
 NAND2_X1 _37868_ (.A1(_11563_),
    .A2(_11695_),
    .ZN(_11696_));
 MUX2_X1 _37869_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [210]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [728]),
    .S(_11639_),
    .Z(_11697_));
 AND2_X1 _37870_ (.A1(_11697_),
    .A2(_11573_),
    .ZN(_11698_));
 OAI21_X1 _37871_ (.A(_11698_),
    .B1(_11619_),
    .B2(_11620_),
    .ZN(_11699_));
 AOI21_X1 _37872_ (.A(_11589_),
    .B1(_11696_),
    .B2(_11699_),
    .ZN(_11700_));
 OR2_X1 _37873_ (.A1(_11693_),
    .A2(_11700_),
    .ZN(_11701_));
 MUX2_X2 _37874_ (.A(_11686_),
    .B(_11701_),
    .S(_08496_),
    .Z(\icache.data_mem_data_li [12]));
 MUX2_X1 _37875_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [275]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [793]),
    .S(_11639_),
    .Z(_11702_));
 AND2_X1 _37876_ (.A1(_11702_),
    .A2(_11671_),
    .ZN(_11703_));
 NAND2_X1 _37877_ (.A1(_11563_),
    .A2(_11703_),
    .ZN(_11704_));
 MUX2_X1 _37878_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [339]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [857]),
    .S(_11639_),
    .Z(_11705_));
 AND2_X2 _37879_ (.A1(_11705_),
    .A2(_11671_),
    .ZN(_11706_));
 OAI21_X1 _37880_ (.A(_11706_),
    .B1(_11619_),
    .B2(_11620_),
    .ZN(_11707_));
 AOI21_X1 _37881_ (.A(_11666_),
    .B1(_11704_),
    .B2(_11707_),
    .ZN(_11708_));
 BUF_X16 _37882_ (.A(_08446_),
    .Z(_11709_));
 BUF_X8 _37883_ (.A(_11709_),
    .Z(_11710_));
 MUX2_X2 _37884_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [403]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [921]),
    .S(_11644_),
    .Z(_11711_));
 BUF_X4 _37885_ (.A(_11266_),
    .Z(_11712_));
 AND2_X1 _37886_ (.A1(_11711_),
    .A2(_11712_),
    .ZN(_11713_));
 NAND2_X1 _37887_ (.A1(_11638_),
    .A2(_11713_),
    .ZN(_11714_));
 MUX2_X1 _37888_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [467]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [985]),
    .S(_11644_),
    .Z(_11715_));
 AND2_X1 _37889_ (.A1(_11715_),
    .A2(_11712_),
    .ZN(_11716_));
 OAI21_X2 _37890_ (.A(_11716_),
    .B1(_11681_),
    .B2(_11683_),
    .ZN(_11717_));
 AOI21_X1 _37891_ (.A(_11710_),
    .B1(_11714_),
    .B2(_11717_),
    .ZN(_11718_));
 OR2_X1 _37892_ (.A1(_11708_),
    .A2(_11718_),
    .ZN(_11719_));
 MUX2_X1 _37893_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [19]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [537]),
    .S(_11448_),
    .Z(_11720_));
 BUF_X16 _37894_ (.A(_11244_),
    .Z(_11721_));
 AND2_X4 _37895_ (.A1(_11720_),
    .A2(_11721_),
    .ZN(_11722_));
 NAND2_X1 _37896_ (.A1(_11638_),
    .A2(_11722_),
    .ZN(_11723_));
 MUX2_X2 _37897_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [83]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [601]),
    .S(_11644_),
    .Z(_11724_));
 AND2_X1 _37898_ (.A1(_11724_),
    .A2(_11712_),
    .ZN(_11725_));
 OAI21_X1 _37899_ (.A(_11725_),
    .B1(_11681_),
    .B2(_11683_),
    .ZN(_11726_));
 AOI21_X1 _37900_ (.A(_11547_),
    .B1(_11723_),
    .B2(_11726_),
    .ZN(_11727_));
 MUX2_X1 _37901_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [147]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [665]),
    .S(_11639_),
    .Z(_11728_));
 AND2_X1 _37902_ (.A1(_11728_),
    .A2(_11671_),
    .ZN(_11729_));
 NAND2_X1 _37903_ (.A1(_11563_),
    .A2(_11729_),
    .ZN(_11730_));
 MUX2_X1 _37904_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [211]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [729]),
    .S(_11639_),
    .Z(_11731_));
 AND2_X1 _37905_ (.A1(_11731_),
    .A2(_11671_),
    .ZN(_11732_));
 OAI21_X1 _37906_ (.A(_11732_),
    .B1(_11619_),
    .B2(_11620_),
    .ZN(_11733_));
 AOI21_X1 _37907_ (.A(_11589_),
    .B1(_11730_),
    .B2(_11733_),
    .ZN(_11734_));
 OR2_X1 _37908_ (.A1(_11727_),
    .A2(_11734_),
    .ZN(_11735_));
 MUX2_X2 _37909_ (.A(_11719_),
    .B(_11735_),
    .S(_08496_),
    .Z(\icache.data_mem_data_li [13]));
 MUX2_X1 _37910_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [276]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [794]),
    .S(_11644_),
    .Z(_11736_));
 AND2_X1 _37911_ (.A1(_11736_),
    .A2(_11712_),
    .ZN(_11737_));
 NAND2_X1 _37912_ (.A1(_11638_),
    .A2(_11737_),
    .ZN(_11738_));
 MUX2_X1 _37913_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [340]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [858]),
    .S(_11644_),
    .Z(_11739_));
 AND2_X1 _37914_ (.A1(_11739_),
    .A2(_11712_),
    .ZN(_11740_));
 OAI21_X1 _37915_ (.A(_11740_),
    .B1(_11681_),
    .B2(_11683_),
    .ZN(_11741_));
 AOI21_X1 _37916_ (.A(_11666_),
    .B1(_11738_),
    .B2(_11741_),
    .ZN(_11742_));
 BUF_X8 _37917_ (.A(_08428_),
    .Z(_11743_));
 MUX2_X2 _37918_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [404]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [922]),
    .S(_11743_),
    .Z(_11744_));
 AND2_X2 _37919_ (.A1(_11744_),
    .A2(_11671_),
    .ZN(_11745_));
 NAND2_X1 _37920_ (.A1(_11638_),
    .A2(_11745_),
    .ZN(_11746_));
 BUF_X8 _37921_ (.A(_11643_),
    .Z(_11747_));
 MUX2_X2 _37922_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [468]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [986]),
    .S(_11747_),
    .Z(_11748_));
 AND2_X2 _37923_ (.A1(_11748_),
    .A2(_11712_),
    .ZN(_11749_));
 OAI21_X1 _37924_ (.A(_11749_),
    .B1(_11681_),
    .B2(_11683_),
    .ZN(_11750_));
 AOI21_X1 _37925_ (.A(_11710_),
    .B1(_11746_),
    .B2(_11750_),
    .ZN(_11751_));
 OR2_X1 _37926_ (.A1(_11742_),
    .A2(_11751_),
    .ZN(_11752_));
 BUF_X8 _37927_ (.A(_11413_),
    .Z(_11753_));
 MUX2_X1 _37928_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [20]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [538]),
    .S(_11347_),
    .Z(_11754_));
 AND2_X4 _37929_ (.A1(_11754_),
    .A2(_11565_),
    .ZN(_11755_));
 NAND2_X1 _37930_ (.A1(_11753_),
    .A2(_11755_),
    .ZN(_11756_));
 MUX2_X1 _37931_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [84]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [602]),
    .S(_11639_),
    .Z(_11757_));
 AND2_X2 _37932_ (.A1(_11757_),
    .A2(_11671_),
    .ZN(_11758_));
 OAI21_X1 _37933_ (.A(_11758_),
    .B1(_11619_),
    .B2(_11620_),
    .ZN(_11759_));
 AOI21_X1 _37934_ (.A(_11547_),
    .B1(_11756_),
    .B2(_11759_),
    .ZN(_11760_));
 MUX2_X1 _37935_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [148]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [666]),
    .S(_11644_),
    .Z(_11761_));
 AND2_X1 _37936_ (.A1(_11761_),
    .A2(_11712_),
    .ZN(_11762_));
 NAND2_X1 _37937_ (.A1(_11753_),
    .A2(_11762_),
    .ZN(_11763_));
 MUX2_X1 _37938_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [212]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [730]),
    .S(_11743_),
    .Z(_11764_));
 AND2_X1 _37939_ (.A1(_11764_),
    .A2(_11671_),
    .ZN(_11765_));
 OAI21_X1 _37940_ (.A(_11765_),
    .B1(_11619_),
    .B2(_11620_),
    .ZN(_11766_));
 AOI21_X1 _37941_ (.A(_11589_),
    .B1(_11763_),
    .B2(_11766_),
    .ZN(_11767_));
 OR2_X1 _37942_ (.A1(_11760_),
    .A2(_11767_),
    .ZN(_11768_));
 BUF_X8 _37943_ (.A(_08495_),
    .Z(_11769_));
 MUX2_X2 _37944_ (.A(_11752_),
    .B(_11768_),
    .S(_11769_),
    .Z(\icache.data_mem_data_li [14]));
 MUX2_X1 _37945_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [277]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [795]),
    .S(_11743_),
    .Z(_11770_));
 AND2_X2 _37946_ (.A1(_11770_),
    .A2(_11671_),
    .ZN(_11771_));
 NAND2_X1 _37947_ (.A1(_11753_),
    .A2(_11771_),
    .ZN(_11772_));
 MUX2_X2 _37948_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [341]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [859]),
    .S(_11743_),
    .Z(_11773_));
 BUF_X4 _37949_ (.A(_11293_),
    .Z(_11774_));
 AND2_X1 _37950_ (.A1(_11773_),
    .A2(_11774_),
    .ZN(_11775_));
 BUF_X4 _37951_ (.A(_11251_),
    .Z(_11776_));
 BUF_X4 _37952_ (.A(_11253_),
    .Z(_11777_));
 OAI21_X2 _37953_ (.A(_11775_),
    .B1(_11776_),
    .B2(_11777_),
    .ZN(_11778_));
 AOI21_X1 _37954_ (.A(_11666_),
    .B1(_11772_),
    .B2(_11778_),
    .ZN(_11779_));
 MUX2_X2 _37955_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [405]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [923]),
    .S(_11743_),
    .Z(_11780_));
 AND2_X2 _37956_ (.A1(_11780_),
    .A2(_11774_),
    .ZN(_11781_));
 NAND2_X1 _37957_ (.A1(_11638_),
    .A2(_11781_),
    .ZN(_11782_));
 MUX2_X2 _37958_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [469]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [987]),
    .S(_11747_),
    .Z(_11783_));
 AND2_X1 _37959_ (.A1(_11783_),
    .A2(_11712_),
    .ZN(_11784_));
 OAI21_X1 _37960_ (.A(_11784_),
    .B1(_11681_),
    .B2(_11683_),
    .ZN(_11785_));
 AOI21_X1 _37961_ (.A(_11710_),
    .B1(_11782_),
    .B2(_11785_),
    .ZN(_11786_));
 OR2_X1 _37962_ (.A1(_11779_),
    .A2(_11786_),
    .ZN(_11787_));
 MUX2_X1 _37963_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [21]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [539]),
    .S(_11448_),
    .Z(_11788_));
 AND2_X4 _37964_ (.A1(_11788_),
    .A2(_11721_),
    .ZN(_11789_));
 NAND2_X1 _37965_ (.A1(_11638_),
    .A2(_11789_),
    .ZN(_11790_));
 MUX2_X2 _37966_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [85]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [603]),
    .S(_11747_),
    .Z(_11791_));
 AND2_X1 _37967_ (.A1(_11791_),
    .A2(_11712_),
    .ZN(_11792_));
 OAI21_X1 _37968_ (.A(_11792_),
    .B1(_11681_),
    .B2(_11683_),
    .ZN(_11793_));
 AOI21_X1 _37969_ (.A(_11547_),
    .B1(_11790_),
    .B2(_11793_),
    .ZN(_11794_));
 MUX2_X2 _37970_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [149]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [667]),
    .S(_11747_),
    .Z(_11795_));
 AND2_X1 _37971_ (.A1(_11795_),
    .A2(_11712_),
    .ZN(_11796_));
 NAND2_X1 _37972_ (.A1(_11753_),
    .A2(_11796_),
    .ZN(_11797_));
 MUX2_X1 _37973_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [213]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [731]),
    .S(_11743_),
    .Z(_11798_));
 AND2_X1 _37974_ (.A1(_11798_),
    .A2(_11671_),
    .ZN(_11799_));
 OAI21_X1 _37975_ (.A(_11799_),
    .B1(_11776_),
    .B2(_11777_),
    .ZN(_11800_));
 AOI21_X1 _37976_ (.A(_11589_),
    .B1(_11797_),
    .B2(_11800_),
    .ZN(_11801_));
 OR2_X1 _37977_ (.A1(_11794_),
    .A2(_11801_),
    .ZN(_11802_));
 MUX2_X2 _37978_ (.A(_11787_),
    .B(_11802_),
    .S(_11769_),
    .Z(\icache.data_mem_data_li [15]));
 MUX2_X1 _37979_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [22]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [540]),
    .S(_11347_),
    .Z(_11803_));
 AND2_X4 _37980_ (.A1(_11803_),
    .A2(_11565_),
    .ZN(_11804_));
 NAND2_X1 _37981_ (.A1(_11753_),
    .A2(_11804_),
    .ZN(_11805_));
 MUX2_X1 _37982_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [86]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [604]),
    .S(_11743_),
    .Z(_11806_));
 AND2_X1 _37983_ (.A1(_11806_),
    .A2(_11774_),
    .ZN(_11807_));
 OAI21_X1 _37984_ (.A(_11807_),
    .B1(_11776_),
    .B2(_11777_),
    .ZN(_11808_));
 AOI21_X1 _37985_ (.A(_11666_),
    .B1(_11805_),
    .B2(_11808_),
    .ZN(_11809_));
 BUF_X4 _37986_ (.A(_11301_),
    .Z(_11810_));
 MUX2_X2 _37987_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [150]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [668]),
    .S(_11747_),
    .Z(_11811_));
 BUF_X4 _37988_ (.A(_11266_),
    .Z(_11812_));
 AND2_X1 _37989_ (.A1(_11811_),
    .A2(_11812_),
    .ZN(_11813_));
 NAND2_X1 _37990_ (.A1(_11810_),
    .A2(_11813_),
    .ZN(_11814_));
 MUX2_X2 _37991_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [214]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [732]),
    .S(_11747_),
    .Z(_11815_));
 AND2_X1 _37992_ (.A1(_11815_),
    .A2(_11812_),
    .ZN(_11816_));
 OAI21_X1 _37993_ (.A(_11816_),
    .B1(_11681_),
    .B2(_11683_),
    .ZN(_11817_));
 AOI21_X1 _37994_ (.A(_11710_),
    .B1(_11814_),
    .B2(_11817_),
    .ZN(_11818_));
 OR2_X1 _37995_ (.A1(_11809_),
    .A2(_11818_),
    .ZN(_11819_));
 MUX2_X1 _37996_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [278]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [796]),
    .S(_11747_),
    .Z(_11820_));
 AND2_X1 _37997_ (.A1(_11820_),
    .A2(_11812_),
    .ZN(_11821_));
 NAND2_X1 _37998_ (.A1(_11810_),
    .A2(_11821_),
    .ZN(_11822_));
 MUX2_X1 _37999_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [342]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [860]),
    .S(_11747_),
    .Z(_11823_));
 AND2_X1 _38000_ (.A1(_11823_),
    .A2(_11812_),
    .ZN(_11824_));
 OAI21_X1 _38001_ (.A(_11824_),
    .B1(_11681_),
    .B2(_11683_),
    .ZN(_11825_));
 AOI21_X1 _38002_ (.A(_11547_),
    .B1(_11822_),
    .B2(_11825_),
    .ZN(_11826_));
 MUX2_X2 _38003_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [406]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [924]),
    .S(_11743_),
    .Z(_11827_));
 AND2_X1 _38004_ (.A1(_11827_),
    .A2(_11774_),
    .ZN(_11828_));
 NAND2_X1 _38005_ (.A1(_11753_),
    .A2(_11828_),
    .ZN(_11829_));
 MUX2_X1 _38006_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [470]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [988]),
    .S(_11743_),
    .Z(_11830_));
 AND2_X1 _38007_ (.A1(_11830_),
    .A2(_11774_),
    .ZN(_11831_));
 OAI21_X1 _38008_ (.A(_11831_),
    .B1(_11776_),
    .B2(_11777_),
    .ZN(_11832_));
 AOI21_X1 _38009_ (.A(_11589_),
    .B1(_11829_),
    .B2(_11832_),
    .ZN(_11833_));
 OR2_X1 _38010_ (.A1(_11826_),
    .A2(_11833_),
    .ZN(_11834_));
 MUX2_X2 _38011_ (.A(_11819_),
    .B(_11834_),
    .S(_08434_),
    .Z(\icache.data_mem_data_li [16]));
 BUF_X16 _38012_ (.A(_08427_),
    .Z(_11835_));
 BUF_X16 _38013_ (.A(_11835_),
    .Z(_11836_));
 MUX2_X2 _38014_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [279]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [797]),
    .S(_11836_),
    .Z(_11837_));
 AND2_X1 _38015_ (.A1(_11837_),
    .A2(_11774_),
    .ZN(_11838_));
 NAND2_X1 _38016_ (.A1(_11753_),
    .A2(_11838_),
    .ZN(_11839_));
 MUX2_X1 _38017_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [343]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [861]),
    .S(_11836_),
    .Z(_11840_));
 AND2_X1 _38018_ (.A1(_11840_),
    .A2(_11774_),
    .ZN(_11841_));
 OAI21_X1 _38019_ (.A(_11841_),
    .B1(_11776_),
    .B2(_11777_),
    .ZN(_11842_));
 AOI21_X1 _38020_ (.A(_11666_),
    .B1(_11839_),
    .B2(_11842_),
    .ZN(_11843_));
 MUX2_X2 _38021_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [407]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [925]),
    .S(_11747_),
    .Z(_11844_));
 AND2_X1 _38022_ (.A1(_11844_),
    .A2(_11812_),
    .ZN(_11845_));
 NAND2_X1 _38023_ (.A1(_11810_),
    .A2(_11845_),
    .ZN(_11846_));
 BUF_X8 _38024_ (.A(_11643_),
    .Z(_11847_));
 MUX2_X1 _38025_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [471]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [989]),
    .S(_11847_),
    .Z(_11848_));
 AND2_X1 _38026_ (.A1(_11848_),
    .A2(_11812_),
    .ZN(_11849_));
 BUF_X4 _38027_ (.A(_11680_),
    .Z(_11850_));
 BUF_X4 _38028_ (.A(_11682_),
    .Z(_11851_));
 OAI21_X1 _38029_ (.A(_11849_),
    .B1(_11850_),
    .B2(_11851_),
    .ZN(_11852_));
 AOI21_X1 _38030_ (.A(_11710_),
    .B1(_11846_),
    .B2(_11852_),
    .ZN(_11853_));
 OR2_X1 _38031_ (.A1(_11843_),
    .A2(_11853_),
    .ZN(_11854_));
 MUX2_X1 _38032_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [23]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [541]),
    .S(_11448_),
    .Z(_11855_));
 AND2_X4 _38033_ (.A1(_11855_),
    .A2(_11721_),
    .ZN(_11856_));
 NAND2_X1 _38034_ (.A1(_11810_),
    .A2(_11856_),
    .ZN(_11857_));
 MUX2_X2 _38035_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [87]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [605]),
    .S(_11747_),
    .Z(_11858_));
 AND2_X1 _38036_ (.A1(_11858_),
    .A2(_11812_),
    .ZN(_11859_));
 OAI21_X1 _38037_ (.A(_11859_),
    .B1(_11850_),
    .B2(_11851_),
    .ZN(_11860_));
 AOI21_X1 _38038_ (.A(_11547_),
    .B1(_11857_),
    .B2(_11860_),
    .ZN(_11861_));
 MUX2_X1 _38039_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [151]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [669]),
    .S(_11743_),
    .Z(_11862_));
 AND2_X2 _38040_ (.A1(_11862_),
    .A2(_11774_),
    .ZN(_11863_));
 NAND2_X1 _38041_ (.A1(_11753_),
    .A2(_11863_),
    .ZN(_11864_));
 MUX2_X2 _38042_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [215]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [733]),
    .S(_11836_),
    .Z(_11865_));
 AND2_X1 _38043_ (.A1(_11865_),
    .A2(_11774_),
    .ZN(_11866_));
 OAI21_X1 _38044_ (.A(_11866_),
    .B1(_11776_),
    .B2(_11777_),
    .ZN(_11867_));
 AOI21_X1 _38045_ (.A(_11589_),
    .B1(_11864_),
    .B2(_11867_),
    .ZN(_11868_));
 OR2_X1 _38046_ (.A1(_11861_),
    .A2(_11868_),
    .ZN(_11869_));
 MUX2_X2 _38047_ (.A(_11854_),
    .B(_11869_),
    .S(_11769_),
    .Z(\icache.data_mem_data_li [17]));
 MUX2_X2 _38048_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [280]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [798]),
    .S(_11847_),
    .Z(_11870_));
 AND2_X1 _38049_ (.A1(_11870_),
    .A2(_11812_),
    .ZN(_11871_));
 NAND2_X1 _38050_ (.A1(_11810_),
    .A2(_11871_),
    .ZN(_11872_));
 MUX2_X1 _38051_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [344]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [862]),
    .S(_11847_),
    .Z(_11873_));
 AND2_X1 _38052_ (.A1(_11873_),
    .A2(_11812_),
    .ZN(_11874_));
 OAI21_X1 _38053_ (.A(_11874_),
    .B1(_11850_),
    .B2(_11851_),
    .ZN(_11875_));
 AOI21_X1 _38054_ (.A(_11666_),
    .B1(_11872_),
    .B2(_11875_),
    .ZN(_11876_));
 MUX2_X1 _38055_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [408]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [926]),
    .S(_11847_),
    .Z(_11877_));
 AND2_X1 _38056_ (.A1(_11877_),
    .A2(_11812_),
    .ZN(_11878_));
 NAND2_X1 _38057_ (.A1(_11810_),
    .A2(_11878_),
    .ZN(_11879_));
 MUX2_X1 _38058_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [472]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [990]),
    .S(_11847_),
    .Z(_11880_));
 BUF_X2 _38059_ (.A(_11266_),
    .Z(_11881_));
 AND2_X1 _38060_ (.A1(_11880_),
    .A2(_11881_),
    .ZN(_11882_));
 OAI21_X1 _38061_ (.A(_11882_),
    .B1(_11850_),
    .B2(_11851_),
    .ZN(_11883_));
 AOI21_X1 _38062_ (.A(_11710_),
    .B1(_11879_),
    .B2(_11883_),
    .ZN(_11884_));
 OR2_X1 _38063_ (.A1(_11876_),
    .A2(_11884_),
    .ZN(_11885_));
 BUF_X8 _38064_ (.A(_11546_),
    .Z(_11886_));
 MUX2_X1 _38065_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [24]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [542]),
    .S(_11347_),
    .Z(_11887_));
 AND2_X4 _38066_ (.A1(_11887_),
    .A2(_11565_),
    .ZN(_11888_));
 NAND2_X1 _38067_ (.A1(_11753_),
    .A2(_11888_),
    .ZN(_11889_));
 MUX2_X1 _38068_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [88]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [606]),
    .S(_11836_),
    .Z(_11890_));
 AND2_X2 _38069_ (.A1(_11890_),
    .A2(_11774_),
    .ZN(_11891_));
 OAI21_X1 _38070_ (.A(_11891_),
    .B1(_11776_),
    .B2(_11777_),
    .ZN(_11892_));
 AOI21_X1 _38071_ (.A(_11886_),
    .B1(_11889_),
    .B2(_11892_),
    .ZN(_11893_));
 MUX2_X2 _38072_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [152]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [670]),
    .S(_11836_),
    .Z(_11894_));
 BUF_X4 _38073_ (.A(_11293_),
    .Z(_11895_));
 AND2_X2 _38074_ (.A1(_11894_),
    .A2(_11895_),
    .ZN(_11896_));
 NAND2_X1 _38075_ (.A1(_11753_),
    .A2(_11896_),
    .ZN(_11897_));
 MUX2_X2 _38076_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [216]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [734]),
    .S(_11836_),
    .Z(_11898_));
 AND2_X1 _38077_ (.A1(_11898_),
    .A2(_11895_),
    .ZN(_11899_));
 OAI21_X1 _38078_ (.A(_11899_),
    .B1(_11776_),
    .B2(_11777_),
    .ZN(_11900_));
 AOI21_X1 _38079_ (.A(_11589_),
    .B1(_11897_),
    .B2(_11900_),
    .ZN(_11901_));
 OR2_X1 _38080_ (.A1(_11893_),
    .A2(_11901_),
    .ZN(_11902_));
 MUX2_X2 _38081_ (.A(_11885_),
    .B(_11902_),
    .S(_11769_),
    .Z(\icache.data_mem_data_li [18]));
 MUX2_X1 _38082_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [281]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [799]),
    .S(_11847_),
    .Z(_11903_));
 AND2_X1 _38083_ (.A1(_11903_),
    .A2(_11881_),
    .ZN(_11904_));
 NAND2_X1 _38084_ (.A1(_11810_),
    .A2(_11904_),
    .ZN(_11905_));
 MUX2_X1 _38085_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [345]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [863]),
    .S(_11847_),
    .Z(_11906_));
 AND2_X1 _38086_ (.A1(_11906_),
    .A2(_11881_),
    .ZN(_11907_));
 OAI21_X1 _38087_ (.A(_11907_),
    .B1(_11850_),
    .B2(_11851_),
    .ZN(_11908_));
 AOI21_X1 _38088_ (.A(_11666_),
    .B1(_11905_),
    .B2(_11908_),
    .ZN(_11909_));
 MUX2_X2 _38089_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [409]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [927]),
    .S(_11847_),
    .Z(_11910_));
 AND2_X1 _38090_ (.A1(_11910_),
    .A2(_11881_),
    .ZN(_11911_));
 NAND2_X1 _38091_ (.A1(_11810_),
    .A2(_11911_),
    .ZN(_11912_));
 MUX2_X1 _38092_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [473]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [991]),
    .S(_11847_),
    .Z(_11913_));
 AND2_X1 _38093_ (.A1(_11913_),
    .A2(_11881_),
    .ZN(_11914_));
 OAI21_X1 _38094_ (.A(_11914_),
    .B1(_11850_),
    .B2(_11851_),
    .ZN(_11915_));
 AOI21_X1 _38095_ (.A(_11710_),
    .B1(_11912_),
    .B2(_11915_),
    .ZN(_11916_));
 OR2_X2 _38096_ (.A1(_11909_),
    .A2(_11916_),
    .ZN(_11917_));
 BUF_X4 _38097_ (.A(_11413_),
    .Z(_11918_));
 BUF_X16 _38098_ (.A(_08427_),
    .Z(_11919_));
 MUX2_X2 _38099_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [25]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [543]),
    .S(_11919_),
    .Z(_11920_));
 AND2_X4 _38100_ (.A1(_11920_),
    .A2(_11565_),
    .ZN(_11921_));
 NAND2_X1 _38101_ (.A1(_11918_),
    .A2(_11921_),
    .ZN(_11922_));
 MUX2_X1 _38102_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [89]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [607]),
    .S(_11836_),
    .Z(_11923_));
 AND2_X2 _38103_ (.A1(_11923_),
    .A2(_11895_),
    .ZN(_11924_));
 OAI21_X1 _38104_ (.A(_11924_),
    .B1(_11776_),
    .B2(_11777_),
    .ZN(_11925_));
 AOI21_X1 _38105_ (.A(_11886_),
    .B1(_11922_),
    .B2(_11925_),
    .ZN(_11926_));
 BUF_X8 _38106_ (.A(_08493_),
    .Z(_11927_));
 MUX2_X1 _38107_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [153]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [671]),
    .S(_11836_),
    .Z(_11928_));
 AND2_X1 _38108_ (.A1(_11928_),
    .A2(_11895_),
    .ZN(_11929_));
 NAND2_X1 _38109_ (.A1(_11918_),
    .A2(_11929_),
    .ZN(_11930_));
 MUX2_X2 _38110_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [217]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [735]),
    .S(_11836_),
    .Z(_11931_));
 AND2_X2 _38111_ (.A1(_11931_),
    .A2(_11895_),
    .ZN(_11932_));
 OAI21_X1 _38112_ (.A(_11932_),
    .B1(_11776_),
    .B2(_11777_),
    .ZN(_11933_));
 AOI21_X1 _38113_ (.A(_11927_),
    .B1(_11930_),
    .B2(_11933_),
    .ZN(_11934_));
 OR2_X1 _38114_ (.A1(_11926_),
    .A2(_11934_),
    .ZN(_11935_));
 MUX2_X2 _38115_ (.A(_11917_),
    .B(_11935_),
    .S(_11769_),
    .Z(\icache.data_mem_data_li [19]));
 MUX2_X1 _38116_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [26]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [544]),
    .S(_11919_),
    .Z(_11936_));
 AND2_X4 _38117_ (.A1(_11936_),
    .A2(_11565_),
    .ZN(_11937_));
 NAND2_X1 _38118_ (.A1(_11918_),
    .A2(_11937_),
    .ZN(_11938_));
 BUF_X8 _38119_ (.A(_11835_),
    .Z(_11939_));
 MUX2_X1 _38120_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [90]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [608]),
    .S(_11939_),
    .Z(_11940_));
 AND2_X1 _38121_ (.A1(_11940_),
    .A2(_11895_),
    .ZN(_11941_));
 BUF_X4 _38122_ (.A(_11251_),
    .Z(_11942_));
 BUF_X4 _38123_ (.A(_11253_),
    .Z(_11943_));
 OAI21_X1 _38124_ (.A(_11941_),
    .B1(_11942_),
    .B2(_11943_),
    .ZN(_11944_));
 AOI21_X1 _38125_ (.A(_11666_),
    .B1(_11938_),
    .B2(_11944_),
    .ZN(_11945_));
 BUF_X16 _38126_ (.A(_11643_),
    .Z(_11946_));
 MUX2_X1 _38127_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [154]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [672]),
    .S(_11946_),
    .Z(_11947_));
 AND2_X1 _38128_ (.A1(_11947_),
    .A2(_11881_),
    .ZN(_11948_));
 NAND2_X1 _38129_ (.A1(_11810_),
    .A2(_11948_),
    .ZN(_11949_));
 MUX2_X2 _38130_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [218]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [736]),
    .S(_11946_),
    .Z(_11950_));
 AND2_X1 _38131_ (.A1(_11950_),
    .A2(_11881_),
    .ZN(_11951_));
 OAI21_X2 _38132_ (.A(_11951_),
    .B1(_11850_),
    .B2(_11851_),
    .ZN(_11952_));
 AOI21_X1 _38133_ (.A(_11710_),
    .B1(_11949_),
    .B2(_11952_),
    .ZN(_11953_));
 OR2_X2 _38134_ (.A1(_11945_),
    .A2(_11953_),
    .ZN(_11954_));
 MUX2_X1 _38135_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [282]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [800]),
    .S(_11847_),
    .Z(_11955_));
 AND2_X1 _38136_ (.A1(_11955_),
    .A2(_11881_),
    .ZN(_11956_));
 NAND2_X1 _38137_ (.A1(_11810_),
    .A2(_11956_),
    .ZN(_11957_));
 MUX2_X1 _38138_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [346]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [864]),
    .S(_11946_),
    .Z(_11958_));
 AND2_X1 _38139_ (.A1(_11958_),
    .A2(_11881_),
    .ZN(_11959_));
 OAI21_X1 _38140_ (.A(_11959_),
    .B1(_11850_),
    .B2(_11851_),
    .ZN(_11960_));
 AOI21_X1 _38141_ (.A(_11886_),
    .B1(_11957_),
    .B2(_11960_),
    .ZN(_11961_));
 MUX2_X2 _38142_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [410]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [928]),
    .S(_11836_),
    .Z(_11962_));
 AND2_X1 _38143_ (.A1(_11962_),
    .A2(_11895_),
    .ZN(_11963_));
 NAND2_X1 _38144_ (.A1(_11918_),
    .A2(_11963_),
    .ZN(_11964_));
 MUX2_X1 _38145_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [474]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [992]),
    .S(_11939_),
    .Z(_11965_));
 AND2_X1 _38146_ (.A1(_11965_),
    .A2(_11895_),
    .ZN(_11966_));
 OAI21_X1 _38147_ (.A(_11966_),
    .B1(_11942_),
    .B2(_11943_),
    .ZN(_11967_));
 AOI21_X1 _38148_ (.A(_11927_),
    .B1(_11964_),
    .B2(_11967_),
    .ZN(_11968_));
 OR2_X2 _38149_ (.A1(_11961_),
    .A2(_11968_),
    .ZN(_11969_));
 MUX2_X2 _38150_ (.A(_11954_),
    .B(_11969_),
    .S(_08434_),
    .Z(\icache.data_mem_data_li [20]));
 BUF_X4 _38151_ (.A(_11301_),
    .Z(_11970_));
 MUX2_X2 _38152_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [283]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [801]),
    .S(_11946_),
    .Z(_11971_));
 AND2_X1 _38153_ (.A1(_11971_),
    .A2(_11881_),
    .ZN(_11972_));
 NAND2_X1 _38154_ (.A1(_11970_),
    .A2(_11972_),
    .ZN(_11973_));
 MUX2_X1 _38155_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [347]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [865]),
    .S(_11946_),
    .Z(_11974_));
 BUF_X4 _38156_ (.A(_11266_),
    .Z(_11975_));
 AND2_X1 _38157_ (.A1(_11974_),
    .A2(_11975_),
    .ZN(_11976_));
 OAI21_X1 _38158_ (.A(_11976_),
    .B1(_11850_),
    .B2(_11851_),
    .ZN(_11977_));
 AOI21_X1 _38159_ (.A(_11666_),
    .B1(_11973_),
    .B2(_11977_),
    .ZN(_11978_));
 MUX2_X2 _38160_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [411]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [929]),
    .S(_11946_),
    .Z(_11979_));
 AND2_X1 _38161_ (.A1(_11979_),
    .A2(_11975_),
    .ZN(_11980_));
 NAND2_X1 _38162_ (.A1(_11970_),
    .A2(_11980_),
    .ZN(_11981_));
 MUX2_X2 _38163_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [475]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [993]),
    .S(_11946_),
    .Z(_11982_));
 AND2_X1 _38164_ (.A1(_11982_),
    .A2(_11975_),
    .ZN(_11983_));
 OAI21_X1 _38165_ (.A(_11983_),
    .B1(_11850_),
    .B2(_11851_),
    .ZN(_11984_));
 AOI21_X1 _38166_ (.A(_11710_),
    .B1(_11981_),
    .B2(_11984_),
    .ZN(_11985_));
 OR2_X2 _38167_ (.A1(_11978_),
    .A2(_11985_),
    .ZN(_11986_));
 MUX2_X2 _38168_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [27]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [545]),
    .S(_11919_),
    .Z(_11987_));
 AND2_X4 _38169_ (.A1(_11987_),
    .A2(_11565_),
    .ZN(_11988_));
 NAND2_X1 _38170_ (.A1(_11918_),
    .A2(_11988_),
    .ZN(_11989_));
 MUX2_X1 _38171_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [91]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [609]),
    .S(_11939_),
    .Z(_11990_));
 AND2_X2 _38172_ (.A1(_11990_),
    .A2(_11895_),
    .ZN(_11991_));
 OAI21_X1 _38173_ (.A(_11991_),
    .B1(_11942_),
    .B2(_11943_),
    .ZN(_11992_));
 AOI21_X1 _38174_ (.A(_11886_),
    .B1(_11989_),
    .B2(_11992_),
    .ZN(_11993_));
 MUX2_X1 _38175_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [155]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [673]),
    .S(_11939_),
    .Z(_11994_));
 AND2_X4 _38176_ (.A1(_11994_),
    .A2(_11895_),
    .ZN(_11995_));
 NAND2_X1 _38177_ (.A1(_11918_),
    .A2(_11995_),
    .ZN(_11996_));
 MUX2_X2 _38178_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [219]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [737]),
    .S(_11939_),
    .Z(_11997_));
 BUF_X2 _38179_ (.A(_11293_),
    .Z(_11998_));
 AND2_X1 _38180_ (.A1(_11997_),
    .A2(_11998_),
    .ZN(_11999_));
 OAI21_X1 _38181_ (.A(_11999_),
    .B1(_11942_),
    .B2(_11943_),
    .ZN(_12000_));
 AOI21_X1 _38182_ (.A(_11927_),
    .B1(_11996_),
    .B2(_12000_),
    .ZN(_12001_));
 OR2_X2 _38183_ (.A1(_11993_),
    .A2(_12001_),
    .ZN(_12002_));
 MUX2_X2 _38184_ (.A(_11986_),
    .B(_12002_),
    .S(_11769_),
    .Z(\icache.data_mem_data_li [21]));
 BUF_X8 _38185_ (.A(_11665_),
    .Z(_12003_));
 MUX2_X1 _38186_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [28]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [546]),
    .S(_11448_),
    .Z(_12004_));
 AND2_X4 _38187_ (.A1(_12004_),
    .A2(_11721_),
    .ZN(_12005_));
 NAND2_X1 _38188_ (.A1(_11970_),
    .A2(_12005_),
    .ZN(_12006_));
 MUX2_X1 _38189_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [92]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [610]),
    .S(_11946_),
    .Z(_12007_));
 AND2_X1 _38190_ (.A1(_12007_),
    .A2(_11975_),
    .ZN(_12008_));
 BUF_X4 _38191_ (.A(_11680_),
    .Z(_12009_));
 BUF_X4 _38192_ (.A(_11682_),
    .Z(_12010_));
 OAI21_X1 _38193_ (.A(_12008_),
    .B1(_12009_),
    .B2(_12010_),
    .ZN(_12011_));
 AOI21_X1 _38194_ (.A(_12003_),
    .B1(_12006_),
    .B2(_12011_),
    .ZN(_12012_));
 MUX2_X2 _38195_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [156]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [674]),
    .S(_11939_),
    .Z(_12013_));
 AND2_X1 _38196_ (.A1(_12013_),
    .A2(_11998_),
    .ZN(_12014_));
 NAND2_X1 _38197_ (.A1(_11970_),
    .A2(_12014_),
    .ZN(_12015_));
 MUX2_X2 _38198_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [220]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [738]),
    .S(_11946_),
    .Z(_12016_));
 AND2_X1 _38199_ (.A1(_12016_),
    .A2(_11975_),
    .ZN(_12017_));
 OAI21_X1 _38200_ (.A(_12017_),
    .B1(_12009_),
    .B2(_12010_),
    .ZN(_12018_));
 AOI21_X1 _38201_ (.A(_11710_),
    .B1(_12015_),
    .B2(_12018_),
    .ZN(_12019_));
 OR2_X4 _38202_ (.A1(_12012_),
    .A2(_12019_),
    .ZN(_12020_));
 MUX2_X1 _38203_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [284]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [802]),
    .S(_11939_),
    .Z(_12021_));
 AND2_X1 _38204_ (.A1(_12021_),
    .A2(_11998_),
    .ZN(_12022_));
 NAND2_X1 _38205_ (.A1(_11918_),
    .A2(_12022_),
    .ZN(_12023_));
 MUX2_X2 _38206_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [348]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [866]),
    .S(_11939_),
    .Z(_12024_));
 AND2_X1 _38207_ (.A1(_12024_),
    .A2(_11998_),
    .ZN(_12025_));
 OAI21_X1 _38208_ (.A(_12025_),
    .B1(_11942_),
    .B2(_11943_),
    .ZN(_12026_));
 AOI21_X1 _38209_ (.A(_11886_),
    .B1(_12023_),
    .B2(_12026_),
    .ZN(_12027_));
 MUX2_X2 _38210_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [412]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [930]),
    .S(_11946_),
    .Z(_12028_));
 AND2_X1 _38211_ (.A1(_12028_),
    .A2(_11975_),
    .ZN(_12029_));
 NAND2_X1 _38212_ (.A1(_11918_),
    .A2(_12029_),
    .ZN(_12030_));
 MUX2_X2 _38213_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [476]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [994]),
    .S(_11939_),
    .Z(_12031_));
 AND2_X1 _38214_ (.A1(_12031_),
    .A2(_11998_),
    .ZN(_12032_));
 OAI21_X1 _38215_ (.A(_12032_),
    .B1(_11942_),
    .B2(_11943_),
    .ZN(_12033_));
 AOI21_X1 _38216_ (.A(_11927_),
    .B1(_12030_),
    .B2(_12033_),
    .ZN(_12034_));
 OR2_X2 _38217_ (.A1(_12027_),
    .A2(_12034_),
    .ZN(_12035_));
 MUX2_X2 _38218_ (.A(_12020_),
    .B(_12035_),
    .S(_08434_),
    .Z(\icache.data_mem_data_li [22]));
 BUF_X8 _38219_ (.A(_11643_),
    .Z(_12036_));
 MUX2_X1 _38220_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [285]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [803]),
    .S(_12036_),
    .Z(_12037_));
 AND2_X1 _38221_ (.A1(_12037_),
    .A2(_11975_),
    .ZN(_12038_));
 NAND2_X1 _38222_ (.A1(_11970_),
    .A2(_12038_),
    .ZN(_12039_));
 MUX2_X1 _38223_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [349]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [867]),
    .S(_12036_),
    .Z(_12040_));
 AND2_X1 _38224_ (.A1(_12040_),
    .A2(_11975_),
    .ZN(_12041_));
 OAI21_X1 _38225_ (.A(_12041_),
    .B1(_12009_),
    .B2(_12010_),
    .ZN(_12042_));
 AOI21_X1 _38226_ (.A(_12003_),
    .B1(_12039_),
    .B2(_12042_),
    .ZN(_12043_));
 BUF_X8 _38227_ (.A(_11709_),
    .Z(_12044_));
 MUX2_X2 _38228_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [413]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [931]),
    .S(_12036_),
    .Z(_12045_));
 AND2_X1 _38229_ (.A1(_12045_),
    .A2(_11975_),
    .ZN(_12046_));
 NAND2_X1 _38230_ (.A1(_11970_),
    .A2(_12046_),
    .ZN(_12047_));
 MUX2_X1 _38231_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [477]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [995]),
    .S(_12036_),
    .Z(_12048_));
 AND2_X2 _38232_ (.A1(_12048_),
    .A2(_11975_),
    .ZN(_12049_));
 OAI21_X1 _38233_ (.A(_12049_),
    .B1(_12009_),
    .B2(_12010_),
    .ZN(_12050_));
 AOI21_X1 _38234_ (.A(_12044_),
    .B1(_12047_),
    .B2(_12050_),
    .ZN(_12051_));
 OR2_X4 _38235_ (.A1(_12043_),
    .A2(_12051_),
    .ZN(_12052_));
 MUX2_X1 _38236_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [29]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [547]),
    .S(_11919_),
    .Z(_12053_));
 AND2_X4 _38237_ (.A1(_12053_),
    .A2(_11565_),
    .ZN(_12054_));
 NAND2_X1 _38238_ (.A1(_11918_),
    .A2(_12054_),
    .ZN(_12055_));
 MUX2_X1 _38239_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [93]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [611]),
    .S(_11939_),
    .Z(_12056_));
 AND2_X1 _38240_ (.A1(_12056_),
    .A2(_11998_),
    .ZN(_12057_));
 OAI21_X1 _38241_ (.A(_12057_),
    .B1(_11942_),
    .B2(_11943_),
    .ZN(_12058_));
 AOI21_X1 _38242_ (.A(_11886_),
    .B1(_12055_),
    .B2(_12058_),
    .ZN(_12059_));
 BUF_X8 _38243_ (.A(_11835_),
    .Z(_12060_));
 MUX2_X1 _38244_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [157]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [675]),
    .S(_12060_),
    .Z(_12061_));
 AND2_X1 _38245_ (.A1(_12061_),
    .A2(_11998_),
    .ZN(_12062_));
 NAND2_X1 _38246_ (.A1(_11918_),
    .A2(_12062_),
    .ZN(_12063_));
 MUX2_X2 _38247_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [221]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [739]),
    .S(_12060_),
    .Z(_12064_));
 AND2_X1 _38248_ (.A1(_12064_),
    .A2(_11998_),
    .ZN(_12065_));
 OAI21_X1 _38249_ (.A(_12065_),
    .B1(_11942_),
    .B2(_11943_),
    .ZN(_12066_));
 AOI21_X1 _38250_ (.A(_11927_),
    .B1(_12063_),
    .B2(_12066_),
    .ZN(_12067_));
 OR2_X4 _38251_ (.A1(_12059_),
    .A2(_12067_),
    .ZN(_12068_));
 MUX2_X2 _38252_ (.A(_12052_),
    .B(_12068_),
    .S(_11769_),
    .Z(\icache.data_mem_data_li [23]));
 BUF_X4 _38253_ (.A(_11413_),
    .Z(_12069_));
 MUX2_X1 _38254_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [286]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [804]),
    .S(_12060_),
    .Z(_12070_));
 BUF_X4 _38255_ (.A(_11293_),
    .Z(_12071_));
 AND2_X1 _38256_ (.A1(_12070_),
    .A2(_12071_),
    .ZN(_12072_));
 NAND2_X1 _38257_ (.A1(_12069_),
    .A2(_12072_),
    .ZN(_12073_));
 MUX2_X1 _38258_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [350]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [868]),
    .S(_12060_),
    .Z(_12074_));
 AND2_X2 _38259_ (.A1(_12074_),
    .A2(_12071_),
    .ZN(_12075_));
 OAI21_X1 _38260_ (.A(_12075_),
    .B1(_11942_),
    .B2(_11943_),
    .ZN(_12076_));
 AOI21_X1 _38261_ (.A(_12003_),
    .B1(_12073_),
    .B2(_12076_),
    .ZN(_12077_));
 MUX2_X1 _38262_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [414]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [932]),
    .S(_12036_),
    .Z(_12078_));
 BUF_X16 _38263_ (.A(_08426_),
    .Z(_12079_));
 BUF_X2 _38264_ (.A(_12079_),
    .Z(_12080_));
 AND2_X1 _38265_ (.A1(_12078_),
    .A2(_12080_),
    .ZN(_12081_));
 NAND2_X1 _38266_ (.A1(_11970_),
    .A2(_12081_),
    .ZN(_12082_));
 MUX2_X2 _38267_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [478]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [996]),
    .S(_12036_),
    .Z(_12083_));
 AND2_X1 _38268_ (.A1(_12083_),
    .A2(_12080_),
    .ZN(_12084_));
 OAI21_X1 _38269_ (.A(_12084_),
    .B1(_12009_),
    .B2(_12010_),
    .ZN(_12085_));
 AOI21_X1 _38270_ (.A(_12044_),
    .B1(_12082_),
    .B2(_12085_),
    .ZN(_12086_));
 OR2_X4 _38271_ (.A1(_12077_),
    .A2(_12086_),
    .ZN(_12087_));
 MUX2_X1 _38272_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [30]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [548]),
    .S(_11448_),
    .Z(_12088_));
 AND2_X4 _38273_ (.A1(_12088_),
    .A2(_11721_),
    .ZN(_12089_));
 NAND2_X1 _38274_ (.A1(_11970_),
    .A2(_12089_),
    .ZN(_12090_));
 MUX2_X1 _38275_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [94]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [612]),
    .S(_12036_),
    .Z(_12091_));
 AND2_X1 _38276_ (.A1(_12091_),
    .A2(_12080_),
    .ZN(_12092_));
 OAI21_X1 _38277_ (.A(_12092_),
    .B1(_12009_),
    .B2(_12010_),
    .ZN(_12093_));
 AOI21_X1 _38278_ (.A(_11886_),
    .B1(_12090_),
    .B2(_12093_),
    .ZN(_12094_));
 MUX2_X1 _38279_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [158]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [676]),
    .S(_12060_),
    .Z(_12095_));
 AND2_X2 _38280_ (.A1(_12095_),
    .A2(_11998_),
    .ZN(_12096_));
 NAND2_X1 _38281_ (.A1(_12069_),
    .A2(_12096_),
    .ZN(_12097_));
 MUX2_X1 _38282_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [222]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [740]),
    .S(_12060_),
    .Z(_12098_));
 AND2_X1 _38283_ (.A1(_12098_),
    .A2(_11998_),
    .ZN(_12099_));
 OAI21_X1 _38284_ (.A(_12099_),
    .B1(_11942_),
    .B2(_11943_),
    .ZN(_12100_));
 AOI21_X1 _38285_ (.A(_11927_),
    .B1(_12097_),
    .B2(_12100_),
    .ZN(_12101_));
 OR2_X4 _38286_ (.A1(_12094_),
    .A2(_12101_),
    .ZN(_12102_));
 MUX2_X2 _38287_ (.A(_12087_),
    .B(_12102_),
    .S(_11769_),
    .Z(\icache.data_mem_data_li [24]));
 MUX2_X2 _38288_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [287]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [805]),
    .S(_12036_),
    .Z(_12103_));
 AND2_X1 _38289_ (.A1(_12103_),
    .A2(_12080_),
    .ZN(_12104_));
 NAND2_X1 _38290_ (.A1(_11970_),
    .A2(_12104_),
    .ZN(_12105_));
 MUX2_X2 _38291_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [351]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [869]),
    .S(_12036_),
    .Z(_12106_));
 AND2_X1 _38292_ (.A1(_12106_),
    .A2(_12080_),
    .ZN(_12107_));
 OAI21_X1 _38293_ (.A(_12107_),
    .B1(_12009_),
    .B2(_12010_),
    .ZN(_12108_));
 AOI21_X1 _38294_ (.A(_12003_),
    .B1(_12105_),
    .B2(_12108_),
    .ZN(_12109_));
 MUX2_X2 _38295_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [415]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [933]),
    .S(_12060_),
    .Z(_12110_));
 AND2_X1 _38296_ (.A1(_12110_),
    .A2(_12071_),
    .ZN(_12111_));
 NAND2_X1 _38297_ (.A1(_11970_),
    .A2(_12111_),
    .ZN(_12112_));
 BUF_X8 _38298_ (.A(_11643_),
    .Z(_12113_));
 MUX2_X2 _38299_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [479]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [997]),
    .S(_12113_),
    .Z(_12114_));
 AND2_X1 _38300_ (.A1(_12114_),
    .A2(_12080_),
    .ZN(_12115_));
 OAI21_X1 _38301_ (.A(_12115_),
    .B1(_12009_),
    .B2(_12010_),
    .ZN(_12116_));
 AOI21_X1 _38302_ (.A(_12044_),
    .B1(_12112_),
    .B2(_12116_),
    .ZN(_12117_));
 OR2_X4 _38303_ (.A1(_12109_),
    .A2(_12117_),
    .ZN(_12118_));
 MUX2_X2 _38304_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [31]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [549]),
    .S(_11919_),
    .Z(_12119_));
 BUF_X16 _38305_ (.A(_11244_),
    .Z(_12120_));
 AND2_X4 _38306_ (.A1(_12119_),
    .A2(_12120_),
    .ZN(_12121_));
 NAND2_X1 _38307_ (.A1(_12069_),
    .A2(_12121_),
    .ZN(_12122_));
 MUX2_X2 _38308_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [95]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [613]),
    .S(_12060_),
    .Z(_12123_));
 AND2_X2 _38309_ (.A1(_12123_),
    .A2(_12071_),
    .ZN(_12124_));
 BUF_X2 _38310_ (.A(_11251_),
    .Z(_12125_));
 BUF_X2 _38311_ (.A(_11253_),
    .Z(_12126_));
 OAI21_X1 _38312_ (.A(_12124_),
    .B1(_12125_),
    .B2(_12126_),
    .ZN(_12127_));
 AOI21_X1 _38313_ (.A(_11886_),
    .B1(_12122_),
    .B2(_12127_),
    .ZN(_12128_));
 MUX2_X1 _38314_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [159]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [677]),
    .S(_12036_),
    .Z(_12129_));
 AND2_X1 _38315_ (.A1(_12129_),
    .A2(_12080_),
    .ZN(_12130_));
 NAND2_X1 _38316_ (.A1(_12069_),
    .A2(_12130_),
    .ZN(_12131_));
 MUX2_X2 _38317_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [223]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [741]),
    .S(_12060_),
    .Z(_12132_));
 AND2_X2 _38318_ (.A1(_12132_),
    .A2(_12071_),
    .ZN(_12133_));
 OAI21_X1 _38319_ (.A(_12133_),
    .B1(_12125_),
    .B2(_12126_),
    .ZN(_12134_));
 AOI21_X1 _38320_ (.A(_11927_),
    .B1(_12131_),
    .B2(_12134_),
    .ZN(_12135_));
 OR2_X4 _38321_ (.A1(_12128_),
    .A2(_12135_),
    .ZN(_12136_));
 MUX2_X2 _38322_ (.A(_12118_),
    .B(_12136_),
    .S(_11769_),
    .Z(\icache.data_mem_data_li [25]));
 BUF_X4 _38323_ (.A(_11301_),
    .Z(_12137_));
 MUX2_X1 _38324_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [288]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [806]),
    .S(_12113_),
    .Z(_12138_));
 AND2_X2 _38325_ (.A1(_12138_),
    .A2(_12080_),
    .ZN(_12139_));
 NAND2_X1 _38326_ (.A1(_12137_),
    .A2(_12139_),
    .ZN(_12140_));
 MUX2_X1 _38327_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [352]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [870]),
    .S(_12113_),
    .Z(_12141_));
 AND2_X1 _38328_ (.A1(_12141_),
    .A2(_12080_),
    .ZN(_12142_));
 OAI21_X1 _38329_ (.A(_12142_),
    .B1(_12009_),
    .B2(_12010_),
    .ZN(_12143_));
 AOI21_X1 _38330_ (.A(_12003_),
    .B1(_12140_),
    .B2(_12143_),
    .ZN(_12144_));
 BUF_X8 _38331_ (.A(_11835_),
    .Z(_12145_));
 MUX2_X1 _38332_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [416]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [934]),
    .S(_12145_),
    .Z(_12146_));
 AND2_X1 _38333_ (.A1(_12146_),
    .A2(_12071_),
    .ZN(_12147_));
 NAND2_X1 _38334_ (.A1(_12137_),
    .A2(_12147_),
    .ZN(_12148_));
 MUX2_X2 _38335_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [480]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [998]),
    .S(_12113_),
    .Z(_12149_));
 BUF_X4 _38336_ (.A(_12079_),
    .Z(_12150_));
 AND2_X1 _38337_ (.A1(_12149_),
    .A2(_12150_),
    .ZN(_12151_));
 OAI21_X1 _38338_ (.A(_12151_),
    .B1(_12009_),
    .B2(_12010_),
    .ZN(_12152_));
 AOI21_X1 _38339_ (.A(_12044_),
    .B1(_12148_),
    .B2(_12152_),
    .ZN(_12153_));
 OR2_X4 _38340_ (.A1(_12144_),
    .A2(_12153_),
    .ZN(_12154_));
 MUX2_X2 _38341_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [32]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [550]),
    .S(_11919_),
    .Z(_12155_));
 AND2_X4 _38342_ (.A1(_12155_),
    .A2(_12120_),
    .ZN(_12156_));
 NAND2_X1 _38343_ (.A1(_12069_),
    .A2(_12156_),
    .ZN(_12157_));
 MUX2_X2 _38344_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [96]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [614]),
    .S(_12060_),
    .Z(_12158_));
 AND2_X1 _38345_ (.A1(_12158_),
    .A2(_12071_),
    .ZN(_12159_));
 OAI21_X1 _38346_ (.A(_12159_),
    .B1(_12125_),
    .B2(_12126_),
    .ZN(_12160_));
 AOI21_X1 _38347_ (.A(_11886_),
    .B1(_12157_),
    .B2(_12160_),
    .ZN(_12161_));
 MUX2_X2 _38348_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [160]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [678]),
    .S(_12113_),
    .Z(_12162_));
 AND2_X2 _38349_ (.A1(_12162_),
    .A2(_12080_),
    .ZN(_12163_));
 NAND2_X1 _38350_ (.A1(_12069_),
    .A2(_12163_),
    .ZN(_12164_));
 MUX2_X1 _38351_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [224]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [742]),
    .S(_12145_),
    .Z(_12165_));
 AND2_X1 _38352_ (.A1(_12165_),
    .A2(_12071_),
    .ZN(_12166_));
 OAI21_X1 _38353_ (.A(_12166_),
    .B1(_12125_),
    .B2(_12126_),
    .ZN(_12167_));
 AOI21_X1 _38354_ (.A(_11927_),
    .B1(_12164_),
    .B2(_12167_),
    .ZN(_12168_));
 OR2_X4 _38355_ (.A1(_12161_),
    .A2(_12168_),
    .ZN(_12169_));
 MUX2_X2 _38356_ (.A(_12154_),
    .B(_12169_),
    .S(_11769_),
    .Z(\icache.data_mem_data_li [26]));
 MUX2_X2 _38357_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [289]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [807]),
    .S(_12113_),
    .Z(_12170_));
 AND2_X1 _38358_ (.A1(_12170_),
    .A2(_12150_),
    .ZN(_12171_));
 NAND2_X1 _38359_ (.A1(_12137_),
    .A2(_12171_),
    .ZN(_12172_));
 MUX2_X2 _38360_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [353]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [871]),
    .S(_12113_),
    .Z(_12173_));
 AND2_X1 _38361_ (.A1(_12173_),
    .A2(_12150_),
    .ZN(_12174_));
 BUF_X4 _38362_ (.A(_11680_),
    .Z(_12175_));
 BUF_X4 _38363_ (.A(_11682_),
    .Z(_12176_));
 OAI21_X1 _38364_ (.A(_12174_),
    .B1(_12175_),
    .B2(_12176_),
    .ZN(_12177_));
 AOI21_X1 _38365_ (.A(_12003_),
    .B1(_12172_),
    .B2(_12177_),
    .ZN(_12178_));
 MUX2_X2 _38366_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [417]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [935]),
    .S(_12113_),
    .Z(_12179_));
 AND2_X1 _38367_ (.A1(_12179_),
    .A2(_12150_),
    .ZN(_12180_));
 NAND2_X1 _38368_ (.A1(_12137_),
    .A2(_12180_),
    .ZN(_12181_));
 MUX2_X1 _38369_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [481]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [999]),
    .S(_12113_),
    .Z(_12182_));
 AND2_X1 _38370_ (.A1(_12182_),
    .A2(_12150_),
    .ZN(_12183_));
 OAI21_X1 _38371_ (.A(_12183_),
    .B1(_12175_),
    .B2(_12176_),
    .ZN(_12184_));
 AOI21_X1 _38372_ (.A(_12044_),
    .B1(_12181_),
    .B2(_12184_),
    .ZN(_12185_));
 OR2_X4 _38373_ (.A1(_12178_),
    .A2(_12185_),
    .ZN(_12186_));
 MUX2_X1 _38374_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [33]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [551]),
    .S(_11919_),
    .Z(_12187_));
 AND2_X4 _38375_ (.A1(_12187_),
    .A2(_12120_),
    .ZN(_12188_));
 NAND2_X1 _38376_ (.A1(_12069_),
    .A2(_12188_),
    .ZN(_12189_));
 MUX2_X1 _38377_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [97]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [615]),
    .S(_12145_),
    .Z(_12190_));
 AND2_X2 _38378_ (.A1(_12190_),
    .A2(_12071_),
    .ZN(_12191_));
 OAI21_X1 _38379_ (.A(_12191_),
    .B1(_12125_),
    .B2(_12126_),
    .ZN(_12192_));
 AOI21_X1 _38380_ (.A(_11886_),
    .B1(_12189_),
    .B2(_12192_),
    .ZN(_12193_));
 MUX2_X1 _38381_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [161]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [679]),
    .S(_12145_),
    .Z(_12194_));
 AND2_X4 _38382_ (.A1(_12194_),
    .A2(_12071_),
    .ZN(_12195_));
 NAND2_X1 _38383_ (.A1(_12069_),
    .A2(_12195_),
    .ZN(_12196_));
 MUX2_X2 _38384_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [225]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [743]),
    .S(_12145_),
    .Z(_12197_));
 BUF_X2 _38385_ (.A(_11293_),
    .Z(_12198_));
 AND2_X1 _38386_ (.A1(_12197_),
    .A2(_12198_),
    .ZN(_12199_));
 OAI21_X1 _38387_ (.A(_12199_),
    .B1(_12125_),
    .B2(_12126_),
    .ZN(_12200_));
 AOI21_X1 _38388_ (.A(_11927_),
    .B1(_12196_),
    .B2(_12200_),
    .ZN(_12201_));
 OR2_X4 _38389_ (.A1(_12193_),
    .A2(_12201_),
    .ZN(_12202_));
 BUF_X8 _38390_ (.A(_08495_),
    .Z(_12203_));
 MUX2_X2 _38391_ (.A(_12186_),
    .B(_12202_),
    .S(_12203_),
    .Z(\icache.data_mem_data_li [27]));
 MUX2_X1 _38392_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [290]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [808]),
    .S(_12113_),
    .Z(_12204_));
 AND2_X1 _38393_ (.A1(_12204_),
    .A2(_12150_),
    .ZN(_12205_));
 NAND2_X1 _38394_ (.A1(_12137_),
    .A2(_12205_),
    .ZN(_12206_));
 BUF_X8 _38395_ (.A(_11643_),
    .Z(_12207_));
 MUX2_X2 _38396_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [354]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [872]),
    .S(_12207_),
    .Z(_12208_));
 AND2_X1 _38397_ (.A1(_12208_),
    .A2(_12150_),
    .ZN(_12209_));
 OAI21_X1 _38398_ (.A(_12209_),
    .B1(_12175_),
    .B2(_12176_),
    .ZN(_12210_));
 AOI21_X1 _38399_ (.A(_12003_),
    .B1(_12206_),
    .B2(_12210_),
    .ZN(_12211_));
 MUX2_X1 _38400_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [418]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [936]),
    .S(_12207_),
    .Z(_12212_));
 AND2_X1 _38401_ (.A1(_12212_),
    .A2(_12150_),
    .ZN(_12213_));
 NAND2_X1 _38402_ (.A1(_12137_),
    .A2(_12213_),
    .ZN(_12214_));
 MUX2_X1 _38403_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [482]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1000]),
    .S(_12207_),
    .Z(_12215_));
 AND2_X1 _38404_ (.A1(_12215_),
    .A2(_12150_),
    .ZN(_12216_));
 OAI21_X1 _38405_ (.A(_12216_),
    .B1(_12175_),
    .B2(_12176_),
    .ZN(_12217_));
 AOI21_X1 _38406_ (.A(_12044_),
    .B1(_12214_),
    .B2(_12217_),
    .ZN(_12218_));
 OR2_X4 _38407_ (.A1(_12211_),
    .A2(_12218_),
    .ZN(_12219_));
 BUF_X8 _38408_ (.A(_11546_),
    .Z(_12220_));
 MUX2_X1 _38409_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [34]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [552]),
    .S(_11919_),
    .Z(_12221_));
 AND2_X4 _38410_ (.A1(_12221_),
    .A2(_12120_),
    .ZN(_12222_));
 NAND2_X1 _38411_ (.A1(_12069_),
    .A2(_12222_),
    .ZN(_12223_));
 MUX2_X2 _38412_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [98]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [616]),
    .S(_12145_),
    .Z(_12224_));
 AND2_X1 _38413_ (.A1(_12224_),
    .A2(_12198_),
    .ZN(_12225_));
 OAI21_X1 _38414_ (.A(_12225_),
    .B1(_12125_),
    .B2(_12126_),
    .ZN(_12226_));
 AOI21_X1 _38415_ (.A(_12220_),
    .B1(_12223_),
    .B2(_12226_),
    .ZN(_12227_));
 MUX2_X2 _38416_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [162]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [680]),
    .S(_12145_),
    .Z(_12228_));
 AND2_X2 _38417_ (.A1(_12228_),
    .A2(_12198_),
    .ZN(_12229_));
 NAND2_X1 _38418_ (.A1(_12069_),
    .A2(_12229_),
    .ZN(_12230_));
 MUX2_X2 _38419_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [226]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [744]),
    .S(_12145_),
    .Z(_12231_));
 AND2_X1 _38420_ (.A1(_12231_),
    .A2(_12198_),
    .ZN(_12232_));
 OAI21_X1 _38421_ (.A(_12232_),
    .B1(_12125_),
    .B2(_12126_),
    .ZN(_12233_));
 AOI21_X1 _38422_ (.A(_11927_),
    .B1(_12230_),
    .B2(_12233_),
    .ZN(_12234_));
 OR2_X4 _38423_ (.A1(_12227_),
    .A2(_12234_),
    .ZN(_12235_));
 MUX2_X2 _38424_ (.A(_12219_),
    .B(_12235_),
    .S(_12203_),
    .Z(\icache.data_mem_data_li [28]));
 BUF_X4 _38425_ (.A(_11413_),
    .Z(_12236_));
 BUF_X8 _38426_ (.A(_11835_),
    .Z(_12237_));
 MUX2_X1 _38427_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [291]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [809]),
    .S(_12237_),
    .Z(_12238_));
 AND2_X1 _38428_ (.A1(_12238_),
    .A2(_12198_),
    .ZN(_12239_));
 NAND2_X1 _38429_ (.A1(_12236_),
    .A2(_12239_),
    .ZN(_12240_));
 MUX2_X2 _38430_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [355]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [873]),
    .S(_12237_),
    .Z(_12241_));
 AND2_X1 _38431_ (.A1(_12241_),
    .A2(_12198_),
    .ZN(_12242_));
 OAI21_X1 _38432_ (.A(_12242_),
    .B1(_12125_),
    .B2(_12126_),
    .ZN(_12243_));
 AOI21_X1 _38433_ (.A(_12003_),
    .B1(_12240_),
    .B2(_12243_),
    .ZN(_12244_));
 MUX2_X1 _38434_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [419]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [937]),
    .S(_12207_),
    .Z(_12245_));
 BUF_X2 _38435_ (.A(_12079_),
    .Z(_12246_));
 AND2_X2 _38436_ (.A1(_12245_),
    .A2(_12246_),
    .ZN(_12247_));
 NAND2_X1 _38437_ (.A1(_12137_),
    .A2(_12247_),
    .ZN(_12248_));
 MUX2_X1 _38438_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [483]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1001]),
    .S(_12207_),
    .Z(_12249_));
 AND2_X1 _38439_ (.A1(_12249_),
    .A2(_12246_),
    .ZN(_12250_));
 OAI21_X2 _38440_ (.A(_12250_),
    .B1(_12175_),
    .B2(_12176_),
    .ZN(_12251_));
 AOI21_X1 _38441_ (.A(_12044_),
    .B1(_12248_),
    .B2(_12251_),
    .ZN(_12252_));
 OR2_X4 _38442_ (.A1(_12244_),
    .A2(_12252_),
    .ZN(_12253_));
 MUX2_X1 _38443_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [35]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [553]),
    .S(_11448_),
    .Z(_12254_));
 AND2_X4 _38444_ (.A1(_12254_),
    .A2(_11721_),
    .ZN(_12255_));
 NAND2_X1 _38445_ (.A1(_12137_),
    .A2(_12255_),
    .ZN(_12256_));
 MUX2_X1 _38446_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [99]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [617]),
    .S(_12207_),
    .Z(_12257_));
 AND2_X2 _38447_ (.A1(_12257_),
    .A2(_12150_),
    .ZN(_12258_));
 OAI21_X1 _38448_ (.A(_12258_),
    .B1(_12175_),
    .B2(_12176_),
    .ZN(_12259_));
 AOI21_X1 _38449_ (.A(_12220_),
    .B1(_12256_),
    .B2(_12259_),
    .ZN(_12260_));
 BUF_X8 _38450_ (.A(_08493_),
    .Z(_12261_));
 MUX2_X2 _38451_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [163]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [681]),
    .S(_12145_),
    .Z(_12262_));
 AND2_X2 _38452_ (.A1(_12262_),
    .A2(_12198_),
    .ZN(_12263_));
 NAND2_X1 _38453_ (.A1(_12236_),
    .A2(_12263_),
    .ZN(_12264_));
 MUX2_X2 _38454_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [227]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [745]),
    .S(_12145_),
    .Z(_12265_));
 AND2_X1 _38455_ (.A1(_12265_),
    .A2(_12198_),
    .ZN(_12266_));
 OAI21_X2 _38456_ (.A(_12266_),
    .B1(_12125_),
    .B2(_12126_),
    .ZN(_12267_));
 AOI21_X1 _38457_ (.A(_12261_),
    .B1(_12264_),
    .B2(_12267_),
    .ZN(_12268_));
 OR2_X4 _38458_ (.A1(_12260_),
    .A2(_12268_),
    .ZN(_12269_));
 MUX2_X2 _38459_ (.A(_12253_),
    .B(_12269_),
    .S(_12203_),
    .Z(\icache.data_mem_data_li [29]));
 MUX2_X1 _38460_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [292]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [810]),
    .S(_12207_),
    .Z(_12270_));
 AND2_X1 _38461_ (.A1(_12270_),
    .A2(_12246_),
    .ZN(_12271_));
 NAND2_X1 _38462_ (.A1(_12137_),
    .A2(_12271_),
    .ZN(_12272_));
 MUX2_X2 _38463_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [356]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [874]),
    .S(_12207_),
    .Z(_12273_));
 AND2_X1 _38464_ (.A1(_12273_),
    .A2(_12246_),
    .ZN(_12274_));
 OAI21_X1 _38465_ (.A(_12274_),
    .B1(_12175_),
    .B2(_12176_),
    .ZN(_12275_));
 AOI21_X1 _38466_ (.A(_12003_),
    .B1(_12272_),
    .B2(_12275_),
    .ZN(_12276_));
 MUX2_X1 _38467_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [420]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [938]),
    .S(_12207_),
    .Z(_12277_));
 AND2_X1 _38468_ (.A1(_12277_),
    .A2(_12246_),
    .ZN(_12278_));
 NAND2_X1 _38469_ (.A1(_12137_),
    .A2(_12278_),
    .ZN(_12279_));
 MUX2_X1 _38470_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [484]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1002]),
    .S(_12207_),
    .Z(_12280_));
 AND2_X1 _38471_ (.A1(_12280_),
    .A2(_12246_),
    .ZN(_12281_));
 OAI21_X1 _38472_ (.A(_12281_),
    .B1(_12175_),
    .B2(_12176_),
    .ZN(_12282_));
 AOI21_X1 _38473_ (.A(_12044_),
    .B1(_12279_),
    .B2(_12282_),
    .ZN(_12283_));
 OR2_X4 _38474_ (.A1(_12276_),
    .A2(_12283_),
    .ZN(_12284_));
 MUX2_X1 _38475_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [36]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [554]),
    .S(_11919_),
    .Z(_12285_));
 AND2_X4 _38476_ (.A1(_12285_),
    .A2(_12120_),
    .ZN(_12286_));
 NAND2_X1 _38477_ (.A1(_12236_),
    .A2(_12286_),
    .ZN(_12287_));
 MUX2_X2 _38478_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [100]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [618]),
    .S(_12237_),
    .Z(_12288_));
 AND2_X1 _38479_ (.A1(_12288_),
    .A2(_12198_),
    .ZN(_12289_));
 BUF_X4 _38480_ (.A(_11251_),
    .Z(_12290_));
 BUF_X4 _38481_ (.A(_11253_),
    .Z(_12291_));
 OAI21_X1 _38482_ (.A(_12289_),
    .B1(_12290_),
    .B2(_12291_),
    .ZN(_12292_));
 AOI21_X1 _38483_ (.A(_12220_),
    .B1(_12287_),
    .B2(_12292_),
    .ZN(_12293_));
 MUX2_X2 _38484_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [164]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [682]),
    .S(_12237_),
    .Z(_12294_));
 AND2_X1 _38485_ (.A1(_12294_),
    .A2(_12198_),
    .ZN(_12295_));
 NAND2_X1 _38486_ (.A1(_12236_),
    .A2(_12295_),
    .ZN(_12296_));
 MUX2_X2 _38487_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [228]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [746]),
    .S(_12237_),
    .Z(_12297_));
 BUF_X16 _38488_ (.A(_08426_),
    .Z(_12298_));
 BUF_X4 _38489_ (.A(_12298_),
    .Z(_12299_));
 AND2_X1 _38490_ (.A1(_12297_),
    .A2(_12299_),
    .ZN(_12300_));
 OAI21_X1 _38491_ (.A(_12300_),
    .B1(_12290_),
    .B2(_12291_),
    .ZN(_12301_));
 AOI21_X1 _38492_ (.A(_12261_),
    .B1(_12296_),
    .B2(_12301_),
    .ZN(_12302_));
 OR2_X4 _38493_ (.A1(_12293_),
    .A2(_12302_),
    .ZN(_12303_));
 MUX2_X2 _38494_ (.A(_12284_),
    .B(_12303_),
    .S(_12203_),
    .Z(\icache.data_mem_data_li [30]));
 BUF_X4 _38495_ (.A(_11301_),
    .Z(_12304_));
 BUF_X16 _38496_ (.A(_08427_),
    .Z(_12305_));
 MUX2_X1 _38497_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [37]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [555]),
    .S(_12305_),
    .Z(_12306_));
 AND2_X4 _38498_ (.A1(_12306_),
    .A2(_11721_),
    .ZN(_12307_));
 NAND2_X1 _38499_ (.A1(_12304_),
    .A2(_12307_),
    .ZN(_12308_));
 BUF_X8 _38500_ (.A(_11643_),
    .Z(_12309_));
 MUX2_X2 _38501_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [101]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [619]),
    .S(_12309_),
    .Z(_12310_));
 AND2_X2 _38502_ (.A1(_12310_),
    .A2(_12246_),
    .ZN(_12311_));
 OAI21_X1 _38503_ (.A(_12311_),
    .B1(_12175_),
    .B2(_12176_),
    .ZN(_12312_));
 AOI21_X1 _38504_ (.A(_12003_),
    .B1(_12308_),
    .B2(_12312_),
    .ZN(_12313_));
 MUX2_X1 _38505_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [165]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [683]),
    .S(_12309_),
    .Z(_12314_));
 AND2_X1 _38506_ (.A1(_12314_),
    .A2(_12246_),
    .ZN(_12315_));
 NAND2_X1 _38507_ (.A1(_12304_),
    .A2(_12315_),
    .ZN(_12316_));
 MUX2_X2 _38508_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [229]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [747]),
    .S(_12309_),
    .Z(_12317_));
 AND2_X1 _38509_ (.A1(_12317_),
    .A2(_12246_),
    .ZN(_12318_));
 OAI21_X1 _38510_ (.A(_12318_),
    .B1(_12175_),
    .B2(_12176_),
    .ZN(_12319_));
 AOI21_X1 _38511_ (.A(_12044_),
    .B1(_12316_),
    .B2(_12319_),
    .ZN(_12320_));
 OR2_X4 _38512_ (.A1(_12313_),
    .A2(_12320_),
    .ZN(_12321_));
 MUX2_X2 _38513_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [293]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [811]),
    .S(_12237_),
    .Z(_12322_));
 AND2_X1 _38514_ (.A1(_12322_),
    .A2(_12299_),
    .ZN(_12323_));
 NAND2_X1 _38515_ (.A1(_12236_),
    .A2(_12323_),
    .ZN(_12324_));
 MUX2_X1 _38516_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [357]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [875]),
    .S(_12237_),
    .Z(_12325_));
 AND2_X1 _38517_ (.A1(_12325_),
    .A2(_12299_),
    .ZN(_12326_));
 OAI21_X1 _38518_ (.A(_12326_),
    .B1(_12290_),
    .B2(_12291_),
    .ZN(_12327_));
 AOI21_X1 _38519_ (.A(_12220_),
    .B1(_12324_),
    .B2(_12327_),
    .ZN(_12328_));
 MUX2_X2 _38520_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [421]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [939]),
    .S(_12237_),
    .Z(_12329_));
 AND2_X1 _38521_ (.A1(_12329_),
    .A2(_12299_),
    .ZN(_12330_));
 NAND2_X1 _38522_ (.A1(_12236_),
    .A2(_12330_),
    .ZN(_12331_));
 MUX2_X2 _38523_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [485]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1003]),
    .S(_12237_),
    .Z(_12332_));
 AND2_X1 _38524_ (.A1(_12332_),
    .A2(_12299_),
    .ZN(_12333_));
 OAI21_X1 _38525_ (.A(_12333_),
    .B1(_12290_),
    .B2(_12291_),
    .ZN(_12334_));
 AOI21_X1 _38526_ (.A(_12261_),
    .B1(_12331_),
    .B2(_12334_),
    .ZN(_12335_));
 OR2_X4 _38527_ (.A1(_12328_),
    .A2(_12335_),
    .ZN(_12336_));
 BUF_X8 _38528_ (.A(_08433_),
    .Z(_12337_));
 MUX2_X2 _38529_ (.A(_12321_),
    .B(_12336_),
    .S(_12337_),
    .Z(\icache.data_mem_data_li [31]));
 BUF_X4 _38530_ (.A(_11665_),
    .Z(_12338_));
 MUX2_X1 _38531_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [38]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [556]),
    .S(_11919_),
    .Z(_12339_));
 AND2_X4 _38532_ (.A1(_12339_),
    .A2(_12120_),
    .ZN(_12340_));
 NAND2_X1 _38533_ (.A1(_12236_),
    .A2(_12340_),
    .ZN(_12341_));
 BUF_X8 _38534_ (.A(_11835_),
    .Z(_12342_));
 MUX2_X2 _38535_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [102]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [620]),
    .S(_12342_),
    .Z(_12343_));
 AND2_X1 _38536_ (.A1(_12343_),
    .A2(_12299_),
    .ZN(_12344_));
 OAI21_X1 _38537_ (.A(_12344_),
    .B1(_12290_),
    .B2(_12291_),
    .ZN(_12345_));
 AOI21_X1 _38538_ (.A(_12338_),
    .B1(_12341_),
    .B2(_12345_),
    .ZN(_12346_));
 MUX2_X2 _38539_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [166]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [684]),
    .S(_12342_),
    .Z(_12347_));
 AND2_X1 _38540_ (.A1(_12347_),
    .A2(_12299_),
    .ZN(_12348_));
 NAND2_X1 _38541_ (.A1(_12304_),
    .A2(_12348_),
    .ZN(_12349_));
 MUX2_X1 _38542_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [230]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [748]),
    .S(_12309_),
    .Z(_12350_));
 BUF_X2 _38543_ (.A(_12079_),
    .Z(_12351_));
 AND2_X1 _38544_ (.A1(_12350_),
    .A2(_12351_),
    .ZN(_12352_));
 BUF_X4 _38545_ (.A(_11680_),
    .Z(_12353_));
 BUF_X4 _38546_ (.A(_11682_),
    .Z(_12354_));
 OAI21_X2 _38547_ (.A(_12352_),
    .B1(_12353_),
    .B2(_12354_),
    .ZN(_12355_));
 AOI21_X1 _38548_ (.A(_12044_),
    .B1(_12349_),
    .B2(_12355_),
    .ZN(_12356_));
 OR2_X4 _38549_ (.A1(_12346_),
    .A2(_12356_),
    .ZN(_12357_));
 MUX2_X2 _38550_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [294]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [812]),
    .S(_12309_),
    .Z(_12358_));
 AND2_X1 _38551_ (.A1(_12358_),
    .A2(_12246_),
    .ZN(_12359_));
 NAND2_X1 _38552_ (.A1(_12304_),
    .A2(_12359_),
    .ZN(_12360_));
 MUX2_X1 _38553_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [358]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [876]),
    .S(_12309_),
    .Z(_12361_));
 AND2_X1 _38554_ (.A1(_12361_),
    .A2(_12351_),
    .ZN(_12362_));
 OAI21_X2 _38555_ (.A(_12362_),
    .B1(_12353_),
    .B2(_12354_),
    .ZN(_12363_));
 AOI21_X1 _38556_ (.A(_12220_),
    .B1(_12360_),
    .B2(_12363_),
    .ZN(_12364_));
 MUX2_X1 _38557_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [422]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [940]),
    .S(_12309_),
    .Z(_12365_));
 AND2_X1 _38558_ (.A1(_12365_),
    .A2(_12351_),
    .ZN(_12366_));
 NAND2_X1 _38559_ (.A1(_12236_),
    .A2(_12366_),
    .ZN(_12367_));
 MUX2_X1 _38560_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [486]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1004]),
    .S(_12237_),
    .Z(_12368_));
 AND2_X1 _38561_ (.A1(_12368_),
    .A2(_12299_),
    .ZN(_12369_));
 OAI21_X1 _38562_ (.A(_12369_),
    .B1(_12290_),
    .B2(_12291_),
    .ZN(_12370_));
 AOI21_X1 _38563_ (.A(_12261_),
    .B1(_12367_),
    .B2(_12370_),
    .ZN(_12371_));
 OR2_X4 _38564_ (.A1(_12364_),
    .A2(_12371_),
    .ZN(_12372_));
 MUX2_X2 _38565_ (.A(_12357_),
    .B(_12372_),
    .S(_12337_),
    .Z(\icache.data_mem_data_li [32]));
 MUX2_X2 _38566_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [295]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [813]),
    .S(_12342_),
    .Z(_12373_));
 BUF_X4 _38567_ (.A(_12298_),
    .Z(_12374_));
 AND2_X2 _38568_ (.A1(_12373_),
    .A2(_12374_),
    .ZN(_12375_));
 NAND2_X1 _38569_ (.A1(_12236_),
    .A2(_12375_),
    .ZN(_12376_));
 MUX2_X1 _38570_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [359]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [877]),
    .S(_12342_),
    .Z(_12377_));
 AND2_X2 _38571_ (.A1(_12377_),
    .A2(_12374_),
    .ZN(_12378_));
 OAI21_X1 _38572_ (.A(_12378_),
    .B1(_12290_),
    .B2(_12291_),
    .ZN(_12379_));
 AOI21_X1 _38573_ (.A(_12338_),
    .B1(_12376_),
    .B2(_12379_),
    .ZN(_12380_));
 BUF_X4 _38574_ (.A(_11709_),
    .Z(_12381_));
 MUX2_X1 _38575_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [423]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [941]),
    .S(_12309_),
    .Z(_12382_));
 AND2_X1 _38576_ (.A1(_12382_),
    .A2(_12351_),
    .ZN(_12383_));
 NAND2_X1 _38577_ (.A1(_12304_),
    .A2(_12383_),
    .ZN(_12384_));
 MUX2_X2 _38578_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [487]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1005]),
    .S(_12309_),
    .Z(_12385_));
 AND2_X2 _38579_ (.A1(_12385_),
    .A2(_12351_),
    .ZN(_12386_));
 OAI21_X1 _38580_ (.A(_12386_),
    .B1(_12353_),
    .B2(_12354_),
    .ZN(_12387_));
 AOI21_X1 _38581_ (.A(_12381_),
    .B1(_12384_),
    .B2(_12387_),
    .ZN(_12388_));
 OR2_X4 _38582_ (.A1(_12380_),
    .A2(_12388_),
    .ZN(_12389_));
 MUX2_X2 _38583_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [39]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [557]),
    .S(_12305_),
    .Z(_12390_));
 AND2_X4 _38584_ (.A1(_12390_),
    .A2(_11721_),
    .ZN(_12391_));
 NAND2_X1 _38585_ (.A1(_12304_),
    .A2(_12391_),
    .ZN(_12392_));
 MUX2_X2 _38586_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [103]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [621]),
    .S(_12309_),
    .Z(_12393_));
 AND2_X2 _38587_ (.A1(_12393_),
    .A2(_12351_),
    .ZN(_12394_));
 OAI21_X2 _38588_ (.A(_12394_),
    .B1(_12353_),
    .B2(_12354_),
    .ZN(_12395_));
 AOI21_X1 _38589_ (.A(_12220_),
    .B1(_12392_),
    .B2(_12395_),
    .ZN(_12396_));
 MUX2_X2 _38590_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [167]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [685]),
    .S(_12342_),
    .Z(_12397_));
 AND2_X1 _38591_ (.A1(_12397_),
    .A2(_12299_),
    .ZN(_12398_));
 NAND2_X1 _38592_ (.A1(_12236_),
    .A2(_12398_),
    .ZN(_12399_));
 MUX2_X2 _38593_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [231]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [749]),
    .S(_12342_),
    .Z(_12400_));
 AND2_X1 _38594_ (.A1(_12400_),
    .A2(_12299_),
    .ZN(_12401_));
 OAI21_X1 _38595_ (.A(_12401_),
    .B1(_12290_),
    .B2(_12291_),
    .ZN(_12402_));
 AOI21_X1 _38596_ (.A(_12261_),
    .B1(_12399_),
    .B2(_12402_),
    .ZN(_12403_));
 OR2_X4 _38597_ (.A1(_12396_),
    .A2(_12403_),
    .ZN(_12404_));
 MUX2_X2 _38598_ (.A(_12389_),
    .B(_12404_),
    .S(_12203_),
    .Z(\icache.data_mem_data_li [33]));
 BUF_X8 _38599_ (.A(_11643_),
    .Z(_12405_));
 MUX2_X2 _38600_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [296]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [814]),
    .S(_12405_),
    .Z(_12406_));
 AND2_X1 _38601_ (.A1(_12406_),
    .A2(_12351_),
    .ZN(_12407_));
 NAND2_X1 _38602_ (.A1(_12304_),
    .A2(_12407_),
    .ZN(_12408_));
 MUX2_X1 _38603_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [360]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [878]),
    .S(_12405_),
    .Z(_12409_));
 AND2_X1 _38604_ (.A1(_12409_),
    .A2(_12351_),
    .ZN(_12410_));
 OAI21_X1 _38605_ (.A(_12410_),
    .B1(_12353_),
    .B2(_12354_),
    .ZN(_12411_));
 AOI21_X1 _38606_ (.A(_12338_),
    .B1(_12408_),
    .B2(_12411_),
    .ZN(_12412_));
 MUX2_X2 _38607_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [424]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [942]),
    .S(_12405_),
    .Z(_12413_));
 AND2_X1 _38608_ (.A1(_12413_),
    .A2(_12351_),
    .ZN(_12414_));
 NAND2_X1 _38609_ (.A1(_12304_),
    .A2(_12414_),
    .ZN(_12415_));
 MUX2_X1 _38610_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [488]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1006]),
    .S(_12405_),
    .Z(_12416_));
 AND2_X1 _38611_ (.A1(_12416_),
    .A2(_12351_),
    .ZN(_12417_));
 OAI21_X1 _38612_ (.A(_12417_),
    .B1(_12353_),
    .B2(_12354_),
    .ZN(_12418_));
 AOI21_X1 _38613_ (.A(_12381_),
    .B1(_12415_),
    .B2(_12418_),
    .ZN(_12419_));
 OR2_X4 _38614_ (.A1(_12412_),
    .A2(_12419_),
    .ZN(_12420_));
 BUF_X16 _38615_ (.A(_08489_),
    .Z(_12421_));
 BUF_X4 _38616_ (.A(_12421_),
    .Z(_12422_));
 BUF_X8 _38617_ (.A(_08427_),
    .Z(_12423_));
 MUX2_X1 _38618_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [40]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [558]),
    .S(_12423_),
    .Z(_12424_));
 AND2_X4 _38619_ (.A1(_12424_),
    .A2(_12120_),
    .ZN(_12425_));
 NAND2_X1 _38620_ (.A1(_12422_),
    .A2(_12425_),
    .ZN(_12426_));
 MUX2_X2 _38621_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [104]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [622]),
    .S(_12342_),
    .Z(_12427_));
 AND2_X2 _38622_ (.A1(_12427_),
    .A2(_12374_),
    .ZN(_12428_));
 OAI21_X1 _38623_ (.A(_12428_),
    .B1(_12290_),
    .B2(_12291_),
    .ZN(_12429_));
 AOI21_X1 _38624_ (.A(_12220_),
    .B1(_12426_),
    .B2(_12429_),
    .ZN(_12430_));
 MUX2_X1 _38625_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [168]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [686]),
    .S(_12342_),
    .Z(_12431_));
 AND2_X2 _38626_ (.A1(_12431_),
    .A2(_12374_),
    .ZN(_12432_));
 NAND2_X1 _38627_ (.A1(_12422_),
    .A2(_12432_),
    .ZN(_12433_));
 MUX2_X1 _38628_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [232]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [750]),
    .S(_12342_),
    .Z(_12434_));
 AND2_X2 _38629_ (.A1(_12434_),
    .A2(_12374_),
    .ZN(_12435_));
 OAI21_X1 _38630_ (.A(_12435_),
    .B1(_12290_),
    .B2(_12291_),
    .ZN(_12436_));
 AOI21_X1 _38631_ (.A(_12261_),
    .B1(_12433_),
    .B2(_12436_),
    .ZN(_12437_));
 OR2_X4 _38632_ (.A1(_12430_),
    .A2(_12437_),
    .ZN(_12438_));
 MUX2_X2 _38633_ (.A(_12420_),
    .B(_12438_),
    .S(_12203_),
    .Z(\icache.data_mem_data_li [34]));
 MUX2_X2 _38634_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [297]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [815]),
    .S(_12405_),
    .Z(_12439_));
 BUF_X2 _38635_ (.A(_12079_),
    .Z(_12440_));
 AND2_X1 _38636_ (.A1(_12439_),
    .A2(_12440_),
    .ZN(_12441_));
 NAND2_X1 _38637_ (.A1(_12304_),
    .A2(_12441_),
    .ZN(_12442_));
 MUX2_X2 _38638_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [361]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [879]),
    .S(_12405_),
    .Z(_12443_));
 AND2_X1 _38639_ (.A1(_12443_),
    .A2(_12440_),
    .ZN(_12444_));
 OAI21_X1 _38640_ (.A(_12444_),
    .B1(_12353_),
    .B2(_12354_),
    .ZN(_12445_));
 AOI21_X1 _38641_ (.A(_12338_),
    .B1(_12442_),
    .B2(_12445_),
    .ZN(_12446_));
 MUX2_X1 _38642_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [425]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [943]),
    .S(_12405_),
    .Z(_12447_));
 AND2_X1 _38643_ (.A1(_12447_),
    .A2(_12440_),
    .ZN(_12448_));
 NAND2_X1 _38644_ (.A1(_12304_),
    .A2(_12448_),
    .ZN(_12449_));
 MUX2_X2 _38645_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [489]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1007]),
    .S(_12405_),
    .Z(_12450_));
 AND2_X1 _38646_ (.A1(_12450_),
    .A2(_12440_),
    .ZN(_12451_));
 OAI21_X1 _38647_ (.A(_12451_),
    .B1(_12353_),
    .B2(_12354_),
    .ZN(_12452_));
 AOI21_X1 _38648_ (.A(_12381_),
    .B1(_12449_),
    .B2(_12452_),
    .ZN(_12453_));
 OR2_X4 _38649_ (.A1(_12446_),
    .A2(_12453_),
    .ZN(_12454_));
 MUX2_X1 _38650_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [41]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [559]),
    .S(_12423_),
    .Z(_12455_));
 AND2_X4 _38651_ (.A1(_12455_),
    .A2(_12120_),
    .ZN(_12456_));
 NAND2_X1 _38652_ (.A1(_12422_),
    .A2(_12456_),
    .ZN(_12457_));
 MUX2_X1 _38653_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [105]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [623]),
    .S(_12342_),
    .Z(_12458_));
 AND2_X2 _38654_ (.A1(_12458_),
    .A2(_12374_),
    .ZN(_12459_));
 BUF_X4 _38655_ (.A(_11251_),
    .Z(_12460_));
 BUF_X4 _38656_ (.A(_11253_),
    .Z(_12461_));
 OAI21_X1 _38657_ (.A(_12459_),
    .B1(_12460_),
    .B2(_12461_),
    .ZN(_12462_));
 AOI21_X1 _38658_ (.A(_12220_),
    .B1(_12457_),
    .B2(_12462_),
    .ZN(_12463_));
 BUF_X8 _38659_ (.A(_11835_),
    .Z(_12464_));
 MUX2_X1 _38660_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [169]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [687]),
    .S(_12464_),
    .Z(_12465_));
 AND2_X2 _38661_ (.A1(_12465_),
    .A2(_12374_),
    .ZN(_12466_));
 NAND2_X1 _38662_ (.A1(_12422_),
    .A2(_12466_),
    .ZN(_12467_));
 MUX2_X1 _38663_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [233]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [751]),
    .S(_12464_),
    .Z(_12468_));
 AND2_X2 _38664_ (.A1(_12468_),
    .A2(_12374_),
    .ZN(_12469_));
 OAI21_X1 _38665_ (.A(_12469_),
    .B1(_12460_),
    .B2(_12461_),
    .ZN(_12470_));
 AOI21_X1 _38666_ (.A(_12261_),
    .B1(_12467_),
    .B2(_12470_),
    .ZN(_12471_));
 OR2_X4 _38667_ (.A1(_12463_),
    .A2(_12471_),
    .ZN(_12472_));
 MUX2_X2 _38668_ (.A(_12454_),
    .B(_12472_),
    .S(_12203_),
    .Z(\icache.data_mem_data_li [35]));
 BUF_X4 _38669_ (.A(_11301_),
    .Z(_12473_));
 MUX2_X2 _38670_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [298]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [816]),
    .S(_12405_),
    .Z(_12474_));
 AND2_X1 _38671_ (.A1(_12474_),
    .A2(_12440_),
    .ZN(_12475_));
 NAND2_X1 _38672_ (.A1(_12473_),
    .A2(_12475_),
    .ZN(_12476_));
 BUF_X8 _38673_ (.A(_11643_),
    .Z(_12477_));
 MUX2_X1 _38674_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [362]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [880]),
    .S(_12477_),
    .Z(_12478_));
 AND2_X1 _38675_ (.A1(_12478_),
    .A2(_12440_),
    .ZN(_12479_));
 OAI21_X1 _38676_ (.A(_12479_),
    .B1(_12353_),
    .B2(_12354_),
    .ZN(_12480_));
 AOI21_X1 _38677_ (.A(_12338_),
    .B1(_12476_),
    .B2(_12480_),
    .ZN(_12481_));
 MUX2_X1 _38678_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [426]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [944]),
    .S(_12464_),
    .Z(_12482_));
 BUF_X4 _38679_ (.A(_12298_),
    .Z(_12483_));
 AND2_X1 _38680_ (.A1(_12482_),
    .A2(_12483_),
    .ZN(_12484_));
 NAND2_X1 _38681_ (.A1(_12473_),
    .A2(_12484_),
    .ZN(_12485_));
 MUX2_X1 _38682_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [490]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1008]),
    .S(_12477_),
    .Z(_12486_));
 AND2_X1 _38683_ (.A1(_12486_),
    .A2(_12440_),
    .ZN(_12487_));
 OAI21_X1 _38684_ (.A(_12487_),
    .B1(_12353_),
    .B2(_12354_),
    .ZN(_12488_));
 AOI21_X1 _38685_ (.A(_12381_),
    .B1(_12485_),
    .B2(_12488_),
    .ZN(_12489_));
 OR2_X4 _38686_ (.A1(_12481_),
    .A2(_12489_),
    .ZN(_12490_));
 MUX2_X2 _38687_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [42]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [560]),
    .S(_12423_),
    .Z(_12491_));
 AND2_X4 _38688_ (.A1(_12491_),
    .A2(_12120_),
    .ZN(_12492_));
 NAND2_X1 _38689_ (.A1(_12422_),
    .A2(_12492_),
    .ZN(_12493_));
 MUX2_X1 _38690_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [106]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [624]),
    .S(_12464_),
    .Z(_12494_));
 AND2_X2 _38691_ (.A1(_12494_),
    .A2(_12374_),
    .ZN(_12495_));
 OAI21_X1 _38692_ (.A(_12495_),
    .B1(_12460_),
    .B2(_12461_),
    .ZN(_12496_));
 AOI21_X1 _38693_ (.A(_12220_),
    .B1(_12493_),
    .B2(_12496_),
    .ZN(_12497_));
 MUX2_X1 _38694_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [170]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [688]),
    .S(_12405_),
    .Z(_12498_));
 AND2_X1 _38695_ (.A1(_12498_),
    .A2(_12440_),
    .ZN(_12499_));
 NAND2_X1 _38696_ (.A1(_12422_),
    .A2(_12499_),
    .ZN(_12500_));
 MUX2_X2 _38697_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [234]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [752]),
    .S(_12464_),
    .Z(_12501_));
 AND2_X2 _38698_ (.A1(_12501_),
    .A2(_12374_),
    .ZN(_12502_));
 OAI21_X1 _38699_ (.A(_12502_),
    .B1(_12460_),
    .B2(_12461_),
    .ZN(_12503_));
 AOI21_X1 _38700_ (.A(_12261_),
    .B1(_12500_),
    .B2(_12503_),
    .ZN(_12504_));
 OR2_X4 _38701_ (.A1(_12497_),
    .A2(_12504_),
    .ZN(_12505_));
 MUX2_X2 _38702_ (.A(_12490_),
    .B(_12505_),
    .S(_12203_),
    .Z(\icache.data_mem_data_li [36]));
 MUX2_X2 _38703_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [299]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [817]),
    .S(_12464_),
    .Z(_12506_));
 AND2_X1 _38704_ (.A1(_12506_),
    .A2(_12483_),
    .ZN(_12507_));
 NAND2_X1 _38705_ (.A1(_12422_),
    .A2(_12507_),
    .ZN(_12508_));
 MUX2_X2 _38706_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [363]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [881]),
    .S(_12464_),
    .Z(_12509_));
 AND2_X2 _38707_ (.A1(_12509_),
    .A2(_12483_),
    .ZN(_12510_));
 OAI21_X1 _38708_ (.A(_12510_),
    .B1(_12460_),
    .B2(_12461_),
    .ZN(_12511_));
 AOI21_X1 _38709_ (.A(_12338_),
    .B1(_12508_),
    .B2(_12511_),
    .ZN(_12512_));
 MUX2_X2 _38710_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [427]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [945]),
    .S(_12477_),
    .Z(_12513_));
 AND2_X1 _38711_ (.A1(_12513_),
    .A2(_12440_),
    .ZN(_12514_));
 NAND2_X1 _38712_ (.A1(_12473_),
    .A2(_12514_),
    .ZN(_12515_));
 MUX2_X1 _38713_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [491]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1009]),
    .S(_12477_),
    .Z(_12516_));
 BUF_X4 _38714_ (.A(_12079_),
    .Z(_12517_));
 AND2_X1 _38715_ (.A1(_12516_),
    .A2(_12517_),
    .ZN(_12518_));
 BUF_X4 _38716_ (.A(_11680_),
    .Z(_12519_));
 BUF_X4 _38717_ (.A(_11682_),
    .Z(_12520_));
 OAI21_X1 _38718_ (.A(_12518_),
    .B1(_12519_),
    .B2(_12520_),
    .ZN(_12521_));
 AOI21_X1 _38719_ (.A(_12381_),
    .B1(_12515_),
    .B2(_12521_),
    .ZN(_12522_));
 OR2_X4 _38720_ (.A1(_12512_),
    .A2(_12522_),
    .ZN(_12523_));
 MUX2_X2 _38721_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [43]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [561]),
    .S(_12305_),
    .Z(_12524_));
 AND2_X4 _38722_ (.A1(_12524_),
    .A2(_11721_),
    .ZN(_12525_));
 NAND2_X1 _38723_ (.A1(_12473_),
    .A2(_12525_),
    .ZN(_12526_));
 MUX2_X1 _38724_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [107]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [625]),
    .S(_12477_),
    .Z(_12527_));
 AND2_X1 _38725_ (.A1(_12527_),
    .A2(_12440_),
    .ZN(_12528_));
 OAI21_X2 _38726_ (.A(_12528_),
    .B1(_12519_),
    .B2(_12520_),
    .ZN(_12529_));
 AOI21_X1 _38727_ (.A(_12220_),
    .B1(_12526_),
    .B2(_12529_),
    .ZN(_12530_));
 MUX2_X1 _38728_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [171]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [689]),
    .S(_12464_),
    .Z(_12531_));
 AND2_X2 _38729_ (.A1(_12531_),
    .A2(_12483_),
    .ZN(_12532_));
 NAND2_X1 _38730_ (.A1(_12422_),
    .A2(_12532_),
    .ZN(_12533_));
 MUX2_X2 _38731_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [235]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [753]),
    .S(_12464_),
    .Z(_12534_));
 AND2_X2 _38732_ (.A1(_12534_),
    .A2(_12483_),
    .ZN(_12535_));
 OAI21_X1 _38733_ (.A(_12535_),
    .B1(_12460_),
    .B2(_12461_),
    .ZN(_12536_));
 AOI21_X1 _38734_ (.A(_12261_),
    .B1(_12533_),
    .B2(_12536_),
    .ZN(_12537_));
 OR2_X4 _38735_ (.A1(_12530_),
    .A2(_12537_),
    .ZN(_12538_));
 MUX2_X2 _38736_ (.A(_12523_),
    .B(_12538_),
    .S(_12203_),
    .Z(\icache.data_mem_data_li [37]));
 BUF_X8 _38737_ (.A(_11835_),
    .Z(_12539_));
 MUX2_X2 _38738_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [300]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [818]),
    .S(_12539_),
    .Z(_12540_));
 AND2_X2 _38739_ (.A1(_12540_),
    .A2(_12483_),
    .ZN(_12541_));
 NAND2_X1 _38740_ (.A1(_12422_),
    .A2(_12541_),
    .ZN(_12542_));
 MUX2_X2 _38741_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [364]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [882]),
    .S(_12539_),
    .Z(_12543_));
 AND2_X2 _38742_ (.A1(_12543_),
    .A2(_12483_),
    .ZN(_12544_));
 OAI21_X1 _38743_ (.A(_12544_),
    .B1(_12460_),
    .B2(_12461_),
    .ZN(_12545_));
 AOI21_X1 _38744_ (.A(_12338_),
    .B1(_12542_),
    .B2(_12545_),
    .ZN(_12546_));
 MUX2_X2 _38745_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [428]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [946]),
    .S(_12477_),
    .Z(_12547_));
 AND2_X2 _38746_ (.A1(_12547_),
    .A2(_12517_),
    .ZN(_12548_));
 NAND2_X1 _38747_ (.A1(_12473_),
    .A2(_12548_),
    .ZN(_12549_));
 MUX2_X1 _38748_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [492]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1010]),
    .S(_12477_),
    .Z(_12550_));
 AND2_X1 _38749_ (.A1(_12550_),
    .A2(_12517_),
    .ZN(_12551_));
 OAI21_X1 _38750_ (.A(_12551_),
    .B1(_12519_),
    .B2(_12520_),
    .ZN(_12552_));
 AOI21_X1 _38751_ (.A(_12381_),
    .B1(_12549_),
    .B2(_12552_),
    .ZN(_12553_));
 OR2_X4 _38752_ (.A1(_12546_),
    .A2(_12553_),
    .ZN(_12554_));
 BUF_X4 _38753_ (.A(_11546_),
    .Z(_12555_));
 MUX2_X1 _38754_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [44]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [562]),
    .S(_12305_),
    .Z(_12556_));
 AND2_X4 _38755_ (.A1(_12556_),
    .A2(_11721_),
    .ZN(_12557_));
 NAND2_X1 _38756_ (.A1(_12473_),
    .A2(_12557_),
    .ZN(_12558_));
 MUX2_X2 _38757_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [108]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [626]),
    .S(_12477_),
    .Z(_12559_));
 AND2_X2 _38758_ (.A1(_12559_),
    .A2(_12517_),
    .ZN(_12560_));
 OAI21_X2 _38759_ (.A(_12560_),
    .B1(_12519_),
    .B2(_12520_),
    .ZN(_12561_));
 AOI21_X1 _38760_ (.A(_12555_),
    .B1(_12558_),
    .B2(_12561_),
    .ZN(_12562_));
 MUX2_X1 _38761_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [172]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [690]),
    .S(_12464_),
    .Z(_12563_));
 AND2_X2 _38762_ (.A1(_12563_),
    .A2(_12483_),
    .ZN(_12564_));
 NAND2_X1 _38763_ (.A1(_12422_),
    .A2(_12564_),
    .ZN(_12565_));
 MUX2_X1 _38764_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [236]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [754]),
    .S(_12539_),
    .Z(_12566_));
 AND2_X2 _38765_ (.A1(_12566_),
    .A2(_12483_),
    .ZN(_12567_));
 OAI21_X1 _38766_ (.A(_12567_),
    .B1(_12460_),
    .B2(_12461_),
    .ZN(_12568_));
 AOI21_X1 _38767_ (.A(_12261_),
    .B1(_12565_),
    .B2(_12568_),
    .ZN(_12569_));
 OR2_X4 _38768_ (.A1(_12562_),
    .A2(_12569_),
    .ZN(_12570_));
 MUX2_X2 _38769_ (.A(_12554_),
    .B(_12570_),
    .S(_12203_),
    .Z(\icache.data_mem_data_li [38]));
 BUF_X4 _38770_ (.A(_12421_),
    .Z(_12571_));
 MUX2_X2 _38771_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [45]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [563]),
    .S(_12423_),
    .Z(_12572_));
 AND2_X4 _38772_ (.A1(_12572_),
    .A2(_12120_),
    .ZN(_12573_));
 NAND2_X1 _38773_ (.A1(_12571_),
    .A2(_12573_),
    .ZN(_12574_));
 MUX2_X1 _38774_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [109]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [627]),
    .S(_12539_),
    .Z(_12575_));
 BUF_X2 _38775_ (.A(_12298_),
    .Z(_12576_));
 AND2_X2 _38776_ (.A1(_12575_),
    .A2(_12576_),
    .ZN(_12577_));
 OAI21_X1 _38777_ (.A(_12577_),
    .B1(_12460_),
    .B2(_12461_),
    .ZN(_12578_));
 AOI21_X1 _38778_ (.A(_12338_),
    .B1(_12574_),
    .B2(_12578_),
    .ZN(_12579_));
 MUX2_X2 _38779_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [173]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [691]),
    .S(_12539_),
    .Z(_12580_));
 AND2_X2 _38780_ (.A1(_12580_),
    .A2(_12576_),
    .ZN(_12581_));
 NAND2_X1 _38781_ (.A1(_12473_),
    .A2(_12581_),
    .ZN(_12582_));
 BUF_X8 _38782_ (.A(_11241_),
    .Z(_12583_));
 MUX2_X1 _38783_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [237]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [755]),
    .S(_12583_),
    .Z(_12584_));
 AND2_X2 _38784_ (.A1(_12584_),
    .A2(_12517_),
    .ZN(_12585_));
 OAI21_X1 _38785_ (.A(_12585_),
    .B1(_12519_),
    .B2(_12520_),
    .ZN(_12586_));
 AOI21_X1 _38786_ (.A(_12381_),
    .B1(_12582_),
    .B2(_12586_),
    .ZN(_12587_));
 OR2_X4 _38787_ (.A1(_12579_),
    .A2(_12587_),
    .ZN(_12588_));
 MUX2_X2 _38788_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [301]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [819]),
    .S(_12477_),
    .Z(_12589_));
 AND2_X2 _38789_ (.A1(_12589_),
    .A2(_12517_),
    .ZN(_12590_));
 NAND2_X1 _38790_ (.A1(_12473_),
    .A2(_12590_),
    .ZN(_12591_));
 MUX2_X2 _38791_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [365]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [883]),
    .S(_12477_),
    .Z(_12592_));
 AND2_X2 _38792_ (.A1(_12592_),
    .A2(_12517_),
    .ZN(_12593_));
 OAI21_X2 _38793_ (.A(_12593_),
    .B1(_12519_),
    .B2(_12520_),
    .ZN(_12594_));
 AOI21_X1 _38794_ (.A(_12555_),
    .B1(_12591_),
    .B2(_12594_),
    .ZN(_12595_));
 BUF_X4 _38795_ (.A(_08493_),
    .Z(_12596_));
 MUX2_X2 _38796_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [429]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [947]),
    .S(_12583_),
    .Z(_12597_));
 AND2_X2 _38797_ (.A1(_12597_),
    .A2(_12517_),
    .ZN(_12598_));
 NAND2_X1 _38798_ (.A1(_12571_),
    .A2(_12598_),
    .ZN(_12599_));
 MUX2_X1 _38799_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [493]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1011]),
    .S(_12539_),
    .Z(_12600_));
 AND2_X2 _38800_ (.A1(_12600_),
    .A2(_12483_),
    .ZN(_12601_));
 OAI21_X1 _38801_ (.A(_12601_),
    .B1(_12460_),
    .B2(_12461_),
    .ZN(_12602_));
 AOI21_X1 _38802_ (.A(_12596_),
    .B1(_12599_),
    .B2(_12602_),
    .ZN(_12603_));
 OR2_X4 _38803_ (.A1(_12595_),
    .A2(_12603_),
    .ZN(_12604_));
 MUX2_X2 _38804_ (.A(_12588_),
    .B(_12604_),
    .S(_12337_),
    .Z(\icache.data_mem_data_li [39]));
 MUX2_X2 _38805_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [302]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [820]),
    .S(_12539_),
    .Z(_12605_));
 AND2_X2 _38806_ (.A1(_12605_),
    .A2(_12576_),
    .ZN(_12606_));
 NAND2_X1 _38807_ (.A1(_12571_),
    .A2(_12606_),
    .ZN(_12607_));
 MUX2_X2 _38808_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [366]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [884]),
    .S(_12539_),
    .Z(_12608_));
 AND2_X2 _38809_ (.A1(_12608_),
    .A2(_12576_),
    .ZN(_12609_));
 BUF_X32 _38810_ (.A(_08483_),
    .Z(_12610_));
 BUF_X4 _38811_ (.A(_12610_),
    .Z(_12611_));
 BUF_X32 _38812_ (.A(_08487_),
    .Z(_12612_));
 BUF_X4 _38813_ (.A(_12612_),
    .Z(_12613_));
 OAI21_X1 _38814_ (.A(_12609_),
    .B1(_12611_),
    .B2(_12613_),
    .ZN(_12614_));
 AOI21_X1 _38815_ (.A(_12338_),
    .B1(_12607_),
    .B2(_12614_),
    .ZN(_12615_));
 MUX2_X2 _38816_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [430]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [948]),
    .S(_12539_),
    .Z(_12616_));
 AND2_X2 _38817_ (.A1(_12616_),
    .A2(_12576_),
    .ZN(_12617_));
 NAND2_X1 _38818_ (.A1(_12473_),
    .A2(_12617_),
    .ZN(_12618_));
 MUX2_X1 _38819_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [494]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1012]),
    .S(_12583_),
    .Z(_12619_));
 BUF_X4 _38820_ (.A(_12079_),
    .Z(_12620_));
 AND2_X2 _38821_ (.A1(_12619_),
    .A2(_12620_),
    .ZN(_12621_));
 OAI21_X1 _38822_ (.A(_12621_),
    .B1(_12519_),
    .B2(_12520_),
    .ZN(_12622_));
 AOI21_X1 _38823_ (.A(_12381_),
    .B1(_12618_),
    .B2(_12622_),
    .ZN(_12623_));
 OR2_X4 _38824_ (.A1(_12615_),
    .A2(_12623_),
    .ZN(_12624_));
 MUX2_X2 _38825_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [46]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [564]),
    .S(_12305_),
    .Z(_12625_));
 AND2_X4 _38826_ (.A1(_12625_),
    .A2(_08500_),
    .ZN(_12626_));
 NAND2_X1 _38827_ (.A1(_12473_),
    .A2(_12626_),
    .ZN(_12627_));
 MUX2_X1 _38828_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [110]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [628]),
    .S(_12583_),
    .Z(_12628_));
 AND2_X2 _38829_ (.A1(_12628_),
    .A2(_12517_),
    .ZN(_12629_));
 OAI21_X2 _38830_ (.A(_12629_),
    .B1(_12519_),
    .B2(_12520_),
    .ZN(_12630_));
 AOI21_X1 _38831_ (.A(_12555_),
    .B1(_12627_),
    .B2(_12630_),
    .ZN(_12631_));
 MUX2_X2 _38832_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [174]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [692]),
    .S(_12583_),
    .Z(_12632_));
 AND2_X2 _38833_ (.A1(_12632_),
    .A2(_12517_),
    .ZN(_12633_));
 NAND2_X1 _38834_ (.A1(_12571_),
    .A2(_12633_),
    .ZN(_12634_));
 MUX2_X2 _38835_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [238]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [756]),
    .S(_12539_),
    .Z(_12635_));
 AND2_X2 _38836_ (.A1(_12635_),
    .A2(_12576_),
    .ZN(_12636_));
 OAI21_X1 _38837_ (.A(_12636_),
    .B1(_12611_),
    .B2(_12613_),
    .ZN(_12637_));
 AOI21_X1 _38838_ (.A(_12596_),
    .B1(_12634_),
    .B2(_12637_),
    .ZN(_12638_));
 OR2_X4 _38839_ (.A1(_12631_),
    .A2(_12638_),
    .ZN(_12639_));
 BUF_X32 _38840_ (.A(_08431_),
    .Z(_12640_));
 BUF_X4 _38841_ (.A(_12640_),
    .Z(_12641_));
 MUX2_X2 _38842_ (.A(_12624_),
    .B(_12639_),
    .S(_12641_),
    .Z(\icache.data_mem_data_li [40]));
 MUX2_X1 _38843_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [47]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [565]),
    .S(_12423_),
    .Z(_12642_));
 BUF_X8 _38844_ (.A(_11244_),
    .Z(_12643_));
 AND2_X4 _38845_ (.A1(_12642_),
    .A2(_12643_),
    .ZN(_12644_));
 NAND2_X1 _38846_ (.A1(_12571_),
    .A2(_12644_),
    .ZN(_12645_));
 BUF_X8 _38847_ (.A(_11835_),
    .Z(_12646_));
 MUX2_X1 _38848_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [111]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [629]),
    .S(_12646_),
    .Z(_12647_));
 AND2_X2 _38849_ (.A1(_12647_),
    .A2(_12576_),
    .ZN(_12648_));
 OAI21_X1 _38850_ (.A(_12648_),
    .B1(_12611_),
    .B2(_12613_),
    .ZN(_12649_));
 AOI21_X1 _38851_ (.A(_12338_),
    .B1(_12645_),
    .B2(_12649_),
    .ZN(_12650_));
 BUF_X4 _38852_ (.A(_11301_),
    .Z(_12651_));
 MUX2_X1 _38853_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [175]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [693]),
    .S(_12646_),
    .Z(_12652_));
 AND2_X1 _38854_ (.A1(_12652_),
    .A2(_12576_),
    .ZN(_12653_));
 NAND2_X1 _38855_ (.A1(_12651_),
    .A2(_12653_),
    .ZN(_12654_));
 MUX2_X1 _38856_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [239]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [757]),
    .S(_12583_),
    .Z(_12655_));
 AND2_X2 _38857_ (.A1(_12655_),
    .A2(_12620_),
    .ZN(_12656_));
 OAI21_X1 _38858_ (.A(_12656_),
    .B1(_12519_),
    .B2(_12520_),
    .ZN(_12657_));
 AOI21_X1 _38859_ (.A(_12381_),
    .B1(_12654_),
    .B2(_12657_),
    .ZN(_12658_));
 OR2_X4 _38860_ (.A1(_12650_),
    .A2(_12658_),
    .ZN(_12659_));
 MUX2_X1 _38861_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [303]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [821]),
    .S(_12583_),
    .Z(_12660_));
 AND2_X2 _38862_ (.A1(_12660_),
    .A2(_12620_),
    .ZN(_12661_));
 NAND2_X1 _38863_ (.A1(_12651_),
    .A2(_12661_),
    .ZN(_12662_));
 MUX2_X2 _38864_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [367]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [885]),
    .S(_12583_),
    .Z(_12663_));
 AND2_X2 _38865_ (.A1(_12663_),
    .A2(_12620_),
    .ZN(_12664_));
 OAI21_X1 _38866_ (.A(_12664_),
    .B1(_12519_),
    .B2(_12520_),
    .ZN(_12665_));
 AOI21_X1 _38867_ (.A(_12555_),
    .B1(_12662_),
    .B2(_12665_),
    .ZN(_12666_));
 MUX2_X1 _38868_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [431]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [949]),
    .S(_12583_),
    .Z(_12667_));
 AND2_X2 _38869_ (.A1(_12667_),
    .A2(_12620_),
    .ZN(_12668_));
 NAND2_X1 _38870_ (.A1(_12571_),
    .A2(_12668_),
    .ZN(_12669_));
 MUX2_X1 _38871_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [495]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1013]),
    .S(_12646_),
    .Z(_12670_));
 AND2_X1 _38872_ (.A1(_12670_),
    .A2(_12576_),
    .ZN(_12671_));
 OAI21_X1 _38873_ (.A(_12671_),
    .B1(_12611_),
    .B2(_12613_),
    .ZN(_12672_));
 AOI21_X1 _38874_ (.A(_12596_),
    .B1(_12669_),
    .B2(_12672_),
    .ZN(_12673_));
 OR2_X4 _38875_ (.A1(_12666_),
    .A2(_12673_),
    .ZN(_12674_));
 MUX2_X2 _38876_ (.A(_12659_),
    .B(_12674_),
    .S(_12337_),
    .Z(\icache.data_mem_data_li [41]));
 BUF_X8 _38877_ (.A(_11665_),
    .Z(_12675_));
 MUX2_X1 _38878_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [48]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [566]),
    .S(_12423_),
    .Z(_12676_));
 AND2_X4 _38879_ (.A1(_12676_),
    .A2(_12643_),
    .ZN(_12677_));
 NAND2_X1 _38880_ (.A1(_12651_),
    .A2(_12677_),
    .ZN(_12678_));
 BUF_X8 _38881_ (.A(_11241_),
    .Z(_12679_));
 MUX2_X1 _38882_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [112]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [630]),
    .S(_12679_),
    .Z(_12680_));
 AND2_X2 _38883_ (.A1(_12680_),
    .A2(_12620_),
    .ZN(_12681_));
 BUF_X4 _38884_ (.A(_11680_),
    .Z(_12682_));
 BUF_X4 _38885_ (.A(_11682_),
    .Z(_12683_));
 OAI21_X1 _38886_ (.A(_12681_),
    .B1(_12682_),
    .B2(_12683_),
    .ZN(_12684_));
 AOI21_X1 _38887_ (.A(_12675_),
    .B1(_12678_),
    .B2(_12684_),
    .ZN(_12685_));
 MUX2_X1 _38888_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [176]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [694]),
    .S(_12646_),
    .Z(_12686_));
 BUF_X4 _38889_ (.A(_12298_),
    .Z(_12687_));
 AND2_X1 _38890_ (.A1(_12686_),
    .A2(_12687_),
    .ZN(_12688_));
 NAND2_X1 _38891_ (.A1(_12651_),
    .A2(_12688_),
    .ZN(_12689_));
 MUX2_X1 _38892_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [240]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [758]),
    .S(_12679_),
    .Z(_12690_));
 AND2_X2 _38893_ (.A1(_12690_),
    .A2(_12620_),
    .ZN(_12691_));
 OAI21_X1 _38894_ (.A(_12691_),
    .B1(_12682_),
    .B2(_12683_),
    .ZN(_12692_));
 AOI21_X1 _38895_ (.A(_12381_),
    .B1(_12689_),
    .B2(_12692_),
    .ZN(_12693_));
 OR2_X4 _38896_ (.A1(_12685_),
    .A2(_12693_),
    .ZN(_12694_));
 MUX2_X2 _38897_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [304]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [822]),
    .S(_12583_),
    .Z(_12695_));
 AND2_X2 _38898_ (.A1(_12695_),
    .A2(_12620_),
    .ZN(_12696_));
 NAND2_X1 _38899_ (.A1(_12571_),
    .A2(_12696_),
    .ZN(_12697_));
 MUX2_X2 _38900_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [368]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [886]),
    .S(_12646_),
    .Z(_12698_));
 AND2_X1 _38901_ (.A1(_12698_),
    .A2(_12576_),
    .ZN(_12699_));
 OAI21_X1 _38902_ (.A(_12699_),
    .B1(_12611_),
    .B2(_12613_),
    .ZN(_12700_));
 AOI21_X1 _38903_ (.A(_12555_),
    .B1(_12697_),
    .B2(_12700_),
    .ZN(_12701_));
 MUX2_X1 _38904_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [432]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [950]),
    .S(_12679_),
    .Z(_12702_));
 AND2_X2 _38905_ (.A1(_12702_),
    .A2(_12620_),
    .ZN(_12703_));
 NAND2_X1 _38906_ (.A1(_12571_),
    .A2(_12703_),
    .ZN(_12704_));
 MUX2_X2 _38907_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [496]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1014]),
    .S(_12646_),
    .Z(_12705_));
 AND2_X1 _38908_ (.A1(_12705_),
    .A2(_12687_),
    .ZN(_12706_));
 OAI21_X1 _38909_ (.A(_12706_),
    .B1(_12611_),
    .B2(_12613_),
    .ZN(_12707_));
 AOI21_X1 _38910_ (.A(_12596_),
    .B1(_12704_),
    .B2(_12707_),
    .ZN(_12708_));
 OR2_X4 _38911_ (.A1(_12701_),
    .A2(_12708_),
    .ZN(_12709_));
 MUX2_X2 _38912_ (.A(_12694_),
    .B(_12709_),
    .S(_12337_),
    .Z(\icache.data_mem_data_li [42]));
 MUX2_X1 _38913_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [49]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [567]),
    .S(_12423_),
    .Z(_12710_));
 AND2_X4 _38914_ (.A1(_12710_),
    .A2(_12643_),
    .ZN(_12711_));
 NAND2_X1 _38915_ (.A1(_12571_),
    .A2(_12711_),
    .ZN(_12712_));
 MUX2_X2 _38916_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [113]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [631]),
    .S(_12646_),
    .Z(_12713_));
 AND2_X2 _38917_ (.A1(_12713_),
    .A2(_12687_),
    .ZN(_12714_));
 OAI21_X1 _38918_ (.A(_12714_),
    .B1(_12611_),
    .B2(_12613_),
    .ZN(_12715_));
 AOI21_X1 _38919_ (.A(_12675_),
    .B1(_12712_),
    .B2(_12715_),
    .ZN(_12716_));
 BUF_X8 _38920_ (.A(_11709_),
    .Z(_12717_));
 MUX2_X1 _38921_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [177]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [695]),
    .S(_12646_),
    .Z(_12718_));
 AND2_X1 _38922_ (.A1(_12718_),
    .A2(_12687_),
    .ZN(_12719_));
 NAND2_X1 _38923_ (.A1(_12651_),
    .A2(_12719_),
    .ZN(_12720_));
 MUX2_X1 _38924_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [241]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [759]),
    .S(_12679_),
    .Z(_12721_));
 BUF_X2 _38925_ (.A(_12079_),
    .Z(_12722_));
 AND2_X1 _38926_ (.A1(_12721_),
    .A2(_12722_),
    .ZN(_12723_));
 OAI21_X2 _38927_ (.A(_12723_),
    .B1(_12682_),
    .B2(_12683_),
    .ZN(_12724_));
 AOI21_X1 _38928_ (.A(_12717_),
    .B1(_12720_),
    .B2(_12724_),
    .ZN(_12725_));
 OR2_X4 _38929_ (.A1(_12716_),
    .A2(_12725_),
    .ZN(_12726_));
 MUX2_X1 _38930_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [305]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [823]),
    .S(_12679_),
    .Z(_12727_));
 AND2_X2 _38931_ (.A1(_12727_),
    .A2(_12620_),
    .ZN(_12728_));
 NAND2_X1 _38932_ (.A1(_12651_),
    .A2(_12728_),
    .ZN(_12729_));
 MUX2_X2 _38933_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [369]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [887]),
    .S(_12679_),
    .Z(_12730_));
 AND2_X1 _38934_ (.A1(_12730_),
    .A2(_12722_),
    .ZN(_12731_));
 OAI21_X2 _38935_ (.A(_12731_),
    .B1(_12682_),
    .B2(_12683_),
    .ZN(_12732_));
 AOI21_X1 _38936_ (.A(_12555_),
    .B1(_12729_),
    .B2(_12732_),
    .ZN(_12733_));
 MUX2_X1 _38937_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [433]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [951]),
    .S(_12679_),
    .Z(_12734_));
 AND2_X2 _38938_ (.A1(_12734_),
    .A2(_12722_),
    .ZN(_12735_));
 NAND2_X1 _38939_ (.A1(_12571_),
    .A2(_12735_),
    .ZN(_12736_));
 MUX2_X1 _38940_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [497]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1015]),
    .S(_12646_),
    .Z(_12737_));
 AND2_X2 _38941_ (.A1(_12737_),
    .A2(_12687_),
    .ZN(_12738_));
 OAI21_X1 _38942_ (.A(_12738_),
    .B1(_12611_),
    .B2(_12613_),
    .ZN(_12739_));
 AOI21_X1 _38943_ (.A(_12596_),
    .B1(_12736_),
    .B2(_12739_),
    .ZN(_12740_));
 OR2_X4 _38944_ (.A1(_12733_),
    .A2(_12740_),
    .ZN(_12741_));
 MUX2_X2 _38945_ (.A(_12726_),
    .B(_12741_),
    .S(_12337_),
    .Z(\icache.data_mem_data_li [43]));
 BUF_X4 _38946_ (.A(_12421_),
    .Z(_12742_));
 BUF_X8 _38947_ (.A(_11835_),
    .Z(_12743_));
 MUX2_X2 _38948_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [306]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [824]),
    .S(_12743_),
    .Z(_12744_));
 AND2_X1 _38949_ (.A1(_12744_),
    .A2(_12687_),
    .ZN(_12745_));
 NAND2_X1 _38950_ (.A1(_12742_),
    .A2(_12745_),
    .ZN(_12746_));
 MUX2_X2 _38951_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [370]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [888]),
    .S(_12743_),
    .Z(_12747_));
 AND2_X1 _38952_ (.A1(_12747_),
    .A2(_12687_),
    .ZN(_12748_));
 OAI21_X1 _38953_ (.A(_12748_),
    .B1(_12611_),
    .B2(_12613_),
    .ZN(_12749_));
 AOI21_X1 _38954_ (.A(_12675_),
    .B1(_12746_),
    .B2(_12749_),
    .ZN(_12750_));
 MUX2_X2 _38955_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [434]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [952]),
    .S(_12679_),
    .Z(_12751_));
 AND2_X1 _38956_ (.A1(_12751_),
    .A2(_12722_),
    .ZN(_12752_));
 NAND2_X1 _38957_ (.A1(_12651_),
    .A2(_12752_),
    .ZN(_12753_));
 MUX2_X1 _38958_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [498]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1016]),
    .S(_12679_),
    .Z(_12754_));
 AND2_X1 _38959_ (.A1(_12754_),
    .A2(_12722_),
    .ZN(_12755_));
 OAI21_X1 _38960_ (.A(_12755_),
    .B1(_12682_),
    .B2(_12683_),
    .ZN(_12756_));
 AOI21_X1 _38961_ (.A(_12717_),
    .B1(_12753_),
    .B2(_12756_),
    .ZN(_12757_));
 OR2_X4 _38962_ (.A1(_12750_),
    .A2(_12757_),
    .ZN(_12758_));
 MUX2_X1 _38963_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [50]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [568]),
    .S(_12305_),
    .Z(_12759_));
 AND2_X4 _38964_ (.A1(_12759_),
    .A2(_08500_),
    .ZN(_12760_));
 NAND2_X1 _38965_ (.A1(_12651_),
    .A2(_12760_),
    .ZN(_12761_));
 MUX2_X1 _38966_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [114]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [632]),
    .S(_12679_),
    .Z(_12762_));
 AND2_X1 _38967_ (.A1(_12762_),
    .A2(_12722_),
    .ZN(_12763_));
 OAI21_X2 _38968_ (.A(_12763_),
    .B1(_12682_),
    .B2(_12683_),
    .ZN(_12764_));
 AOI21_X1 _38969_ (.A(_12555_),
    .B1(_12761_),
    .B2(_12764_),
    .ZN(_12765_));
 MUX2_X1 _38970_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [178]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [696]),
    .S(_12646_),
    .Z(_12766_));
 AND2_X2 _38971_ (.A1(_12766_),
    .A2(_12687_),
    .ZN(_12767_));
 NAND2_X1 _38972_ (.A1(_12742_),
    .A2(_12767_),
    .ZN(_12768_));
 MUX2_X2 _38973_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [242]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [760]),
    .S(_12743_),
    .Z(_12769_));
 AND2_X1 _38974_ (.A1(_12769_),
    .A2(_12687_),
    .ZN(_12770_));
 OAI21_X1 _38975_ (.A(_12770_),
    .B1(_12611_),
    .B2(_12613_),
    .ZN(_12771_));
 AOI21_X1 _38976_ (.A(_12596_),
    .B1(_12768_),
    .B2(_12771_),
    .ZN(_12772_));
 OR2_X4 _38977_ (.A1(_12765_),
    .A2(_12772_),
    .ZN(_12773_));
 MUX2_X2 _38978_ (.A(_12758_),
    .B(_12773_),
    .S(_12641_),
    .Z(\icache.data_mem_data_li [44]));
 MUX2_X2 _38979_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [307]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [825]),
    .S(_12743_),
    .Z(_12774_));
 BUF_X4 _38980_ (.A(_12298_),
    .Z(_12775_));
 AND2_X1 _38981_ (.A1(_12774_),
    .A2(_12775_),
    .ZN(_12776_));
 NAND2_X1 _38982_ (.A1(_12742_),
    .A2(_12776_),
    .ZN(_12777_));
 MUX2_X2 _38983_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [371]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [889]),
    .S(_12743_),
    .Z(_12778_));
 AND2_X1 _38984_ (.A1(_12778_),
    .A2(_12775_),
    .ZN(_12779_));
 BUF_X4 _38985_ (.A(_12610_),
    .Z(_12780_));
 BUF_X4 _38986_ (.A(_12612_),
    .Z(_12781_));
 OAI21_X1 _38987_ (.A(_12779_),
    .B1(_12780_),
    .B2(_12781_),
    .ZN(_12782_));
 AOI21_X1 _38988_ (.A(_12675_),
    .B1(_12777_),
    .B2(_12782_),
    .ZN(_12783_));
 BUF_X8 _38989_ (.A(_11241_),
    .Z(_12784_));
 MUX2_X2 _38990_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [435]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [953]),
    .S(_12784_),
    .Z(_12785_));
 AND2_X1 _38991_ (.A1(_12785_),
    .A2(_12722_),
    .ZN(_12786_));
 NAND2_X1 _38992_ (.A1(_12651_),
    .A2(_12786_),
    .ZN(_12787_));
 MUX2_X2 _38993_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [499]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1017]),
    .S(_12784_),
    .Z(_12788_));
 AND2_X1 _38994_ (.A1(_12788_),
    .A2(_12722_),
    .ZN(_12789_));
 OAI21_X1 _38995_ (.A(_12789_),
    .B1(_12682_),
    .B2(_12683_),
    .ZN(_12790_));
 AOI21_X1 _38996_ (.A(_12717_),
    .B1(_12787_),
    .B2(_12790_),
    .ZN(_12791_));
 OR2_X4 _38997_ (.A1(_12783_),
    .A2(_12791_),
    .ZN(_12792_));
 MUX2_X2 _38998_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [51]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [569]),
    .S(_12305_),
    .Z(_12793_));
 AND2_X4 _38999_ (.A1(_12793_),
    .A2(_08500_),
    .ZN(_12794_));
 NAND2_X1 _39000_ (.A1(_12651_),
    .A2(_12794_),
    .ZN(_12795_));
 MUX2_X2 _39001_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [115]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [633]),
    .S(_12784_),
    .Z(_12796_));
 AND2_X1 _39002_ (.A1(_12796_),
    .A2(_12722_),
    .ZN(_12797_));
 OAI21_X2 _39003_ (.A(_12797_),
    .B1(_12682_),
    .B2(_12683_),
    .ZN(_12798_));
 AOI21_X1 _39004_ (.A(_12555_),
    .B1(_12795_),
    .B2(_12798_),
    .ZN(_12799_));
 MUX2_X1 _39005_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [179]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [697]),
    .S(_12743_),
    .Z(_12800_));
 AND2_X1 _39006_ (.A1(_12800_),
    .A2(_12687_),
    .ZN(_12801_));
 NAND2_X1 _39007_ (.A1(_12742_),
    .A2(_12801_),
    .ZN(_12802_));
 MUX2_X2 _39008_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [243]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [761]),
    .S(_12743_),
    .Z(_12803_));
 AND2_X1 _39009_ (.A1(_12803_),
    .A2(_12775_),
    .ZN(_12804_));
 OAI21_X1 _39010_ (.A(_12804_),
    .B1(_12780_),
    .B2(_12781_),
    .ZN(_12805_));
 AOI21_X1 _39011_ (.A(_12596_),
    .B1(_12802_),
    .B2(_12805_),
    .ZN(_12806_));
 OR2_X4 _39012_ (.A1(_12799_),
    .A2(_12806_),
    .ZN(_12807_));
 MUX2_X2 _39013_ (.A(_12792_),
    .B(_12807_),
    .S(_12641_),
    .Z(\icache.data_mem_data_li [45]));
 BUF_X4 _39014_ (.A(_11301_),
    .Z(_12808_));
 MUX2_X1 _39015_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [308]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [826]),
    .S(_12784_),
    .Z(_12809_));
 BUF_X4 _39016_ (.A(_12079_),
    .Z(_12810_));
 AND2_X1 _39017_ (.A1(_12809_),
    .A2(_12810_),
    .ZN(_12811_));
 NAND2_X1 _39018_ (.A1(_12808_),
    .A2(_12811_),
    .ZN(_12812_));
 MUX2_X1 _39019_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [372]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [890]),
    .S(_12784_),
    .Z(_12813_));
 AND2_X2 _39020_ (.A1(_12813_),
    .A2(_12810_),
    .ZN(_12814_));
 OAI21_X1 _39021_ (.A(_12814_),
    .B1(_12682_),
    .B2(_12683_),
    .ZN(_12815_));
 AOI21_X1 _39022_ (.A(_12675_),
    .B1(_12812_),
    .B2(_12815_),
    .ZN(_12816_));
 MUX2_X2 _39023_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [436]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [954]),
    .S(_12743_),
    .Z(_12817_));
 AND2_X1 _39024_ (.A1(_12817_),
    .A2(_12775_),
    .ZN(_12818_));
 NAND2_X1 _39025_ (.A1(_12808_),
    .A2(_12818_),
    .ZN(_12819_));
 MUX2_X2 _39026_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [500]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1018]),
    .S(_12784_),
    .Z(_12820_));
 AND2_X1 _39027_ (.A1(_12820_),
    .A2(_12810_),
    .ZN(_12821_));
 OAI21_X1 _39028_ (.A(_12821_),
    .B1(_12682_),
    .B2(_12683_),
    .ZN(_12822_));
 AOI21_X1 _39029_ (.A(_12717_),
    .B1(_12819_),
    .B2(_12822_),
    .ZN(_12823_));
 OR2_X4 _39030_ (.A1(_12816_),
    .A2(_12823_),
    .ZN(_12824_));
 MUX2_X2 _39031_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [52]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [570]),
    .S(_12423_),
    .Z(_12825_));
 AND2_X4 _39032_ (.A1(_12825_),
    .A2(_12643_),
    .ZN(_12826_));
 NAND2_X1 _39033_ (.A1(_12742_),
    .A2(_12826_),
    .ZN(_12827_));
 MUX2_X2 _39034_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [116]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [634]),
    .S(_12743_),
    .Z(_12828_));
 AND2_X1 _39035_ (.A1(_12828_),
    .A2(_12775_),
    .ZN(_12829_));
 OAI21_X1 _39036_ (.A(_12829_),
    .B1(_12780_),
    .B2(_12781_),
    .ZN(_12830_));
 AOI21_X1 _39037_ (.A(_12555_),
    .B1(_12827_),
    .B2(_12830_),
    .ZN(_12831_));
 MUX2_X1 _39038_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [180]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [698]),
    .S(_12784_),
    .Z(_12832_));
 AND2_X1 _39039_ (.A1(_12832_),
    .A2(_12722_),
    .ZN(_12833_));
 NAND2_X1 _39040_ (.A1(_12742_),
    .A2(_12833_),
    .ZN(_12834_));
 MUX2_X2 _39041_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [244]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [762]),
    .S(_12743_),
    .Z(_12835_));
 AND2_X1 _39042_ (.A1(_12835_),
    .A2(_12775_),
    .ZN(_12836_));
 OAI21_X1 _39043_ (.A(_12836_),
    .B1(_12780_),
    .B2(_12781_),
    .ZN(_12837_));
 AOI21_X1 _39044_ (.A(_12596_),
    .B1(_12834_),
    .B2(_12837_),
    .ZN(_12838_));
 OR2_X4 _39045_ (.A1(_12831_),
    .A2(_12838_),
    .ZN(_12839_));
 MUX2_X2 _39046_ (.A(_12824_),
    .B(_12839_),
    .S(_12641_),
    .Z(\icache.data_mem_data_li [46]));
 BUF_X8 _39047_ (.A(_11263_),
    .Z(_12840_));
 MUX2_X1 _39048_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [309]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [827]),
    .S(_12840_),
    .Z(_12841_));
 AND2_X1 _39049_ (.A1(_12841_),
    .A2(_12775_),
    .ZN(_12842_));
 NAND2_X1 _39050_ (.A1(_12742_),
    .A2(_12842_),
    .ZN(_12843_));
 MUX2_X2 _39051_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [373]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [891]),
    .S(_12840_),
    .Z(_12844_));
 AND2_X1 _39052_ (.A1(_12844_),
    .A2(_12775_),
    .ZN(_12845_));
 OAI21_X1 _39053_ (.A(_12845_),
    .B1(_12780_),
    .B2(_12781_),
    .ZN(_12846_));
 AOI21_X1 _39054_ (.A(_12675_),
    .B1(_12843_),
    .B2(_12846_),
    .ZN(_12847_));
 MUX2_X1 _39055_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [437]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [955]),
    .S(_12840_),
    .Z(_12848_));
 AND2_X1 _39056_ (.A1(_12848_),
    .A2(_12775_),
    .ZN(_12849_));
 NAND2_X1 _39057_ (.A1(_12808_),
    .A2(_12849_),
    .ZN(_12850_));
 MUX2_X2 _39058_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [501]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1019]),
    .S(_12784_),
    .Z(_12851_));
 AND2_X1 _39059_ (.A1(_12851_),
    .A2(_12810_),
    .ZN(_12852_));
 BUF_X4 _39060_ (.A(_11680_),
    .Z(_12853_));
 BUF_X4 _39061_ (.A(_11682_),
    .Z(_12854_));
 OAI21_X1 _39062_ (.A(_12852_),
    .B1(_12853_),
    .B2(_12854_),
    .ZN(_12855_));
 AOI21_X1 _39063_ (.A(_12717_),
    .B1(_12850_),
    .B2(_12855_),
    .ZN(_12856_));
 OR2_X4 _39064_ (.A1(_12847_),
    .A2(_12856_),
    .ZN(_12857_));
 MUX2_X2 _39065_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [53]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [571]),
    .S(_12305_),
    .Z(_12858_));
 AND2_X4 _39066_ (.A1(_12858_),
    .A2(_08500_),
    .ZN(_12859_));
 NAND2_X1 _39067_ (.A1(_12808_),
    .A2(_12859_),
    .ZN(_12860_));
 MUX2_X1 _39068_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [117]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [635]),
    .S(_12784_),
    .Z(_12861_));
 AND2_X1 _39069_ (.A1(_12861_),
    .A2(_12810_),
    .ZN(_12862_));
 OAI21_X1 _39070_ (.A(_12862_),
    .B1(_12853_),
    .B2(_12854_),
    .ZN(_12863_));
 AOI21_X1 _39071_ (.A(_12555_),
    .B1(_12860_),
    .B2(_12863_),
    .ZN(_12864_));
 MUX2_X1 _39072_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [181]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [699]),
    .S(_12784_),
    .Z(_12865_));
 AND2_X1 _39073_ (.A1(_12865_),
    .A2(_12810_),
    .ZN(_12866_));
 NAND2_X1 _39074_ (.A1(_12742_),
    .A2(_12866_),
    .ZN(_12867_));
 MUX2_X2 _39075_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [245]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [763]),
    .S(_12840_),
    .Z(_12868_));
 AND2_X1 _39076_ (.A1(_12868_),
    .A2(_12775_),
    .ZN(_12869_));
 OAI21_X1 _39077_ (.A(_12869_),
    .B1(_12780_),
    .B2(_12781_),
    .ZN(_12870_));
 AOI21_X1 _39078_ (.A(_12596_),
    .B1(_12867_),
    .B2(_12870_),
    .ZN(_12871_));
 OR2_X4 _39079_ (.A1(_12864_),
    .A2(_12871_),
    .ZN(_12872_));
 MUX2_X2 _39080_ (.A(_12857_),
    .B(_12872_),
    .S(_12641_),
    .Z(\icache.data_mem_data_li [47]));
 MUX2_X2 _39081_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [54]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [572]),
    .S(_12423_),
    .Z(_12873_));
 AND2_X4 _39082_ (.A1(_12873_),
    .A2(_12643_),
    .ZN(_12874_));
 NAND2_X1 _39083_ (.A1(_12742_),
    .A2(_12874_),
    .ZN(_12875_));
 MUX2_X2 _39084_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [118]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [636]),
    .S(_12840_),
    .Z(_12876_));
 BUF_X4 _39085_ (.A(_12298_),
    .Z(_12877_));
 AND2_X1 _39086_ (.A1(_12876_),
    .A2(_12877_),
    .ZN(_12878_));
 OAI21_X1 _39087_ (.A(_12878_),
    .B1(_12780_),
    .B2(_12781_),
    .ZN(_12879_));
 AOI21_X1 _39088_ (.A(_12675_),
    .B1(_12875_),
    .B2(_12879_),
    .ZN(_12880_));
 BUF_X8 _39089_ (.A(_11241_),
    .Z(_12881_));
 MUX2_X2 _39090_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [182]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [700]),
    .S(_12881_),
    .Z(_12882_));
 AND2_X2 _39091_ (.A1(_12882_),
    .A2(_12810_),
    .ZN(_12883_));
 NAND2_X1 _39092_ (.A1(_12808_),
    .A2(_12883_),
    .ZN(_12884_));
 MUX2_X2 _39093_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [246]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [764]),
    .S(_12881_),
    .Z(_12885_));
 AND2_X1 _39094_ (.A1(_12885_),
    .A2(_12810_),
    .ZN(_12886_));
 OAI21_X1 _39095_ (.A(_12886_),
    .B1(_12853_),
    .B2(_12854_),
    .ZN(_12887_));
 AOI21_X1 _39096_ (.A(_12717_),
    .B1(_12884_),
    .B2(_12887_),
    .ZN(_12888_));
 OR2_X4 _39097_ (.A1(_12880_),
    .A2(_12888_),
    .ZN(_12889_));
 BUF_X8 _39098_ (.A(_11546_),
    .Z(_12890_));
 MUX2_X2 _39099_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [310]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [828]),
    .S(_12881_),
    .Z(_12891_));
 AND2_X1 _39100_ (.A1(_12891_),
    .A2(_12810_),
    .ZN(_12892_));
 NAND2_X1 _39101_ (.A1(_12808_),
    .A2(_12892_),
    .ZN(_12893_));
 MUX2_X1 _39102_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [374]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [892]),
    .S(_12881_),
    .Z(_12894_));
 AND2_X1 _39103_ (.A1(_12894_),
    .A2(_12810_),
    .ZN(_12895_));
 OAI21_X2 _39104_ (.A(_12895_),
    .B1(_12853_),
    .B2(_12854_),
    .ZN(_12896_));
 AOI21_X1 _39105_ (.A(_12890_),
    .B1(_12893_),
    .B2(_12896_),
    .ZN(_12897_));
 MUX2_X1 _39106_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [438]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [956]),
    .S(_12840_),
    .Z(_12898_));
 AND2_X1 _39107_ (.A1(_12898_),
    .A2(_12877_),
    .ZN(_12899_));
 NAND2_X1 _39108_ (.A1(_12742_),
    .A2(_12899_),
    .ZN(_12900_));
 MUX2_X1 _39109_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [502]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1020]),
    .S(_12840_),
    .Z(_12901_));
 AND2_X1 _39110_ (.A1(_12901_),
    .A2(_12877_),
    .ZN(_12902_));
 OAI21_X1 _39111_ (.A(_12902_),
    .B1(_12780_),
    .B2(_12781_),
    .ZN(_12903_));
 AOI21_X1 _39112_ (.A(_12596_),
    .B1(_12900_),
    .B2(_12903_),
    .ZN(_12904_));
 OR2_X4 _39113_ (.A1(_12897_),
    .A2(_12904_),
    .ZN(_12905_));
 MUX2_X2 _39114_ (.A(_12889_),
    .B(_12905_),
    .S(_12337_),
    .Z(\icache.data_mem_data_li [48]));
 BUF_X4 _39115_ (.A(_12421_),
    .Z(_12906_));
 MUX2_X2 _39116_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [311]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [829]),
    .S(_12840_),
    .Z(_12907_));
 AND2_X1 _39117_ (.A1(_12907_),
    .A2(_12877_),
    .ZN(_12908_));
 NAND2_X1 _39118_ (.A1(_12906_),
    .A2(_12908_),
    .ZN(_12909_));
 BUF_X16 _39119_ (.A(_11263_),
    .Z(_12910_));
 MUX2_X2 _39120_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [375]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [893]),
    .S(_12910_),
    .Z(_12911_));
 AND2_X1 _39121_ (.A1(_12911_),
    .A2(_12877_),
    .ZN(_12912_));
 OAI21_X1 _39122_ (.A(_12912_),
    .B1(_12780_),
    .B2(_12781_),
    .ZN(_12913_));
 AOI21_X1 _39123_ (.A(_12675_),
    .B1(_12909_),
    .B2(_12913_),
    .ZN(_12914_));
 MUX2_X2 _39124_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [439]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [957]),
    .S(_12881_),
    .Z(_12915_));
 BUF_X4 _39125_ (.A(_12079_),
    .Z(_12916_));
 AND2_X1 _39126_ (.A1(_12915_),
    .A2(_12916_),
    .ZN(_12917_));
 NAND2_X1 _39127_ (.A1(_12808_),
    .A2(_12917_),
    .ZN(_12918_));
 MUX2_X2 _39128_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [503]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1021]),
    .S(_12881_),
    .Z(_12919_));
 AND2_X1 _39129_ (.A1(_12919_),
    .A2(_12916_),
    .ZN(_12920_));
 OAI21_X1 _39130_ (.A(_12920_),
    .B1(_12853_),
    .B2(_12854_),
    .ZN(_12921_));
 AOI21_X1 _39131_ (.A(_12717_),
    .B1(_12918_),
    .B2(_12921_),
    .ZN(_12922_));
 OR2_X4 _39132_ (.A1(_12914_),
    .A2(_12922_),
    .ZN(_12923_));
 MUX2_X1 _39133_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [55]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [573]),
    .S(_12305_),
    .Z(_12924_));
 AND2_X4 _39134_ (.A1(_12924_),
    .A2(_08500_),
    .ZN(_12925_));
 NAND2_X1 _39135_ (.A1(_12808_),
    .A2(_12925_),
    .ZN(_12926_));
 MUX2_X2 _39136_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [119]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [637]),
    .S(_12881_),
    .Z(_12927_));
 AND2_X1 _39137_ (.A1(_12927_),
    .A2(_12916_),
    .ZN(_12928_));
 OAI21_X1 _39138_ (.A(_12928_),
    .B1(_12853_),
    .B2(_12854_),
    .ZN(_12929_));
 AOI21_X1 _39139_ (.A(_12890_),
    .B1(_12926_),
    .B2(_12929_),
    .ZN(_12930_));
 BUF_X8 _39140_ (.A(_08493_),
    .Z(_12931_));
 MUX2_X1 _39141_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [183]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [701]),
    .S(_12840_),
    .Z(_12932_));
 AND2_X1 _39142_ (.A1(_12932_),
    .A2(_12877_),
    .ZN(_12933_));
 NAND2_X1 _39143_ (.A1(_12906_),
    .A2(_12933_),
    .ZN(_12934_));
 MUX2_X1 _39144_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [247]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [765]),
    .S(_12840_),
    .Z(_12935_));
 AND2_X2 _39145_ (.A1(_12935_),
    .A2(_12877_),
    .ZN(_12936_));
 OAI21_X1 _39146_ (.A(_12936_),
    .B1(_12780_),
    .B2(_12781_),
    .ZN(_12937_));
 AOI21_X1 _39147_ (.A(_12931_),
    .B1(_12934_),
    .B2(_12937_),
    .ZN(_12938_));
 OR2_X4 _39148_ (.A1(_12930_),
    .A2(_12938_),
    .ZN(_12939_));
 MUX2_X2 _39149_ (.A(_12923_),
    .B(_12939_),
    .S(_12641_),
    .Z(\icache.data_mem_data_li [49]));
 MUX2_X2 _39150_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [312]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [830]),
    .S(_12881_),
    .Z(_12940_));
 AND2_X1 _39151_ (.A1(_12940_),
    .A2(_12916_),
    .ZN(_12941_));
 NAND2_X1 _39152_ (.A1(_12808_),
    .A2(_12941_),
    .ZN(_12942_));
 MUX2_X1 _39153_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [376]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [894]),
    .S(_12881_),
    .Z(_12943_));
 AND2_X2 _39154_ (.A1(_12943_),
    .A2(_12916_),
    .ZN(_12944_));
 OAI21_X1 _39155_ (.A(_12944_),
    .B1(_12853_),
    .B2(_12854_),
    .ZN(_12945_));
 AOI21_X1 _39156_ (.A(_12675_),
    .B1(_12942_),
    .B2(_12945_),
    .ZN(_12946_));
 MUX2_X2 _39157_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [440]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [958]),
    .S(_12881_),
    .Z(_12947_));
 AND2_X1 _39158_ (.A1(_12947_),
    .A2(_12916_),
    .ZN(_12948_));
 NAND2_X1 _39159_ (.A1(_12808_),
    .A2(_12948_),
    .ZN(_12949_));
 BUF_X8 _39160_ (.A(_11241_),
    .Z(_12950_));
 MUX2_X2 _39161_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [504]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1022]),
    .S(_12950_),
    .Z(_12951_));
 AND2_X2 _39162_ (.A1(_12951_),
    .A2(_12916_),
    .ZN(_12952_));
 OAI21_X1 _39163_ (.A(_12952_),
    .B1(_12853_),
    .B2(_12854_),
    .ZN(_12953_));
 AOI21_X1 _39164_ (.A(_12717_),
    .B1(_12949_),
    .B2(_12953_),
    .ZN(_12954_));
 OR2_X4 _39165_ (.A1(_12946_),
    .A2(_12954_),
    .ZN(_12955_));
 MUX2_X2 _39166_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [56]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [574]),
    .S(_12423_),
    .Z(_12956_));
 AND2_X4 _39167_ (.A1(_12956_),
    .A2(_12643_),
    .ZN(_12957_));
 NAND2_X1 _39168_ (.A1(_12906_),
    .A2(_12957_),
    .ZN(_12958_));
 MUX2_X2 _39169_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [120]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [638]),
    .S(_12910_),
    .Z(_12959_));
 AND2_X1 _39170_ (.A1(_12959_),
    .A2(_12877_),
    .ZN(_12960_));
 BUF_X4 _39171_ (.A(_12610_),
    .Z(_12961_));
 BUF_X4 _39172_ (.A(_12612_),
    .Z(_12962_));
 OAI21_X1 _39173_ (.A(_12960_),
    .B1(_12961_),
    .B2(_12962_),
    .ZN(_12963_));
 AOI21_X1 _39174_ (.A(_12890_),
    .B1(_12958_),
    .B2(_12963_),
    .ZN(_12964_));
 MUX2_X2 _39175_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [184]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [702]),
    .S(_12910_),
    .Z(_12965_));
 AND2_X2 _39176_ (.A1(_12965_),
    .A2(_12877_),
    .ZN(_12966_));
 NAND2_X1 _39177_ (.A1(_12906_),
    .A2(_12966_),
    .ZN(_12967_));
 MUX2_X1 _39178_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [248]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [766]),
    .S(_12910_),
    .Z(_12968_));
 AND2_X1 _39179_ (.A1(_12968_),
    .A2(_12877_),
    .ZN(_12969_));
 OAI21_X1 _39180_ (.A(_12969_),
    .B1(_12961_),
    .B2(_12962_),
    .ZN(_12970_));
 AOI21_X1 _39181_ (.A(_12931_),
    .B1(_12967_),
    .B2(_12970_),
    .ZN(_12971_));
 OR2_X4 _39182_ (.A1(_12964_),
    .A2(_12971_),
    .ZN(_12972_));
 MUX2_X2 _39183_ (.A(_12955_),
    .B(_12972_),
    .S(_12641_),
    .Z(\icache.data_mem_data_li [50]));
 BUF_X32 _39184_ (.A(_08489_),
    .Z(_12973_));
 BUF_X4 _39185_ (.A(_12973_),
    .Z(_12974_));
 MUX2_X2 _39186_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [313]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [831]),
    .S(_12950_),
    .Z(_12975_));
 AND2_X1 _39187_ (.A1(_12975_),
    .A2(_12916_),
    .ZN(_12976_));
 NAND2_X1 _39188_ (.A1(_12974_),
    .A2(_12976_),
    .ZN(_12977_));
 MUX2_X1 _39189_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [377]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [895]),
    .S(_12950_),
    .Z(_12978_));
 AND2_X1 _39190_ (.A1(_12978_),
    .A2(_12916_),
    .ZN(_12979_));
 OAI21_X1 _39191_ (.A(_12979_),
    .B1(_12853_),
    .B2(_12854_),
    .ZN(_12980_));
 AOI21_X1 _39192_ (.A(_12675_),
    .B1(_12977_),
    .B2(_12980_),
    .ZN(_12981_));
 MUX2_X2 _39193_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [441]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [959]),
    .S(_12950_),
    .Z(_12982_));
 AND2_X1 _39194_ (.A1(_12982_),
    .A2(_12916_),
    .ZN(_12983_));
 NAND2_X1 _39195_ (.A1(_12974_),
    .A2(_12983_),
    .ZN(_12984_));
 MUX2_X2 _39196_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [505]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1023]),
    .S(_12950_),
    .Z(_12985_));
 BUF_X2 _39197_ (.A(_11244_),
    .Z(_12986_));
 AND2_X1 _39198_ (.A1(_12985_),
    .A2(_12986_),
    .ZN(_12987_));
 OAI21_X1 _39199_ (.A(_12987_),
    .B1(_12853_),
    .B2(_12854_),
    .ZN(_12988_));
 AOI21_X1 _39200_ (.A(_12717_),
    .B1(_12984_),
    .B2(_12988_),
    .ZN(_12989_));
 OR2_X4 _39201_ (.A1(_12981_),
    .A2(_12989_),
    .ZN(_12990_));
 MUX2_X1 _39202_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [57]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [575]),
    .S(_11311_),
    .Z(_12991_));
 AND2_X4 _39203_ (.A1(_12991_),
    .A2(_12643_),
    .ZN(_12992_));
 NAND2_X1 _39204_ (.A1(_12906_),
    .A2(_12992_),
    .ZN(_12993_));
 MUX2_X2 _39205_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [121]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [639]),
    .S(_12910_),
    .Z(_12994_));
 BUF_X2 _39206_ (.A(_12298_),
    .Z(_12995_));
 AND2_X1 _39207_ (.A1(_12994_),
    .A2(_12995_),
    .ZN(_12996_));
 OAI21_X1 _39208_ (.A(_12996_),
    .B1(_12961_),
    .B2(_12962_),
    .ZN(_12997_));
 AOI21_X1 _39209_ (.A(_12890_),
    .B1(_12993_),
    .B2(_12997_),
    .ZN(_12998_));
 MUX2_X1 _39210_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [185]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [703]),
    .S(_12910_),
    .Z(_12999_));
 AND2_X1 _39211_ (.A1(_12999_),
    .A2(_12995_),
    .ZN(_13000_));
 NAND2_X1 _39212_ (.A1(_12906_),
    .A2(_13000_),
    .ZN(_13001_));
 MUX2_X2 _39213_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [249]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [767]),
    .S(_12910_),
    .Z(_13002_));
 AND2_X1 _39214_ (.A1(_13002_),
    .A2(_12995_),
    .ZN(_13003_));
 OAI21_X1 _39215_ (.A(_13003_),
    .B1(_12961_),
    .B2(_12962_),
    .ZN(_13004_));
 AOI21_X1 _39216_ (.A(_12931_),
    .B1(_13001_),
    .B2(_13004_),
    .ZN(_13005_));
 OR2_X4 _39217_ (.A1(_12998_),
    .A2(_13005_),
    .ZN(_13006_));
 MUX2_X2 _39218_ (.A(_12990_),
    .B(_13006_),
    .S(_12641_),
    .Z(\icache.data_mem_data_li [51]));
 BUF_X8 _39219_ (.A(_11665_),
    .Z(_13007_));
 MUX2_X1 _39220_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [58]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [576]),
    .S(_11311_),
    .Z(_13008_));
 AND2_X4 _39221_ (.A1(_13008_),
    .A2(_12643_),
    .ZN(_13009_));
 NAND2_X1 _39222_ (.A1(_12906_),
    .A2(_13009_),
    .ZN(_13010_));
 MUX2_X2 _39223_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [122]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [640]),
    .S(_12910_),
    .Z(_13011_));
 AND2_X1 _39224_ (.A1(_13011_),
    .A2(_12995_),
    .ZN(_13012_));
 OAI21_X2 _39225_ (.A(_13012_),
    .B1(_12961_),
    .B2(_12962_),
    .ZN(_13013_));
 AOI21_X1 _39226_ (.A(_13007_),
    .B1(_13010_),
    .B2(_13013_),
    .ZN(_13014_));
 MUX2_X2 _39227_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [186]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [704]),
    .S(_12950_),
    .Z(_13015_));
 AND2_X1 _39228_ (.A1(_13015_),
    .A2(_12986_),
    .ZN(_13016_));
 NAND2_X1 _39229_ (.A1(_12974_),
    .A2(_13016_),
    .ZN(_13017_));
 MUX2_X2 _39230_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [250]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [768]),
    .S(_12950_),
    .Z(_13018_));
 AND2_X1 _39231_ (.A1(_13018_),
    .A2(_12986_),
    .ZN(_13019_));
 BUF_X4 _39232_ (.A(_11680_),
    .Z(_13020_));
 BUF_X4 _39233_ (.A(_11682_),
    .Z(_13021_));
 OAI21_X1 _39234_ (.A(_13019_),
    .B1(_13020_),
    .B2(_13021_),
    .ZN(_13022_));
 AOI21_X1 _39235_ (.A(_12717_),
    .B1(_13017_),
    .B2(_13022_),
    .ZN(_13023_));
 OR2_X4 _39236_ (.A1(_13014_),
    .A2(_13023_),
    .ZN(_13024_));
 MUX2_X2 _39237_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [314]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [832]),
    .S(_12950_),
    .Z(_13025_));
 AND2_X1 _39238_ (.A1(_13025_),
    .A2(_12986_),
    .ZN(_13026_));
 NAND2_X1 _39239_ (.A1(_12974_),
    .A2(_13026_),
    .ZN(_13027_));
 MUX2_X1 _39240_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [378]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [896]),
    .S(_12950_),
    .Z(_13028_));
 AND2_X1 _39241_ (.A1(_13028_),
    .A2(_12986_),
    .ZN(_13029_));
 OAI21_X1 _39242_ (.A(_13029_),
    .B1(_13020_),
    .B2(_13021_),
    .ZN(_13030_));
 AOI21_X1 _39243_ (.A(_12890_),
    .B1(_13027_),
    .B2(_13030_),
    .ZN(_13031_));
 MUX2_X1 _39244_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [442]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [960]),
    .S(_12910_),
    .Z(_13032_));
 AND2_X1 _39245_ (.A1(_13032_),
    .A2(_12995_),
    .ZN(_13033_));
 NAND2_X1 _39246_ (.A1(_12906_),
    .A2(_13033_),
    .ZN(_13034_));
 MUX2_X2 _39247_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [506]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1024]),
    .S(_12910_),
    .Z(_13035_));
 AND2_X1 _39248_ (.A1(_13035_),
    .A2(_12995_),
    .ZN(_13036_));
 OAI21_X1 _39249_ (.A(_13036_),
    .B1(_12961_),
    .B2(_12962_),
    .ZN(_13037_));
 AOI21_X1 _39250_ (.A(_12931_),
    .B1(_13034_),
    .B2(_13037_),
    .ZN(_13038_));
 OR2_X4 _39251_ (.A1(_13031_),
    .A2(_13038_),
    .ZN(_13039_));
 MUX2_X2 _39252_ (.A(_13024_),
    .B(_13039_),
    .S(_12337_),
    .Z(\icache.data_mem_data_li [52]));
 MUX2_X2 _39253_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [315]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [833]),
    .S(_12950_),
    .Z(_13040_));
 AND2_X1 _39254_ (.A1(_13040_),
    .A2(_12986_),
    .ZN(_13041_));
 NAND2_X1 _39255_ (.A1(_12974_),
    .A2(_13041_),
    .ZN(_13042_));
 BUF_X8 _39256_ (.A(_11241_),
    .Z(_13043_));
 MUX2_X1 _39257_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [379]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [897]),
    .S(_13043_),
    .Z(_13044_));
 AND2_X1 _39258_ (.A1(_13044_),
    .A2(_12986_),
    .ZN(_13045_));
 OAI21_X1 _39259_ (.A(_13045_),
    .B1(_13020_),
    .B2(_13021_),
    .ZN(_13046_));
 AOI21_X1 _39260_ (.A(_13007_),
    .B1(_13042_),
    .B2(_13046_),
    .ZN(_13047_));
 BUF_X8 _39261_ (.A(_11709_),
    .Z(_13048_));
 MUX2_X2 _39262_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [443]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [961]),
    .S(_13043_),
    .Z(_13049_));
 AND2_X1 _39263_ (.A1(_13049_),
    .A2(_12986_),
    .ZN(_13050_));
 NAND2_X1 _39264_ (.A1(_12974_),
    .A2(_13050_),
    .ZN(_13051_));
 MUX2_X1 _39265_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [507]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1025]),
    .S(_13043_),
    .Z(_13052_));
 AND2_X1 _39266_ (.A1(_13052_),
    .A2(_12986_),
    .ZN(_13053_));
 OAI21_X1 _39267_ (.A(_13053_),
    .B1(_13020_),
    .B2(_13021_),
    .ZN(_13054_));
 AOI21_X1 _39268_ (.A(_13048_),
    .B1(_13051_),
    .B2(_13054_),
    .ZN(_13055_));
 OR2_X4 _39269_ (.A1(_13047_),
    .A2(_13055_),
    .ZN(_13056_));
 MUX2_X2 _39270_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [59]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [577]),
    .S(_11311_),
    .Z(_13057_));
 AND2_X4 _39271_ (.A1(_13057_),
    .A2(_12643_),
    .ZN(_13058_));
 NAND2_X1 _39272_ (.A1(_12906_),
    .A2(_13058_),
    .ZN(_13059_));
 BUF_X16 _39273_ (.A(_11263_),
    .Z(_13060_));
 MUX2_X2 _39274_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [123]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [641]),
    .S(_13060_),
    .Z(_13061_));
 AND2_X1 _39275_ (.A1(_13061_),
    .A2(_12995_),
    .ZN(_13062_));
 OAI21_X1 _39276_ (.A(_13062_),
    .B1(_12961_),
    .B2(_12962_),
    .ZN(_13063_));
 AOI21_X1 _39277_ (.A(_12890_),
    .B1(_13059_),
    .B2(_13063_),
    .ZN(_13064_));
 MUX2_X2 _39278_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [187]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [705]),
    .S(_13060_),
    .Z(_13065_));
 AND2_X1 _39279_ (.A1(_13065_),
    .A2(_12995_),
    .ZN(_13066_));
 NAND2_X1 _39280_ (.A1(_12906_),
    .A2(_13066_),
    .ZN(_13067_));
 MUX2_X2 _39281_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [251]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [769]),
    .S(_13060_),
    .Z(_13068_));
 AND2_X1 _39282_ (.A1(_13068_),
    .A2(_12995_),
    .ZN(_13069_));
 OAI21_X1 _39283_ (.A(_13069_),
    .B1(_12961_),
    .B2(_12962_),
    .ZN(_13070_));
 AOI21_X1 _39284_ (.A(_12931_),
    .B1(_13067_),
    .B2(_13070_),
    .ZN(_13071_));
 OR2_X4 _39285_ (.A1(_13064_),
    .A2(_13071_),
    .ZN(_13072_));
 MUX2_X2 _39286_ (.A(_13056_),
    .B(_13072_),
    .S(_12641_),
    .Z(\icache.data_mem_data_li [53]));
 MUX2_X2 _39287_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [60]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [578]),
    .S(_12305_),
    .Z(_13073_));
 AND2_X4 _39288_ (.A1(_13073_),
    .A2(_08500_),
    .ZN(_13074_));
 NAND2_X1 _39289_ (.A1(_12974_),
    .A2(_13074_),
    .ZN(_13075_));
 MUX2_X1 _39290_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [124]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [642]),
    .S(_13043_),
    .Z(_13076_));
 BUF_X4 _39291_ (.A(_11244_),
    .Z(_13077_));
 AND2_X1 _39292_ (.A1(_13076_),
    .A2(_13077_),
    .ZN(_13078_));
 OAI21_X1 _39293_ (.A(_13078_),
    .B1(_13020_),
    .B2(_13021_),
    .ZN(_13079_));
 AOI21_X1 _39294_ (.A(_13007_),
    .B1(_13075_),
    .B2(_13079_),
    .ZN(_13080_));
 MUX2_X2 _39295_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [188]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [706]),
    .S(_13060_),
    .Z(_13081_));
 BUF_X4 _39296_ (.A(_12298_),
    .Z(_13082_));
 AND2_X1 _39297_ (.A1(_13081_),
    .A2(_13082_),
    .ZN(_13083_));
 NAND2_X1 _39298_ (.A1(_12974_),
    .A2(_13083_),
    .ZN(_13084_));
 MUX2_X2 _39299_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [252]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [770]),
    .S(_13043_),
    .Z(_13085_));
 AND2_X2 _39300_ (.A1(_13085_),
    .A2(_13077_),
    .ZN(_13086_));
 OAI21_X1 _39301_ (.A(_13086_),
    .B1(_13020_),
    .B2(_13021_),
    .ZN(_13087_));
 AOI21_X1 _39302_ (.A(_13048_),
    .B1(_13084_),
    .B2(_13087_),
    .ZN(_13088_));
 OR2_X4 _39303_ (.A1(_13080_),
    .A2(_13088_),
    .ZN(_13089_));
 BUF_X4 _39304_ (.A(_12421_),
    .Z(_13090_));
 MUX2_X2 _39305_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [316]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [834]),
    .S(_13060_),
    .Z(_13091_));
 AND2_X1 _39306_ (.A1(_13091_),
    .A2(_12995_),
    .ZN(_13092_));
 NAND2_X1 _39307_ (.A1(_13090_),
    .A2(_13092_),
    .ZN(_13093_));
 MUX2_X2 _39308_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [380]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [898]),
    .S(_13060_),
    .Z(_13094_));
 AND2_X1 _39309_ (.A1(_13094_),
    .A2(_13082_),
    .ZN(_13095_));
 OAI21_X1 _39310_ (.A(_13095_),
    .B1(_12961_),
    .B2(_12962_),
    .ZN(_13096_));
 AOI21_X1 _39311_ (.A(_12890_),
    .B1(_13093_),
    .B2(_13096_),
    .ZN(_13097_));
 MUX2_X2 _39312_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [444]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [962]),
    .S(_13043_),
    .Z(_13098_));
 AND2_X2 _39313_ (.A1(_13098_),
    .A2(_12986_),
    .ZN(_13099_));
 NAND2_X1 _39314_ (.A1(_13090_),
    .A2(_13099_),
    .ZN(_13100_));
 MUX2_X2 _39315_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [508]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1026]),
    .S(_13060_),
    .Z(_13101_));
 AND2_X1 _39316_ (.A1(_13101_),
    .A2(_13082_),
    .ZN(_13102_));
 OAI21_X1 _39317_ (.A(_13102_),
    .B1(_12961_),
    .B2(_12962_),
    .ZN(_13103_));
 AOI21_X1 _39318_ (.A(_12931_),
    .B1(_13100_),
    .B2(_13103_),
    .ZN(_13104_));
 OR2_X4 _39319_ (.A1(_13097_),
    .A2(_13104_),
    .ZN(_13105_));
 MUX2_X2 _39320_ (.A(_13089_),
    .B(_13105_),
    .S(_12337_),
    .Z(\icache.data_mem_data_li [54]));
 MUX2_X2 _39321_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [317]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [835]),
    .S(_13043_),
    .Z(_13106_));
 AND2_X1 _39322_ (.A1(_13106_),
    .A2(_13077_),
    .ZN(_13107_));
 NAND2_X1 _39323_ (.A1(_12974_),
    .A2(_13107_),
    .ZN(_13108_));
 MUX2_X1 _39324_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [381]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [899]),
    .S(_13043_),
    .Z(_13109_));
 AND2_X1 _39325_ (.A1(_13109_),
    .A2(_13077_),
    .ZN(_13110_));
 OAI21_X1 _39326_ (.A(_13110_),
    .B1(_13020_),
    .B2(_13021_),
    .ZN(_13111_));
 AOI21_X1 _39327_ (.A(_13007_),
    .B1(_13108_),
    .B2(_13111_),
    .ZN(_13112_));
 MUX2_X2 _39328_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [445]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [963]),
    .S(_13043_),
    .Z(_13113_));
 AND2_X1 _39329_ (.A1(_13113_),
    .A2(_13077_),
    .ZN(_13114_));
 NAND2_X1 _39330_ (.A1(_12974_),
    .A2(_13114_),
    .ZN(_13115_));
 MUX2_X1 _39331_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [509]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1027]),
    .S(_13043_),
    .Z(_13116_));
 AND2_X1 _39332_ (.A1(_13116_),
    .A2(_13077_),
    .ZN(_13117_));
 OAI21_X1 _39333_ (.A(_13117_),
    .B1(_13020_),
    .B2(_13021_),
    .ZN(_13118_));
 AOI21_X1 _39334_ (.A(_13048_),
    .B1(_13115_),
    .B2(_13118_),
    .ZN(_13119_));
 OR2_X4 _39335_ (.A1(_13112_),
    .A2(_13119_),
    .ZN(_13120_));
 MUX2_X2 _39336_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [61]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [579]),
    .S(_11311_),
    .Z(_13121_));
 AND2_X4 _39337_ (.A1(_13121_),
    .A2(_12643_),
    .ZN(_13122_));
 NAND2_X1 _39338_ (.A1(_13090_),
    .A2(_13122_),
    .ZN(_13123_));
 MUX2_X1 _39339_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [125]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [643]),
    .S(_13060_),
    .Z(_13124_));
 AND2_X1 _39340_ (.A1(_13124_),
    .A2(_13082_),
    .ZN(_13125_));
 BUF_X4 _39341_ (.A(_12610_),
    .Z(_13126_));
 BUF_X4 _39342_ (.A(_12612_),
    .Z(_13127_));
 OAI21_X1 _39343_ (.A(_13125_),
    .B1(_13126_),
    .B2(_13127_),
    .ZN(_13128_));
 AOI21_X1 _39344_ (.A(_12890_),
    .B1(_13123_),
    .B2(_13128_),
    .ZN(_13129_));
 MUX2_X2 _39345_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [189]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [707]),
    .S(_13060_),
    .Z(_13130_));
 AND2_X1 _39346_ (.A1(_13130_),
    .A2(_13082_),
    .ZN(_13131_));
 NAND2_X1 _39347_ (.A1(_13090_),
    .A2(_13131_),
    .ZN(_13132_));
 MUX2_X2 _39348_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [253]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [771]),
    .S(_13060_),
    .Z(_13133_));
 AND2_X2 _39349_ (.A1(_13133_),
    .A2(_13082_),
    .ZN(_13134_));
 OAI21_X1 _39350_ (.A(_13134_),
    .B1(_13126_),
    .B2(_13127_),
    .ZN(_13135_));
 AOI21_X1 _39351_ (.A(_12931_),
    .B1(_13132_),
    .B2(_13135_),
    .ZN(_13136_));
 OR2_X4 _39352_ (.A1(_13129_),
    .A2(_13136_),
    .ZN(_13137_));
 MUX2_X2 _39353_ (.A(_13120_),
    .B(_13137_),
    .S(_12641_),
    .Z(\icache.data_mem_data_li [55]));
 BUF_X16 _39354_ (.A(_11263_),
    .Z(_13138_));
 MUX2_X2 _39355_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [318]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [836]),
    .S(_13138_),
    .Z(_13139_));
 AND2_X1 _39356_ (.A1(_13139_),
    .A2(_13082_),
    .ZN(_13140_));
 NAND2_X1 _39357_ (.A1(_13090_),
    .A2(_13140_),
    .ZN(_13141_));
 MUX2_X2 _39358_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [382]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [900]),
    .S(_13138_),
    .Z(_13142_));
 AND2_X1 _39359_ (.A1(_13142_),
    .A2(_13082_),
    .ZN(_13143_));
 OAI21_X1 _39360_ (.A(_13143_),
    .B1(_13126_),
    .B2(_13127_),
    .ZN(_13144_));
 AOI21_X1 _39361_ (.A(_13007_),
    .B1(_13141_),
    .B2(_13144_),
    .ZN(_13145_));
 BUF_X4 _39362_ (.A(_12973_),
    .Z(_13146_));
 BUF_X8 _39363_ (.A(_11241_),
    .Z(_13147_));
 MUX2_X1 _39364_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [446]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [964]),
    .S(_13147_),
    .Z(_13148_));
 AND2_X1 _39365_ (.A1(_13148_),
    .A2(_13077_),
    .ZN(_13149_));
 NAND2_X1 _39366_ (.A1(_13146_),
    .A2(_13149_),
    .ZN(_13150_));
 MUX2_X1 _39367_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [510]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1028]),
    .S(_13147_),
    .Z(_13151_));
 AND2_X1 _39368_ (.A1(_13151_),
    .A2(_13077_),
    .ZN(_13152_));
 OAI21_X1 _39369_ (.A(_13152_),
    .B1(_13020_),
    .B2(_13021_),
    .ZN(_13153_));
 AOI21_X1 _39370_ (.A(_13048_),
    .B1(_13150_),
    .B2(_13153_),
    .ZN(_13154_));
 OR2_X4 _39371_ (.A1(_13145_),
    .A2(_13154_),
    .ZN(_13155_));
 MUX2_X2 _39372_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [62]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [580]),
    .S(_08428_),
    .Z(_13156_));
 AND2_X4 _39373_ (.A1(_13156_),
    .A2(_08500_),
    .ZN(_13157_));
 NAND2_X1 _39374_ (.A1(_13146_),
    .A2(_13157_),
    .ZN(_13158_));
 MUX2_X2 _39375_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [126]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [644]),
    .S(_13147_),
    .Z(_13159_));
 AND2_X1 _39376_ (.A1(_13159_),
    .A2(_13077_),
    .ZN(_13160_));
 OAI21_X1 _39377_ (.A(_13160_),
    .B1(_13020_),
    .B2(_13021_),
    .ZN(_13161_));
 AOI21_X1 _39378_ (.A(_12890_),
    .B1(_13158_),
    .B2(_13161_),
    .ZN(_13162_));
 MUX2_X2 _39379_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [190]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [708]),
    .S(_13138_),
    .Z(_13163_));
 AND2_X1 _39380_ (.A1(_13163_),
    .A2(_13082_),
    .ZN(_13164_));
 NAND2_X1 _39381_ (.A1(_13090_),
    .A2(_13164_),
    .ZN(_13165_));
 MUX2_X2 _39382_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [254]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [772]),
    .S(_13138_),
    .Z(_13166_));
 AND2_X1 _39383_ (.A1(_13166_),
    .A2(_13082_),
    .ZN(_13167_));
 OAI21_X1 _39384_ (.A(_13167_),
    .B1(_13126_),
    .B2(_13127_),
    .ZN(_13168_));
 AOI21_X1 _39385_ (.A(_12931_),
    .B1(_13165_),
    .B2(_13168_),
    .ZN(_13169_));
 OR2_X4 _39386_ (.A1(_13162_),
    .A2(_13169_),
    .ZN(_13170_));
 BUF_X32 _39387_ (.A(_12640_),
    .Z(_13171_));
 MUX2_X2 _39388_ (.A(_13155_),
    .B(_13170_),
    .S(_13171_),
    .Z(\icache.data_mem_data_li [56]));
 MUX2_X2 _39389_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [319]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [837]),
    .S(_13147_),
    .Z(_13172_));
 BUF_X4 _39390_ (.A(_11244_),
    .Z(_13173_));
 AND2_X1 _39391_ (.A1(_13172_),
    .A2(_13173_),
    .ZN(_13174_));
 NAND2_X1 _39392_ (.A1(_13146_),
    .A2(_13174_),
    .ZN(_13175_));
 MUX2_X1 _39393_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [383]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [901]),
    .S(_13147_),
    .Z(_13176_));
 AND2_X1 _39394_ (.A1(_13176_),
    .A2(_13173_),
    .ZN(_13177_));
 BUF_X4 _39395_ (.A(_11680_),
    .Z(_13178_));
 BUF_X4 _39396_ (.A(_11682_),
    .Z(_13179_));
 OAI21_X1 _39397_ (.A(_13177_),
    .B1(_13178_),
    .B2(_13179_),
    .ZN(_13180_));
 AOI21_X1 _39398_ (.A(_13007_),
    .B1(_13175_),
    .B2(_13180_),
    .ZN(_13181_));
 MUX2_X1 _39399_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [447]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [965]),
    .S(_13138_),
    .Z(_13182_));
 BUF_X4 _39400_ (.A(_12298_),
    .Z(_13183_));
 AND2_X1 _39401_ (.A1(_13182_),
    .A2(_13183_),
    .ZN(_13184_));
 NAND2_X1 _39402_ (.A1(_13146_),
    .A2(_13184_),
    .ZN(_13185_));
 MUX2_X1 _39403_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [511]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1029]),
    .S(_13147_),
    .Z(_13186_));
 AND2_X1 _39404_ (.A1(_13186_),
    .A2(_13173_),
    .ZN(_13187_));
 OAI21_X1 _39405_ (.A(_13187_),
    .B1(_13178_),
    .B2(_13179_),
    .ZN(_13188_));
 AOI21_X1 _39406_ (.A(_13048_),
    .B1(_13185_),
    .B2(_13188_),
    .ZN(_13189_));
 OR2_X4 _39407_ (.A1(_13181_),
    .A2(_13189_),
    .ZN(_13190_));
 MUX2_X2 _39408_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [63]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [581]),
    .S(_11311_),
    .Z(_13191_));
 AND2_X4 _39409_ (.A1(_13191_),
    .A2(_11313_),
    .ZN(_13192_));
 NAND2_X1 _39410_ (.A1(_13090_),
    .A2(_13192_),
    .ZN(_13193_));
 MUX2_X2 _39411_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [127]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [645]),
    .S(_13138_),
    .Z(_13194_));
 AND2_X1 _39412_ (.A1(_13194_),
    .A2(_13183_),
    .ZN(_13195_));
 OAI21_X1 _39413_ (.A(_13195_),
    .B1(_13126_),
    .B2(_13127_),
    .ZN(_13196_));
 AOI21_X1 _39414_ (.A(_12890_),
    .B1(_13193_),
    .B2(_13196_),
    .ZN(_13197_));
 MUX2_X1 _39415_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [191]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [709]),
    .S(_13147_),
    .Z(_13198_));
 AND2_X1 _39416_ (.A1(_13198_),
    .A2(_13077_),
    .ZN(_13199_));
 NAND2_X1 _39417_ (.A1(_13090_),
    .A2(_13199_),
    .ZN(_13200_));
 MUX2_X2 _39418_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [255]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [773]),
    .S(_13138_),
    .Z(_13201_));
 AND2_X1 _39419_ (.A1(_13201_),
    .A2(_13183_),
    .ZN(_13202_));
 OAI21_X1 _39420_ (.A(_13202_),
    .B1(_13126_),
    .B2(_13127_),
    .ZN(_13203_));
 AOI21_X1 _39421_ (.A(_12931_),
    .B1(_13200_),
    .B2(_13203_),
    .ZN(_13204_));
 OR2_X4 _39422_ (.A1(_13197_),
    .A2(_13204_),
    .ZN(_13205_));
 MUX2_X2 _39423_ (.A(_13190_),
    .B(_13205_),
    .S(_13171_),
    .Z(\icache.data_mem_data_li [57]));
 MUX2_X1 _39424_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [320]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [838]),
    .S(_13147_),
    .Z(_13206_));
 AND2_X1 _39425_ (.A1(_13206_),
    .A2(_13173_),
    .ZN(_13207_));
 NAND2_X1 _39426_ (.A1(_13146_),
    .A2(_13207_),
    .ZN(_13208_));
 MUX2_X1 _39427_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [384]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [902]),
    .S(_13147_),
    .Z(_13209_));
 AND2_X1 _39428_ (.A1(_13209_),
    .A2(_13173_),
    .ZN(_13210_));
 OAI21_X1 _39429_ (.A(_13210_),
    .B1(_13178_),
    .B2(_13179_),
    .ZN(_13211_));
 AOI21_X1 _39430_ (.A(_13007_),
    .B1(_13208_),
    .B2(_13211_),
    .ZN(_13212_));
 MUX2_X2 _39431_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [448]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [966]),
    .S(_13138_),
    .Z(_13213_));
 AND2_X1 _39432_ (.A1(_13213_),
    .A2(_13183_),
    .ZN(_13214_));
 NAND2_X1 _39433_ (.A1(_13146_),
    .A2(_13214_),
    .ZN(_13215_));
 BUF_X16 _39434_ (.A(_11241_),
    .Z(_13216_));
 MUX2_X1 _39435_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [512]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1030]),
    .S(_13216_),
    .Z(_13217_));
 AND2_X1 _39436_ (.A1(_13217_),
    .A2(_13173_),
    .ZN(_13218_));
 OAI21_X1 _39437_ (.A(_13218_),
    .B1(_13178_),
    .B2(_13179_),
    .ZN(_13219_));
 AOI21_X1 _39438_ (.A(_13048_),
    .B1(_13215_),
    .B2(_13219_),
    .ZN(_13220_));
 OR2_X2 _39439_ (.A1(_13212_),
    .A2(_13220_),
    .ZN(_13221_));
 BUF_X8 _39440_ (.A(_11546_),
    .Z(_13222_));
 MUX2_X1 _39441_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [64]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [582]),
    .S(_11311_),
    .Z(_13223_));
 AND2_X4 _39442_ (.A1(_13223_),
    .A2(_11313_),
    .ZN(_13224_));
 NAND2_X1 _39443_ (.A1(_13090_),
    .A2(_13224_),
    .ZN(_13225_));
 MUX2_X2 _39444_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [128]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [646]),
    .S(_13138_),
    .Z(_13226_));
 AND2_X1 _39445_ (.A1(_13226_),
    .A2(_13183_),
    .ZN(_13227_));
 OAI21_X1 _39446_ (.A(_13227_),
    .B1(_13126_),
    .B2(_13127_),
    .ZN(_13228_));
 AOI21_X1 _39447_ (.A(_13222_),
    .B1(_13225_),
    .B2(_13228_),
    .ZN(_13229_));
 MUX2_X2 _39448_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [192]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [710]),
    .S(_13147_),
    .Z(_13230_));
 AND2_X1 _39449_ (.A1(_13230_),
    .A2(_13173_),
    .ZN(_13231_));
 NAND2_X1 _39450_ (.A1(_13090_),
    .A2(_13231_),
    .ZN(_13232_));
 MUX2_X2 _39451_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [256]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [774]),
    .S(_13138_),
    .Z(_13233_));
 AND2_X1 _39452_ (.A1(_13233_),
    .A2(_13183_),
    .ZN(_13234_));
 OAI21_X1 _39453_ (.A(_13234_),
    .B1(_13126_),
    .B2(_13127_),
    .ZN(_13235_));
 AOI21_X1 _39454_ (.A(_12931_),
    .B1(_13232_),
    .B2(_13235_),
    .ZN(_13236_));
 OR2_X4 _39455_ (.A1(_13229_),
    .A2(_13236_),
    .ZN(_13237_));
 MUX2_X2 _39456_ (.A(_13221_),
    .B(_13237_),
    .S(_13171_),
    .Z(\icache.data_mem_data_li [58]));
 MUX2_X2 _39457_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [321]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [839]),
    .S(_13216_),
    .Z(_13238_));
 AND2_X1 _39458_ (.A1(_13238_),
    .A2(_13173_),
    .ZN(_13239_));
 NAND2_X1 _39459_ (.A1(_13146_),
    .A2(_13239_),
    .ZN(_13240_));
 MUX2_X2 _39460_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [385]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [903]),
    .S(_13216_),
    .Z(_13241_));
 AND2_X1 _39461_ (.A1(_13241_),
    .A2(_13173_),
    .ZN(_13242_));
 OAI21_X1 _39462_ (.A(_13242_),
    .B1(_13178_),
    .B2(_13179_),
    .ZN(_13243_));
 AOI21_X1 _39463_ (.A(_13007_),
    .B1(_13240_),
    .B2(_13243_),
    .ZN(_13244_));
 MUX2_X2 _39464_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [449]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [967]),
    .S(_13216_),
    .Z(_13245_));
 AND2_X1 _39465_ (.A1(_13245_),
    .A2(_13173_),
    .ZN(_13246_));
 NAND2_X1 _39466_ (.A1(_13146_),
    .A2(_13246_),
    .ZN(_13247_));
 MUX2_X1 _39467_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [513]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1031]),
    .S(_13216_),
    .Z(_13248_));
 BUF_X4 _39468_ (.A(_11244_),
    .Z(_13249_));
 AND2_X1 _39469_ (.A1(_13248_),
    .A2(_13249_),
    .ZN(_13250_));
 OAI21_X1 _39470_ (.A(_13250_),
    .B1(_13178_),
    .B2(_13179_),
    .ZN(_13251_));
 AOI21_X1 _39471_ (.A(_13048_),
    .B1(_13247_),
    .B2(_13251_),
    .ZN(_13252_));
 OR2_X4 _39472_ (.A1(_13244_),
    .A2(_13252_),
    .ZN(_13253_));
 BUF_X4 _39473_ (.A(_12421_),
    .Z(_13254_));
 MUX2_X2 _39474_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [65]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [583]),
    .S(_11311_),
    .Z(_13255_));
 AND2_X4 _39475_ (.A1(_13255_),
    .A2(_11313_),
    .ZN(_13256_));
 NAND2_X1 _39476_ (.A1(_13254_),
    .A2(_13256_),
    .ZN(_13257_));
 BUF_X16 _39477_ (.A(_11263_),
    .Z(_13258_));
 MUX2_X2 _39478_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [129]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [647]),
    .S(_13258_),
    .Z(_13259_));
 AND2_X1 _39479_ (.A1(_13259_),
    .A2(_13183_),
    .ZN(_13260_));
 OAI21_X2 _39480_ (.A(_13260_),
    .B1(_13126_),
    .B2(_13127_),
    .ZN(_13261_));
 AOI21_X1 _39481_ (.A(_13222_),
    .B1(_13257_),
    .B2(_13261_),
    .ZN(_13262_));
 BUF_X8 _39482_ (.A(_08493_),
    .Z(_13263_));
 MUX2_X2 _39483_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [193]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [711]),
    .S(_13258_),
    .Z(_13264_));
 AND2_X1 _39484_ (.A1(_13264_),
    .A2(_13183_),
    .ZN(_13265_));
 NAND2_X1 _39485_ (.A1(_13254_),
    .A2(_13265_),
    .ZN(_13266_));
 MUX2_X2 _39486_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [257]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [775]),
    .S(_13258_),
    .Z(_13267_));
 AND2_X1 _39487_ (.A1(_13267_),
    .A2(_13183_),
    .ZN(_13268_));
 OAI21_X2 _39488_ (.A(_13268_),
    .B1(_13126_),
    .B2(_13127_),
    .ZN(_13269_));
 AOI21_X1 _39489_ (.A(_13263_),
    .B1(_13266_),
    .B2(_13269_),
    .ZN(_13270_));
 OR2_X4 _39490_ (.A1(_13262_),
    .A2(_13270_),
    .ZN(_13271_));
 MUX2_X2 _39491_ (.A(_13253_),
    .B(_13271_),
    .S(_13171_),
    .Z(\icache.data_mem_data_li [59]));
 MUX2_X2 _39492_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [322]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [840]),
    .S(_13216_),
    .Z(_13272_));
 AND2_X1 _39493_ (.A1(_13272_),
    .A2(_13249_),
    .ZN(_13273_));
 NAND2_X1 _39494_ (.A1(_13146_),
    .A2(_13273_),
    .ZN(_13274_));
 MUX2_X2 _39495_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [386]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [904]),
    .S(_13216_),
    .Z(_13275_));
 AND2_X1 _39496_ (.A1(_13275_),
    .A2(_13249_),
    .ZN(_13276_));
 OAI21_X1 _39497_ (.A(_13276_),
    .B1(_13178_),
    .B2(_13179_),
    .ZN(_13277_));
 AOI21_X1 _39498_ (.A(_13007_),
    .B1(_13274_),
    .B2(_13277_),
    .ZN(_13278_));
 MUX2_X2 _39499_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [450]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [968]),
    .S(_13216_),
    .Z(_13279_));
 AND2_X1 _39500_ (.A1(_13279_),
    .A2(_13249_),
    .ZN(_13280_));
 NAND2_X1 _39501_ (.A1(_13146_),
    .A2(_13280_),
    .ZN(_13281_));
 MUX2_X2 _39502_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [514]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1032]),
    .S(_13216_),
    .Z(_13282_));
 AND2_X1 _39503_ (.A1(_13282_),
    .A2(_13249_),
    .ZN(_13283_));
 OAI21_X1 _39504_ (.A(_13283_),
    .B1(_13178_),
    .B2(_13179_),
    .ZN(_13284_));
 AOI21_X1 _39505_ (.A(_13048_),
    .B1(_13281_),
    .B2(_13284_),
    .ZN(_13285_));
 OR2_X2 _39506_ (.A1(_13278_),
    .A2(_13285_),
    .ZN(_13286_));
 MUX2_X1 _39507_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [66]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [584]),
    .S(_11311_),
    .Z(_13287_));
 AND2_X4 _39508_ (.A1(_13287_),
    .A2(_11313_),
    .ZN(_13288_));
 NAND2_X1 _39509_ (.A1(_13254_),
    .A2(_13288_),
    .ZN(_13289_));
 MUX2_X1 _39510_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [130]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [648]),
    .S(_13258_),
    .Z(_13290_));
 AND2_X1 _39511_ (.A1(_13290_),
    .A2(_13183_),
    .ZN(_13291_));
 BUF_X4 _39512_ (.A(_12610_),
    .Z(_13292_));
 BUF_X4 _39513_ (.A(_12612_),
    .Z(_13293_));
 OAI21_X2 _39514_ (.A(_13291_),
    .B1(_13292_),
    .B2(_13293_),
    .ZN(_13294_));
 AOI21_X1 _39515_ (.A(_13222_),
    .B1(_13289_),
    .B2(_13294_),
    .ZN(_13295_));
 MUX2_X1 _39516_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [194]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [712]),
    .S(_13258_),
    .Z(_13296_));
 BUF_X4 _39517_ (.A(_11266_),
    .Z(_13297_));
 AND2_X1 _39518_ (.A1(_13296_),
    .A2(_13297_),
    .ZN(_13298_));
 NAND2_X1 _39519_ (.A1(_13254_),
    .A2(_13298_),
    .ZN(_13299_));
 MUX2_X2 _39520_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [258]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [776]),
    .S(_13258_),
    .Z(_13300_));
 AND2_X1 _39521_ (.A1(_13300_),
    .A2(_13297_),
    .ZN(_13301_));
 OAI21_X1 _39522_ (.A(_13301_),
    .B1(_13292_),
    .B2(_13293_),
    .ZN(_13302_));
 AOI21_X1 _39523_ (.A(_13263_),
    .B1(_13299_),
    .B2(_13302_),
    .ZN(_13303_));
 OR2_X2 _39524_ (.A1(_13295_),
    .A2(_13303_),
    .ZN(_13304_));
 MUX2_X2 _39525_ (.A(_13286_),
    .B(_13304_),
    .S(_13171_),
    .Z(\icache.data_mem_data_li [60]));
 MUX2_X2 _39526_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [323]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [841]),
    .S(_13258_),
    .Z(_13305_));
 AND2_X1 _39527_ (.A1(_13305_),
    .A2(_13297_),
    .ZN(_13306_));
 NAND2_X1 _39528_ (.A1(_13254_),
    .A2(_13306_),
    .ZN(_13307_));
 MUX2_X2 _39529_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [387]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [905]),
    .S(_13258_),
    .Z(_13308_));
 AND2_X1 _39530_ (.A1(_13308_),
    .A2(_13297_),
    .ZN(_13309_));
 OAI21_X1 _39531_ (.A(_13309_),
    .B1(_13292_),
    .B2(_13293_),
    .ZN(_13310_));
 AOI21_X1 _39532_ (.A(_13007_),
    .B1(_13307_),
    .B2(_13310_),
    .ZN(_13311_));
 BUF_X4 _39533_ (.A(_12973_),
    .Z(_13312_));
 MUX2_X2 _39534_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [451]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [969]),
    .S(_11242_),
    .Z(_13313_));
 AND2_X1 _39535_ (.A1(_13313_),
    .A2(_13249_),
    .ZN(_13314_));
 NAND2_X1 _39536_ (.A1(_13312_),
    .A2(_13314_),
    .ZN(_13315_));
 MUX2_X2 _39537_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [515]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1033]),
    .S(_11242_),
    .Z(_13316_));
 AND2_X1 _39538_ (.A1(_13316_),
    .A2(_13249_),
    .ZN(_13317_));
 OAI21_X1 _39539_ (.A(_13317_),
    .B1(_13178_),
    .B2(_13179_),
    .ZN(_13318_));
 AOI21_X1 _39540_ (.A(_13048_),
    .B1(_13315_),
    .B2(_13318_),
    .ZN(_13319_));
 OR2_X2 _39541_ (.A1(_13311_),
    .A2(_13319_),
    .ZN(_13320_));
 MUX2_X1 _39542_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [67]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [585]),
    .S(_08428_),
    .Z(_13321_));
 AND2_X4 _39543_ (.A1(_13321_),
    .A2(_08500_),
    .ZN(_13322_));
 NAND2_X1 _39544_ (.A1(_13312_),
    .A2(_13322_),
    .ZN(_13323_));
 MUX2_X1 _39545_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [131]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [649]),
    .S(_13216_),
    .Z(_13324_));
 AND2_X1 _39546_ (.A1(_13324_),
    .A2(_13249_),
    .ZN(_13325_));
 OAI21_X2 _39547_ (.A(_13325_),
    .B1(_13178_),
    .B2(_13179_),
    .ZN(_13326_));
 AOI21_X1 _39548_ (.A(_13222_),
    .B1(_13323_),
    .B2(_13326_),
    .ZN(_13327_));
 MUX2_X2 _39549_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [195]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [713]),
    .S(_13258_),
    .Z(_13328_));
 AND2_X1 _39550_ (.A1(_13328_),
    .A2(_13297_),
    .ZN(_13329_));
 NAND2_X1 _39551_ (.A1(_13254_),
    .A2(_13329_),
    .ZN(_13330_));
 MUX2_X2 _39552_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [259]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [777]),
    .S(_13258_),
    .Z(_13331_));
 AND2_X1 _39553_ (.A1(_13331_),
    .A2(_13297_),
    .ZN(_13332_));
 OAI21_X1 _39554_ (.A(_13332_),
    .B1(_13292_),
    .B2(_13293_),
    .ZN(_13333_));
 AOI21_X1 _39555_ (.A(_13263_),
    .B1(_13330_),
    .B2(_13333_),
    .ZN(_13334_));
 OR2_X2 _39556_ (.A1(_13327_),
    .A2(_13334_),
    .ZN(_13335_));
 MUX2_X2 _39557_ (.A(_13320_),
    .B(_13335_),
    .S(_13171_),
    .Z(\icache.data_mem_data_li [61]));
 BUF_X8 _39558_ (.A(_11665_),
    .Z(_13336_));
 MUX2_X1 _39559_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [324]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [842]),
    .S(_11242_),
    .Z(_13337_));
 AND2_X1 _39560_ (.A1(_13337_),
    .A2(_13249_),
    .ZN(_13338_));
 NAND2_X1 _39561_ (.A1(_13312_),
    .A2(_13338_),
    .ZN(_13339_));
 MUX2_X2 _39562_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [388]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [906]),
    .S(_11242_),
    .Z(_13340_));
 AND2_X1 _39563_ (.A1(_13340_),
    .A2(_13249_),
    .ZN(_13341_));
 BUF_X32 _39564_ (.A(_08483_),
    .Z(_13342_));
 BUF_X4 _39565_ (.A(_13342_),
    .Z(_13343_));
 BUF_X32 _39566_ (.A(_08487_),
    .Z(_13344_));
 BUF_X4 _39567_ (.A(_13344_),
    .Z(_13345_));
 OAI21_X1 _39568_ (.A(_13341_),
    .B1(_13343_),
    .B2(_13345_),
    .ZN(_13346_));
 AOI21_X1 _39569_ (.A(_13336_),
    .B1(_13339_),
    .B2(_13346_),
    .ZN(_13347_));
 MUX2_X1 _39570_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [452]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [970]),
    .S(_11242_),
    .Z(_13348_));
 AND2_X4 _39571_ (.A1(_13348_),
    .A2(_11245_),
    .ZN(_13349_));
 NAND2_X1 _39572_ (.A1(_13312_),
    .A2(_13349_),
    .ZN(_13350_));
 MUX2_X1 _39573_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [516]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1034]),
    .S(_11242_),
    .Z(_13351_));
 AND2_X1 _39574_ (.A1(_13351_),
    .A2(_11245_),
    .ZN(_13352_));
 OAI21_X1 _39575_ (.A(_13352_),
    .B1(_13343_),
    .B2(_13345_),
    .ZN(_13353_));
 AOI21_X1 _39576_ (.A(_13048_),
    .B1(_13350_),
    .B2(_13353_),
    .ZN(_13354_));
 OR2_X1 _39577_ (.A1(_13347_),
    .A2(_13354_),
    .ZN(_13355_));
 MUX2_X1 _39578_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [68]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [586]),
    .S(_11311_),
    .Z(_13356_));
 AND2_X4 _39579_ (.A1(_13356_),
    .A2(_11313_),
    .ZN(_13357_));
 NAND2_X1 _39580_ (.A1(_13254_),
    .A2(_13357_),
    .ZN(_13358_));
 MUX2_X1 _39581_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [132]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [650]),
    .S(_11276_),
    .Z(_13359_));
 AND2_X1 _39582_ (.A1(_13359_),
    .A2(_13297_),
    .ZN(_13360_));
 OAI21_X1 _39583_ (.A(_13360_),
    .B1(_13292_),
    .B2(_13293_),
    .ZN(_13361_));
 AOI21_X1 _39584_ (.A(_13222_),
    .B1(_13358_),
    .B2(_13361_),
    .ZN(_13362_));
 MUX2_X2 _39585_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [196]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [714]),
    .S(_11276_),
    .Z(_13363_));
 AND2_X1 _39586_ (.A1(_13363_),
    .A2(_13297_),
    .ZN(_13364_));
 NAND2_X1 _39587_ (.A1(_13254_),
    .A2(_13364_),
    .ZN(_13365_));
 MUX2_X2 _39588_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [260]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [778]),
    .S(_11276_),
    .Z(_13366_));
 AND2_X1 _39589_ (.A1(_13366_),
    .A2(_13297_),
    .ZN(_13367_));
 OAI21_X1 _39590_ (.A(_13367_),
    .B1(_13292_),
    .B2(_13293_),
    .ZN(_13368_));
 AOI21_X1 _39591_ (.A(_13263_),
    .B1(_13365_),
    .B2(_13368_),
    .ZN(_13369_));
 OR2_X1 _39592_ (.A1(_13362_),
    .A2(_13369_),
    .ZN(_13370_));
 MUX2_X2 _39593_ (.A(_13355_),
    .B(_13370_),
    .S(_13171_),
    .Z(\icache.data_mem_data_li [62]));
 MUX2_X2 _39594_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [69]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [587]),
    .S(_08428_),
    .Z(_13371_));
 AND2_X4 _39595_ (.A1(_13371_),
    .A2(_08500_),
    .ZN(_13372_));
 NAND2_X1 _39596_ (.A1(_13312_),
    .A2(_13372_),
    .ZN(_13373_));
 MUX2_X1 _39597_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [133]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [651]),
    .S(_11242_),
    .Z(_13374_));
 AND2_X1 _39598_ (.A1(_13374_),
    .A2(_11245_),
    .ZN(_13375_));
 OAI21_X1 _39599_ (.A(_13375_),
    .B1(_13343_),
    .B2(_13345_),
    .ZN(_13376_));
 AOI21_X1 _39600_ (.A(_13336_),
    .B1(_13373_),
    .B2(_13376_),
    .ZN(_13377_));
 BUF_X8 _39601_ (.A(_11709_),
    .Z(_13378_));
 MUX2_X2 _39602_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [197]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [715]),
    .S(_11242_),
    .Z(_13379_));
 AND2_X1 _39603_ (.A1(_13379_),
    .A2(_11245_),
    .ZN(_13380_));
 NAND2_X1 _39604_ (.A1(_13312_),
    .A2(_13380_),
    .ZN(_13381_));
 MUX2_X1 _39605_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [261]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [779]),
    .S(_11242_),
    .Z(_13382_));
 AND2_X1 _39606_ (.A1(_13382_),
    .A2(_11245_),
    .ZN(_13383_));
 OAI21_X1 _39607_ (.A(_13383_),
    .B1(_13343_),
    .B2(_13345_),
    .ZN(_13384_));
 AOI21_X1 _39608_ (.A(_13378_),
    .B1(_13381_),
    .B2(_13384_),
    .ZN(_13385_));
 OR2_X1 _39609_ (.A1(_13377_),
    .A2(_13385_),
    .ZN(_13386_));
 MUX2_X2 _39610_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [325]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [843]),
    .S(_11276_),
    .Z(_13387_));
 AND2_X1 _39611_ (.A1(_13387_),
    .A2(_13297_),
    .ZN(_13388_));
 NAND2_X1 _39612_ (.A1(_13254_),
    .A2(_13388_),
    .ZN(_13389_));
 MUX2_X2 _39613_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [389]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [907]),
    .S(_11276_),
    .Z(_13390_));
 AND2_X1 _39614_ (.A1(_13390_),
    .A2(_11267_),
    .ZN(_13391_));
 OAI21_X1 _39615_ (.A(_13391_),
    .B1(_13292_),
    .B2(_13293_),
    .ZN(_13392_));
 AOI21_X1 _39616_ (.A(_13222_),
    .B1(_13389_),
    .B2(_13392_),
    .ZN(_13393_));
 MUX2_X2 _39617_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [453]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [971]),
    .S(_11276_),
    .Z(_13394_));
 AND2_X1 _39618_ (.A1(_13394_),
    .A2(_11267_),
    .ZN(_13395_));
 NAND2_X1 _39619_ (.A1(_13254_),
    .A2(_13395_),
    .ZN(_13396_));
 MUX2_X2 _39620_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [517]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1035]),
    .S(_11276_),
    .Z(_13397_));
 AND2_X1 _39621_ (.A1(_13397_),
    .A2(_11267_),
    .ZN(_13398_));
 OAI21_X1 _39622_ (.A(_13398_),
    .B1(_13292_),
    .B2(_13293_),
    .ZN(_13399_));
 AOI21_X1 _39623_ (.A(_13263_),
    .B1(_13396_),
    .B2(_13399_),
    .ZN(_13400_));
 OR2_X1 _39624_ (.A1(_13393_),
    .A2(_13400_),
    .ZN(_13401_));
 MUX2_X2 _39625_ (.A(_13386_),
    .B(_13401_),
    .S(_12337_),
    .Z(\icache.data_mem_data_li [63]));
 NAND2_X1 _39626_ (.A1(_13312_),
    .A2(_11281_),
    .ZN(_13402_));
 OAI21_X1 _39627_ (.A(_11278_),
    .B1(_13343_),
    .B2(_13345_),
    .ZN(_13403_));
 AOI21_X1 _39628_ (.A(_13336_),
    .B1(_13402_),
    .B2(_13403_),
    .ZN(_13404_));
 NAND2_X1 _39629_ (.A1(_13312_),
    .A2(_11288_),
    .ZN(_13405_));
 OAI21_X1 _39630_ (.A(_11285_),
    .B1(_13343_),
    .B2(_13345_),
    .ZN(_13406_));
 AOI21_X1 _39631_ (.A(_13378_),
    .B1(_13405_),
    .B2(_13406_),
    .ZN(_13407_));
 OR2_X4 _39632_ (.A1(_13404_),
    .A2(_13407_),
    .ZN(_13408_));
 BUF_X4 _39633_ (.A(_12421_),
    .Z(_13409_));
 NAND2_X1 _39634_ (.A1(_13409_),
    .A2(_11250_),
    .ZN(_13410_));
 OAI21_X1 _39635_ (.A(_11246_),
    .B1(_13292_),
    .B2(_13293_),
    .ZN(_13411_));
 AOI21_X1 _39636_ (.A(_13222_),
    .B1(_13410_),
    .B2(_13411_),
    .ZN(_13412_));
 NAND2_X1 _39637_ (.A1(_13409_),
    .A2(_11268_),
    .ZN(_13413_));
 OAI21_X1 _39638_ (.A(_11261_),
    .B1(_13292_),
    .B2(_13293_),
    .ZN(_13414_));
 AOI21_X1 _39639_ (.A(_13263_),
    .B1(_13413_),
    .B2(_13414_),
    .ZN(_13415_));
 OR2_X4 _39640_ (.A1(_13412_),
    .A2(_13415_),
    .ZN(_13416_));
 MUX2_X2 _39641_ (.A(_13408_),
    .B(_13416_),
    .S(_13171_),
    .Z(\icache.data_mem_data_li [64]));
 NAND2_X1 _39642_ (.A1(_13409_),
    .A2(_11298_),
    .ZN(_13417_));
 BUF_X4 _39643_ (.A(_12610_),
    .Z(_13418_));
 BUF_X4 _39644_ (.A(_12612_),
    .Z(_13419_));
 OAI21_X1 _39645_ (.A(_11295_),
    .B1(_13418_),
    .B2(_13419_),
    .ZN(_13420_));
 AOI21_X1 _39646_ (.A(_13336_),
    .B1(_13417_),
    .B2(_13420_),
    .ZN(_13421_));
 NAND2_X1 _39647_ (.A1(_13312_),
    .A2(_11307_),
    .ZN(_13422_));
 OAI21_X1 _39648_ (.A(_11304_),
    .B1(_13343_),
    .B2(_13345_),
    .ZN(_13423_));
 AOI21_X1 _39649_ (.A(_13378_),
    .B1(_13422_),
    .B2(_13423_),
    .ZN(_13424_));
 OR2_X4 _39650_ (.A1(_13421_),
    .A2(_13424_),
    .ZN(_13425_));
 NAND2_X1 _39651_ (.A1(_13312_),
    .A2(_11317_),
    .ZN(_13426_));
 OAI21_X2 _39652_ (.A(_11314_),
    .B1(_13343_),
    .B2(_13345_),
    .ZN(_13427_));
 AOI21_X1 _39653_ (.A(_13222_),
    .B1(_13426_),
    .B2(_13427_),
    .ZN(_13428_));
 NAND2_X1 _39654_ (.A1(_13409_),
    .A2(_11324_),
    .ZN(_13429_));
 OAI21_X1 _39655_ (.A(_11321_),
    .B1(_13418_),
    .B2(_13419_),
    .ZN(_13430_));
 AOI21_X1 _39656_ (.A(_13263_),
    .B1(_13429_),
    .B2(_13430_),
    .ZN(_13431_));
 OR2_X4 _39657_ (.A1(_13428_),
    .A2(_13431_),
    .ZN(_13432_));
 MUX2_X2 _39658_ (.A(_13425_),
    .B(_13432_),
    .S(_13171_),
    .Z(\icache.data_mem_data_li [65]));
 BUF_X4 _39659_ (.A(_12973_),
    .Z(_13433_));
 NAND2_X1 _39660_ (.A1(_13433_),
    .A2(_11334_),
    .ZN(_13434_));
 OAI21_X1 _39661_ (.A(_11331_),
    .B1(_13343_),
    .B2(_13345_),
    .ZN(_13435_));
 AOI21_X1 _39662_ (.A(_13336_),
    .B1(_13434_),
    .B2(_13435_),
    .ZN(_13436_));
 NAND2_X1 _39663_ (.A1(_13433_),
    .A2(_11343_),
    .ZN(_13437_));
 OAI21_X1 _39664_ (.A(_11340_),
    .B1(_13343_),
    .B2(_13345_),
    .ZN(_13438_));
 AOI21_X1 _39665_ (.A(_13378_),
    .B1(_13437_),
    .B2(_13438_),
    .ZN(_13439_));
 OR2_X4 _39666_ (.A1(_13436_),
    .A2(_13439_),
    .ZN(_13440_));
 NAND2_X1 _39667_ (.A1(_13409_),
    .A2(_11352_),
    .ZN(_13441_));
 OAI21_X2 _39668_ (.A(_11349_),
    .B1(_13418_),
    .B2(_13419_),
    .ZN(_13442_));
 AOI21_X1 _39669_ (.A(_13222_),
    .B1(_13441_),
    .B2(_13442_),
    .ZN(_13443_));
 NAND2_X1 _39670_ (.A1(_13409_),
    .A2(_11360_),
    .ZN(_13444_));
 OAI21_X1 _39671_ (.A(_11356_),
    .B1(_13418_),
    .B2(_13419_),
    .ZN(_13445_));
 AOI21_X1 _39672_ (.A(_13263_),
    .B1(_13444_),
    .B2(_13445_),
    .ZN(_13446_));
 OR2_X4 _39673_ (.A1(_13443_),
    .A2(_13446_),
    .ZN(_13447_));
 MUX2_X2 _39674_ (.A(_13440_),
    .B(_13447_),
    .S(_13171_),
    .Z(\icache.data_mem_data_li [66]));
 NAND2_X1 _39675_ (.A1(_13433_),
    .A2(_11368_),
    .ZN(_13448_));
 BUF_X4 _39676_ (.A(_13342_),
    .Z(_13449_));
 BUF_X4 _39677_ (.A(_13344_),
    .Z(_13450_));
 OAI21_X1 _39678_ (.A(_11365_),
    .B1(_13449_),
    .B2(_13450_),
    .ZN(_13451_));
 AOI21_X1 _39679_ (.A(_13336_),
    .B1(_13448_),
    .B2(_13451_),
    .ZN(_13452_));
 NAND2_X1 _39680_ (.A1(_13433_),
    .A2(_11377_),
    .ZN(_13453_));
 OAI21_X1 _39681_ (.A(_11374_),
    .B1(_13449_),
    .B2(_13450_),
    .ZN(_13454_));
 AOI21_X1 _39682_ (.A(_13378_),
    .B1(_13453_),
    .B2(_13454_),
    .ZN(_13455_));
 OR2_X4 _39683_ (.A1(_13452_),
    .A2(_13455_),
    .ZN(_13456_));
 NAND2_X1 _39684_ (.A1(_13409_),
    .A2(_11385_),
    .ZN(_13457_));
 OAI21_X2 _39685_ (.A(_11382_),
    .B1(_13418_),
    .B2(_13419_),
    .ZN(_13458_));
 AOI21_X1 _39686_ (.A(_13222_),
    .B1(_13457_),
    .B2(_13458_),
    .ZN(_13459_));
 NAND2_X1 _39687_ (.A1(_13409_),
    .A2(_11392_),
    .ZN(_13460_));
 OAI21_X2 _39688_ (.A(_11389_),
    .B1(_13418_),
    .B2(_13419_),
    .ZN(_13461_));
 AOI21_X2 _39689_ (.A(_13263_),
    .B1(_13460_),
    .B2(_13461_),
    .ZN(_13462_));
 OR2_X4 _39690_ (.A1(_13459_),
    .A2(_13462_),
    .ZN(_13463_));
 BUF_X4 _39691_ (.A(_12640_),
    .Z(_13464_));
 MUX2_X2 _39692_ (.A(_13456_),
    .B(_13463_),
    .S(_13464_),
    .Z(\icache.data_mem_data_li [67]));
 NAND2_X1 _39693_ (.A1(_13409_),
    .A2(_11419_),
    .ZN(_13465_));
 OAI21_X1 _39694_ (.A(_11416_),
    .B1(_13418_),
    .B2(_13419_),
    .ZN(_13466_));
 AOI21_X1 _39695_ (.A(_13336_),
    .B1(_13465_),
    .B2(_13466_),
    .ZN(_13467_));
 NAND2_X1 _39696_ (.A1(_13433_),
    .A2(_11426_),
    .ZN(_13468_));
 OAI21_X1 _39697_ (.A(_11423_),
    .B1(_13449_),
    .B2(_13450_),
    .ZN(_13469_));
 AOI21_X1 _39698_ (.A(_13378_),
    .B1(_13468_),
    .B2(_13469_),
    .ZN(_13470_));
 OR2_X4 _39699_ (.A1(_13467_),
    .A2(_13470_),
    .ZN(_13471_));
 BUF_X16 _39700_ (.A(_08447_),
    .Z(_13472_));
 BUF_X8 _39701_ (.A(_13472_),
    .Z(_13473_));
 NAND2_X1 _39702_ (.A1(_13433_),
    .A2(_11401_),
    .ZN(_13474_));
 OAI21_X2 _39703_ (.A(_11397_),
    .B1(_13449_),
    .B2(_13450_),
    .ZN(_13475_));
 AOI21_X2 _39704_ (.A(_13473_),
    .B1(_13474_),
    .B2(_13475_),
    .ZN(_13476_));
 NAND2_X1 _39705_ (.A1(_13409_),
    .A2(_11409_),
    .ZN(_13477_));
 OAI21_X1 _39706_ (.A(_11406_),
    .B1(_13418_),
    .B2(_13419_),
    .ZN(_13478_));
 AOI21_X1 _39707_ (.A(_13263_),
    .B1(_13477_),
    .B2(_13478_),
    .ZN(_13479_));
 OR2_X4 _39708_ (.A1(_13476_),
    .A2(_13479_),
    .ZN(_13480_));
 BUF_X32 _39709_ (.A(_08432_),
    .Z(_13481_));
 BUF_X32 _39710_ (.A(_13481_),
    .Z(_13482_));
 MUX2_X2 _39711_ (.A(_13471_),
    .B(_13480_),
    .S(_13482_),
    .Z(\icache.data_mem_data_li [68]));
 BUF_X4 _39712_ (.A(_12421_),
    .Z(_13483_));
 NAND2_X2 _39713_ (.A1(_13483_),
    .A2(_11435_),
    .ZN(_13484_));
 OAI21_X1 _39714_ (.A(_11431_),
    .B1(_13418_),
    .B2(_13419_),
    .ZN(_13485_));
 AOI21_X1 _39715_ (.A(_13336_),
    .B1(_13484_),
    .B2(_13485_),
    .ZN(_13486_));
 NAND2_X1 _39716_ (.A1(_13433_),
    .A2(_11444_),
    .ZN(_13487_));
 OAI21_X1 _39717_ (.A(_11441_),
    .B1(_13449_),
    .B2(_13450_),
    .ZN(_13488_));
 AOI21_X1 _39718_ (.A(_13378_),
    .B1(_13487_),
    .B2(_13488_),
    .ZN(_13489_));
 OR2_X4 _39719_ (.A1(_13486_),
    .A2(_13489_),
    .ZN(_13490_));
 NAND2_X1 _39720_ (.A1(_13433_),
    .A2(_11453_),
    .ZN(_13491_));
 OAI21_X1 _39721_ (.A(_11450_),
    .B1(_13449_),
    .B2(_13450_),
    .ZN(_13492_));
 AOI21_X1 _39722_ (.A(_13473_),
    .B1(_13491_),
    .B2(_13492_),
    .ZN(_13493_));
 BUF_X32 _39723_ (.A(_08446_),
    .Z(_13494_));
 BUF_X8 _39724_ (.A(_13494_),
    .Z(_13495_));
 NAND2_X1 _39725_ (.A1(_13483_),
    .A2(_11460_),
    .ZN(_13496_));
 OAI21_X1 _39726_ (.A(_11457_),
    .B1(_13418_),
    .B2(_13419_),
    .ZN(_13497_));
 AOI21_X1 _39727_ (.A(_13495_),
    .B1(_13496_),
    .B2(_13497_),
    .ZN(_13498_));
 OR2_X4 _39728_ (.A1(_13493_),
    .A2(_13498_),
    .ZN(_13499_));
 MUX2_X2 _39729_ (.A(_13490_),
    .B(_13499_),
    .S(_13464_),
    .Z(\icache.data_mem_data_li [69]));
 NAND2_X1 _39730_ (.A1(_13483_),
    .A2(_11469_),
    .ZN(_13500_));
 BUF_X4 _39731_ (.A(_12610_),
    .Z(_13501_));
 BUF_X4 _39732_ (.A(_12612_),
    .Z(_13502_));
 OAI21_X1 _39733_ (.A(_11465_),
    .B1(_13501_),
    .B2(_13502_),
    .ZN(_13503_));
 AOI21_X1 _39734_ (.A(_13336_),
    .B1(_13500_),
    .B2(_13503_),
    .ZN(_13504_));
 NAND2_X1 _39735_ (.A1(_13433_),
    .A2(_11478_),
    .ZN(_13505_));
 OAI21_X1 _39736_ (.A(_11475_),
    .B1(_13449_),
    .B2(_13450_),
    .ZN(_13506_));
 AOI21_X1 _39737_ (.A(_13378_),
    .B1(_13505_),
    .B2(_13506_),
    .ZN(_13507_));
 OR2_X4 _39738_ (.A1(_13504_),
    .A2(_13507_),
    .ZN(_13508_));
 NAND2_X1 _39739_ (.A1(_13433_),
    .A2(_11486_),
    .ZN(_13509_));
 OAI21_X1 _39740_ (.A(_11483_),
    .B1(_13449_),
    .B2(_13450_),
    .ZN(_13510_));
 AOI21_X1 _39741_ (.A(_13473_),
    .B1(_13509_),
    .B2(_13510_),
    .ZN(_13511_));
 NAND2_X1 _39742_ (.A1(_13483_),
    .A2(_11493_),
    .ZN(_13512_));
 OAI21_X2 _39743_ (.A(_11490_),
    .B1(_13501_),
    .B2(_13502_),
    .ZN(_13513_));
 AOI21_X2 _39744_ (.A(_13495_),
    .B1(_13512_),
    .B2(_13513_),
    .ZN(_13514_));
 OR2_X4 _39745_ (.A1(_13511_),
    .A2(_13514_),
    .ZN(_13515_));
 MUX2_X2 _39746_ (.A(_13508_),
    .B(_13515_),
    .S(_13464_),
    .Z(\icache.data_mem_data_li [70]));
 BUF_X4 _39747_ (.A(_12973_),
    .Z(_13516_));
 NAND2_X1 _39748_ (.A1(_13516_),
    .A2(_11519_),
    .ZN(_13517_));
 OAI21_X1 _39749_ (.A(_11516_),
    .B1(_13449_),
    .B2(_13450_),
    .ZN(_13518_));
 AOI21_X1 _39750_ (.A(_13336_),
    .B1(_13517_),
    .B2(_13518_),
    .ZN(_13519_));
 NAND2_X1 _39751_ (.A1(_13516_),
    .A2(_11526_),
    .ZN(_13520_));
 OAI21_X1 _39752_ (.A(_11523_),
    .B1(_13449_),
    .B2(_13450_),
    .ZN(_13521_));
 AOI21_X1 _39753_ (.A(_13378_),
    .B1(_13520_),
    .B2(_13521_),
    .ZN(_13522_));
 OR2_X4 _39754_ (.A1(_13519_),
    .A2(_13522_),
    .ZN(_13523_));
 NAND2_X1 _39755_ (.A1(_13483_),
    .A2(_11501_),
    .ZN(_13524_));
 OAI21_X1 _39756_ (.A(_11498_),
    .B1(_13501_),
    .B2(_13502_),
    .ZN(_13525_));
 AOI21_X1 _39757_ (.A(_13473_),
    .B1(_13524_),
    .B2(_13525_),
    .ZN(_13526_));
 NAND2_X1 _39758_ (.A1(_13483_),
    .A2(_11509_),
    .ZN(_13527_));
 OAI21_X1 _39759_ (.A(_11505_),
    .B1(_13501_),
    .B2(_13502_),
    .ZN(_13528_));
 AOI21_X1 _39760_ (.A(_13495_),
    .B1(_13527_),
    .B2(_13528_),
    .ZN(_13529_));
 OR2_X4 _39761_ (.A1(_13526_),
    .A2(_13529_),
    .ZN(_13530_));
 MUX2_X2 _39762_ (.A(_13523_),
    .B(_13530_),
    .S(_13464_),
    .Z(\icache.data_mem_data_li [71]));
 BUF_X8 _39763_ (.A(_11665_),
    .Z(_13531_));
 NAND2_X1 _39764_ (.A1(_13516_),
    .A2(_11552_),
    .ZN(_13532_));
 BUF_X4 _39765_ (.A(_13342_),
    .Z(_13533_));
 BUF_X4 _39766_ (.A(_13344_),
    .Z(_13534_));
 OAI21_X2 _39767_ (.A(_11549_),
    .B1(_13533_),
    .B2(_13534_),
    .ZN(_13535_));
 AOI21_X2 _39768_ (.A(_13531_),
    .B1(_13532_),
    .B2(_13535_),
    .ZN(_13536_));
 NAND2_X1 _39769_ (.A1(_13516_),
    .A2(_11559_),
    .ZN(_13537_));
 OAI21_X1 _39770_ (.A(_11556_),
    .B1(_13533_),
    .B2(_13534_),
    .ZN(_13538_));
 AOI21_X1 _39771_ (.A(_13378_),
    .B1(_13537_),
    .B2(_13538_),
    .ZN(_13539_));
 OR2_X4 _39772_ (.A1(_13536_),
    .A2(_13539_),
    .ZN(_13540_));
 NAND2_X1 _39773_ (.A1(_13483_),
    .A2(_11535_),
    .ZN(_13541_));
 OAI21_X2 _39774_ (.A(_11531_),
    .B1(_13501_),
    .B2(_13502_),
    .ZN(_13542_));
 AOI21_X2 _39775_ (.A(_13473_),
    .B1(_13541_),
    .B2(_13542_),
    .ZN(_13543_));
 NAND2_X1 _39776_ (.A1(_13483_),
    .A2(_11542_),
    .ZN(_13544_));
 OAI21_X1 _39777_ (.A(_11539_),
    .B1(_13501_),
    .B2(_13502_),
    .ZN(_13545_));
 AOI21_X1 _39778_ (.A(_13495_),
    .B1(_13544_),
    .B2(_13545_),
    .ZN(_13546_));
 OR2_X4 _39779_ (.A1(_13543_),
    .A2(_13546_),
    .ZN(_13547_));
 MUX2_X2 _39780_ (.A(_13540_),
    .B(_13547_),
    .S(_13482_),
    .Z(\icache.data_mem_data_li [72]));
 NAND2_X1 _39781_ (.A1(_13516_),
    .A2(_11586_),
    .ZN(_13548_));
 OAI21_X1 _39782_ (.A(_11583_),
    .B1(_13533_),
    .B2(_13534_),
    .ZN(_13549_));
 AOI21_X1 _39783_ (.A(_13531_),
    .B1(_13548_),
    .B2(_13549_),
    .ZN(_13550_));
 BUF_X8 _39784_ (.A(_11709_),
    .Z(_13551_));
 NAND2_X1 _39785_ (.A1(_13516_),
    .A2(_11594_),
    .ZN(_13552_));
 OAI21_X1 _39786_ (.A(_11591_),
    .B1(_13533_),
    .B2(_13534_),
    .ZN(_13553_));
 AOI21_X1 _39787_ (.A(_13551_),
    .B1(_13552_),
    .B2(_13553_),
    .ZN(_13554_));
 OR2_X4 _39788_ (.A1(_13550_),
    .A2(_13554_),
    .ZN(_13555_));
 NAND2_X1 _39789_ (.A1(_13483_),
    .A2(_11569_),
    .ZN(_13556_));
 OAI21_X1 _39790_ (.A(_11566_),
    .B1(_13501_),
    .B2(_13502_),
    .ZN(_13557_));
 AOI21_X1 _39791_ (.A(_13473_),
    .B1(_13556_),
    .B2(_13557_),
    .ZN(_13558_));
 NAND2_X1 _39792_ (.A1(_13483_),
    .A2(_11578_),
    .ZN(_13559_));
 OAI21_X1 _39793_ (.A(_11574_),
    .B1(_13501_),
    .B2(_13502_),
    .ZN(_13560_));
 AOI21_X1 _39794_ (.A(_13495_),
    .B1(_13559_),
    .B2(_13560_),
    .ZN(_13561_));
 OR2_X4 _39795_ (.A1(_13558_),
    .A2(_13561_),
    .ZN(_13562_));
 MUX2_X2 _39796_ (.A(_13555_),
    .B(_13562_),
    .S(_13464_),
    .Z(\icache.data_mem_data_li [73]));
 NAND2_X1 _39797_ (.A1(_13516_),
    .A2(_11618_),
    .ZN(_13563_));
 OAI21_X1 _39798_ (.A(_11615_),
    .B1(_13533_),
    .B2(_13534_),
    .ZN(_13564_));
 AOI21_X1 _39799_ (.A(_13531_),
    .B1(_13563_),
    .B2(_13564_),
    .ZN(_13565_));
 NAND2_X1 _39800_ (.A1(_13516_),
    .A2(_11627_),
    .ZN(_13566_));
 OAI21_X2 _39801_ (.A(_11624_),
    .B1(_13533_),
    .B2(_13534_),
    .ZN(_13567_));
 AOI21_X1 _39802_ (.A(_13551_),
    .B1(_13566_),
    .B2(_13567_),
    .ZN(_13568_));
 OR2_X4 _39803_ (.A1(_13565_),
    .A2(_13568_),
    .ZN(_13569_));
 BUF_X4 _39804_ (.A(_12421_),
    .Z(_13570_));
 NAND2_X1 _39805_ (.A1(_13570_),
    .A2(_11603_),
    .ZN(_13571_));
 OAI21_X1 _39806_ (.A(_11599_),
    .B1(_13501_),
    .B2(_13502_),
    .ZN(_13572_));
 AOI21_X1 _39807_ (.A(_13473_),
    .B1(_13571_),
    .B2(_13572_),
    .ZN(_13573_));
 NAND2_X1 _39808_ (.A1(_13570_),
    .A2(_11610_),
    .ZN(_13574_));
 OAI21_X1 _39809_ (.A(_11607_),
    .B1(_13501_),
    .B2(_13502_),
    .ZN(_13575_));
 AOI21_X1 _39810_ (.A(_13495_),
    .B1(_13574_),
    .B2(_13575_),
    .ZN(_13576_));
 OR2_X4 _39811_ (.A1(_13573_),
    .A2(_13576_),
    .ZN(_13577_));
 MUX2_X2 _39812_ (.A(_13569_),
    .B(_13577_),
    .S(_13464_),
    .Z(\icache.data_mem_data_li [74]));
 NAND2_X1 _39813_ (.A1(_13516_),
    .A2(_11654_),
    .ZN(_13578_));
 OAI21_X1 _39814_ (.A(_11651_),
    .B1(_13533_),
    .B2(_13534_),
    .ZN(_13579_));
 AOI21_X1 _39815_ (.A(_13531_),
    .B1(_13578_),
    .B2(_13579_),
    .ZN(_13580_));
 NAND2_X1 _39816_ (.A1(_13516_),
    .A2(_11661_),
    .ZN(_13581_));
 OAI21_X1 _39817_ (.A(_11658_),
    .B1(_13533_),
    .B2(_13534_),
    .ZN(_13582_));
 AOI21_X1 _39818_ (.A(_13551_),
    .B1(_13581_),
    .B2(_13582_),
    .ZN(_13583_));
 OR2_X4 _39819_ (.A1(_13580_),
    .A2(_13583_),
    .ZN(_13584_));
 NAND2_X1 _39820_ (.A1(_13570_),
    .A2(_11635_),
    .ZN(_13585_));
 BUF_X4 _39821_ (.A(_12610_),
    .Z(_13586_));
 BUF_X4 _39822_ (.A(_12612_),
    .Z(_13587_));
 OAI21_X1 _39823_ (.A(_11632_),
    .B1(_13586_),
    .B2(_13587_),
    .ZN(_13588_));
 AOI21_X1 _39824_ (.A(_13473_),
    .B1(_13585_),
    .B2(_13588_),
    .ZN(_13589_));
 NAND2_X1 _39825_ (.A1(_13570_),
    .A2(_11646_),
    .ZN(_13590_));
 OAI21_X1 _39826_ (.A(_11641_),
    .B1(_13586_),
    .B2(_13587_),
    .ZN(_13591_));
 AOI21_X1 _39827_ (.A(_13495_),
    .B1(_13590_),
    .B2(_13591_),
    .ZN(_13592_));
 OR2_X4 _39828_ (.A1(_13589_),
    .A2(_13592_),
    .ZN(_13593_));
 MUX2_X2 _39829_ (.A(_13584_),
    .B(_13593_),
    .S(_13464_),
    .Z(\icache.data_mem_data_li [75]));
 NAND2_X1 _39830_ (.A1(_13570_),
    .A2(_11672_),
    .ZN(_13594_));
 OAI21_X1 _39831_ (.A(_11668_),
    .B1(_13586_),
    .B2(_13587_),
    .ZN(_13595_));
 AOI21_X1 _39832_ (.A(_13531_),
    .B1(_13594_),
    .B2(_13595_),
    .ZN(_13596_));
 BUF_X4 _39833_ (.A(_12973_),
    .Z(_13597_));
 NAND2_X1 _39834_ (.A1(_13597_),
    .A2(_11679_),
    .ZN(_13598_));
 OAI21_X1 _39835_ (.A(_11676_),
    .B1(_13533_),
    .B2(_13534_),
    .ZN(_13599_));
 AOI21_X1 _39836_ (.A(_13551_),
    .B1(_13598_),
    .B2(_13599_),
    .ZN(_13600_));
 OR2_X4 _39837_ (.A1(_13596_),
    .A2(_13600_),
    .ZN(_13601_));
 NAND2_X1 _39838_ (.A1(_13597_),
    .A2(_11691_),
    .ZN(_13602_));
 OAI21_X1 _39839_ (.A(_11688_),
    .B1(_13533_),
    .B2(_13534_),
    .ZN(_13603_));
 AOI21_X1 _39840_ (.A(_13473_),
    .B1(_13602_),
    .B2(_13603_),
    .ZN(_13604_));
 NAND2_X1 _39841_ (.A1(_13570_),
    .A2(_11698_),
    .ZN(_13605_));
 OAI21_X1 _39842_ (.A(_11695_),
    .B1(_13586_),
    .B2(_13587_),
    .ZN(_13606_));
 AOI21_X1 _39843_ (.A(_13495_),
    .B1(_13605_),
    .B2(_13606_),
    .ZN(_13607_));
 OR2_X4 _39844_ (.A1(_13604_),
    .A2(_13607_),
    .ZN(_13608_));
 MUX2_X2 _39845_ (.A(_13601_),
    .B(_13608_),
    .S(_13464_),
    .Z(\icache.data_mem_data_li [76]));
 NAND2_X1 _39846_ (.A1(_13570_),
    .A2(_11706_),
    .ZN(_13609_));
 OAI21_X1 _39847_ (.A(_11703_),
    .B1(_13586_),
    .B2(_13587_),
    .ZN(_13610_));
 AOI21_X1 _39848_ (.A(_13531_),
    .B1(_13609_),
    .B2(_13610_),
    .ZN(_13611_));
 NAND2_X1 _39849_ (.A1(_13597_),
    .A2(_11716_),
    .ZN(_13612_));
 BUF_X4 _39850_ (.A(_13342_),
    .Z(_13613_));
 BUF_X4 _39851_ (.A(_13344_),
    .Z(_13614_));
 OAI21_X1 _39852_ (.A(_11713_),
    .B1(_13613_),
    .B2(_13614_),
    .ZN(_13615_));
 AOI21_X1 _39853_ (.A(_13551_),
    .B1(_13612_),
    .B2(_13615_),
    .ZN(_13616_));
 OR2_X4 _39854_ (.A1(_13611_),
    .A2(_13616_),
    .ZN(_13617_));
 NAND2_X1 _39855_ (.A1(_13597_),
    .A2(_11725_),
    .ZN(_13618_));
 OAI21_X2 _39856_ (.A(_11722_),
    .B1(_13613_),
    .B2(_13614_),
    .ZN(_13619_));
 AOI21_X1 _39857_ (.A(_13473_),
    .B1(_13618_),
    .B2(_13619_),
    .ZN(_13620_));
 NAND2_X1 _39858_ (.A1(_13570_),
    .A2(_11732_),
    .ZN(_13621_));
 OAI21_X1 _39859_ (.A(_11729_),
    .B1(_13586_),
    .B2(_13587_),
    .ZN(_13622_));
 AOI21_X1 _39860_ (.A(_13495_),
    .B1(_13621_),
    .B2(_13622_),
    .ZN(_13623_));
 OR2_X4 _39861_ (.A1(_13620_),
    .A2(_13623_),
    .ZN(_13624_));
 MUX2_X2 _39862_ (.A(_13617_),
    .B(_13624_),
    .S(_13464_),
    .Z(\icache.data_mem_data_li [77]));
 NAND2_X1 _39863_ (.A1(_13570_),
    .A2(_11758_),
    .ZN(_13625_));
 OAI21_X1 _39864_ (.A(_11755_),
    .B1(_13586_),
    .B2(_13587_),
    .ZN(_13626_));
 AOI21_X1 _39865_ (.A(_13531_),
    .B1(_13625_),
    .B2(_13626_),
    .ZN(_13627_));
 NAND2_X1 _39866_ (.A1(_13597_),
    .A2(_11765_),
    .ZN(_13628_));
 OAI21_X2 _39867_ (.A(_11762_),
    .B1(_13613_),
    .B2(_13614_),
    .ZN(_13629_));
 AOI21_X1 _39868_ (.A(_13551_),
    .B1(_13628_),
    .B2(_13629_),
    .ZN(_13630_));
 OR2_X4 _39869_ (.A1(_13627_),
    .A2(_13630_),
    .ZN(_13631_));
 BUF_X8 _39870_ (.A(_13472_),
    .Z(_13632_));
 NAND2_X1 _39871_ (.A1(_13597_),
    .A2(_11740_),
    .ZN(_13633_));
 OAI21_X1 _39872_ (.A(_11737_),
    .B1(_13613_),
    .B2(_13614_),
    .ZN(_13634_));
 AOI21_X1 _39873_ (.A(_13632_),
    .B1(_13633_),
    .B2(_13634_),
    .ZN(_13635_));
 NAND2_X1 _39874_ (.A1(_13570_),
    .A2(_11749_),
    .ZN(_13636_));
 OAI21_X1 _39875_ (.A(_11745_),
    .B1(_13586_),
    .B2(_13587_),
    .ZN(_13637_));
 AOI21_X1 _39876_ (.A(_13495_),
    .B1(_13636_),
    .B2(_13637_),
    .ZN(_13638_));
 OR2_X4 _39877_ (.A1(_13635_),
    .A2(_13638_),
    .ZN(_13639_));
 MUX2_X2 _39878_ (.A(_13631_),
    .B(_13639_),
    .S(_13482_),
    .Z(\icache.data_mem_data_li [78]));
 NAND2_X1 _39879_ (.A1(_13597_),
    .A2(_11792_),
    .ZN(_13640_));
 OAI21_X1 _39880_ (.A(_11789_),
    .B1(_13613_),
    .B2(_13614_),
    .ZN(_13641_));
 AOI21_X1 _39881_ (.A(_13531_),
    .B1(_13640_),
    .B2(_13641_),
    .ZN(_13642_));
 NAND2_X1 _39882_ (.A1(_13597_),
    .A2(_11799_),
    .ZN(_13643_));
 OAI21_X1 _39883_ (.A(_11796_),
    .B1(_13613_),
    .B2(_13614_),
    .ZN(_13644_));
 AOI21_X1 _39884_ (.A(_13551_),
    .B1(_13643_),
    .B2(_13644_),
    .ZN(_13645_));
 OR2_X4 _39885_ (.A1(_13642_),
    .A2(_13645_),
    .ZN(_13646_));
 BUF_X4 _39886_ (.A(_12421_),
    .Z(_13647_));
 NAND2_X1 _39887_ (.A1(_13647_),
    .A2(_11775_),
    .ZN(_13648_));
 OAI21_X2 _39888_ (.A(_11771_),
    .B1(_13586_),
    .B2(_13587_),
    .ZN(_13649_));
 AOI21_X1 _39889_ (.A(_13632_),
    .B1(_13648_),
    .B2(_13649_),
    .ZN(_13650_));
 BUF_X8 _39890_ (.A(_13494_),
    .Z(_13651_));
 NAND2_X1 _39891_ (.A1(_13647_),
    .A2(_11784_),
    .ZN(_13652_));
 OAI21_X2 _39892_ (.A(_11781_),
    .B1(_13586_),
    .B2(_13587_),
    .ZN(_13653_));
 AOI21_X1 _39893_ (.A(_13651_),
    .B1(_13652_),
    .B2(_13653_),
    .ZN(_13654_));
 OR2_X4 _39894_ (.A1(_13650_),
    .A2(_13654_),
    .ZN(_13655_));
 MUX2_X2 _39895_ (.A(_13646_),
    .B(_13655_),
    .S(_13482_),
    .Z(\icache.data_mem_data_li [79]));
 NAND2_X1 _39896_ (.A1(_13647_),
    .A2(_11807_),
    .ZN(_13656_));
 BUF_X4 _39897_ (.A(_12610_),
    .Z(_13657_));
 BUF_X4 _39898_ (.A(_12612_),
    .Z(_13658_));
 OAI21_X1 _39899_ (.A(_11804_),
    .B1(_13657_),
    .B2(_13658_),
    .ZN(_13659_));
 AOI21_X1 _39900_ (.A(_13531_),
    .B1(_13656_),
    .B2(_13659_),
    .ZN(_13660_));
 NAND2_X1 _39901_ (.A1(_13597_),
    .A2(_11816_),
    .ZN(_13661_));
 OAI21_X1 _39902_ (.A(_11813_),
    .B1(_13613_),
    .B2(_13614_),
    .ZN(_13662_));
 AOI21_X1 _39903_ (.A(_13551_),
    .B1(_13661_),
    .B2(_13662_),
    .ZN(_13663_));
 OR2_X4 _39904_ (.A1(_13660_),
    .A2(_13663_),
    .ZN(_13664_));
 NAND2_X1 _39905_ (.A1(_13597_),
    .A2(_11824_),
    .ZN(_13665_));
 OAI21_X1 _39906_ (.A(_11821_),
    .B1(_13613_),
    .B2(_13614_),
    .ZN(_13666_));
 AOI21_X1 _39907_ (.A(_13632_),
    .B1(_13665_),
    .B2(_13666_),
    .ZN(_13667_));
 NAND2_X1 _39908_ (.A1(_13647_),
    .A2(_11831_),
    .ZN(_13668_));
 OAI21_X1 _39909_ (.A(_11828_),
    .B1(_13657_),
    .B2(_13658_),
    .ZN(_13669_));
 AOI21_X1 _39910_ (.A(_13651_),
    .B1(_13668_),
    .B2(_13669_),
    .ZN(_13670_));
 OR2_X4 _39911_ (.A1(_13667_),
    .A2(_13670_),
    .ZN(_13671_));
 MUX2_X2 _39912_ (.A(_13664_),
    .B(_13671_),
    .S(_13482_),
    .Z(\icache.data_mem_data_li [80]));
 NAND2_X1 _39913_ (.A1(_13647_),
    .A2(_11841_),
    .ZN(_13672_));
 OAI21_X1 _39914_ (.A(_11838_),
    .B1(_13657_),
    .B2(_13658_),
    .ZN(_13673_));
 AOI21_X1 _39915_ (.A(_13531_),
    .B1(_13672_),
    .B2(_13673_),
    .ZN(_13674_));
 BUF_X4 _39916_ (.A(_12973_),
    .Z(_13675_));
 NAND2_X1 _39917_ (.A1(_13675_),
    .A2(_11849_),
    .ZN(_13676_));
 OAI21_X2 _39918_ (.A(_11845_),
    .B1(_13613_),
    .B2(_13614_),
    .ZN(_13677_));
 AOI21_X1 _39919_ (.A(_13551_),
    .B1(_13676_),
    .B2(_13677_),
    .ZN(_13678_));
 OR2_X4 _39920_ (.A1(_13674_),
    .A2(_13678_),
    .ZN(_13679_));
 NAND2_X2 _39921_ (.A1(_13675_),
    .A2(_11859_),
    .ZN(_13680_));
 OAI21_X1 _39922_ (.A(_11856_),
    .B1(_13613_),
    .B2(_13614_),
    .ZN(_13681_));
 AOI21_X1 _39923_ (.A(_13632_),
    .B1(_13680_),
    .B2(_13681_),
    .ZN(_13682_));
 NAND2_X1 _39924_ (.A1(_13647_),
    .A2(_11866_),
    .ZN(_13683_));
 OAI21_X1 _39925_ (.A(_11863_),
    .B1(_13657_),
    .B2(_13658_),
    .ZN(_13684_));
 AOI21_X1 _39926_ (.A(_13651_),
    .B1(_13683_),
    .B2(_13684_),
    .ZN(_13685_));
 OR2_X4 _39927_ (.A1(_13682_),
    .A2(_13685_),
    .ZN(_13686_));
 MUX2_X2 _39928_ (.A(_13679_),
    .B(_13686_),
    .S(_13464_),
    .Z(\icache.data_mem_data_li [81]));
 BUF_X8 _39929_ (.A(_11665_),
    .Z(_13687_));
 NAND2_X1 _39930_ (.A1(_13675_),
    .A2(_11874_),
    .ZN(_13688_));
 BUF_X4 _39931_ (.A(_13342_),
    .Z(_13689_));
 BUF_X4 _39932_ (.A(_13344_),
    .Z(_13690_));
 OAI21_X1 _39933_ (.A(_11871_),
    .B1(_13689_),
    .B2(_13690_),
    .ZN(_13691_));
 AOI21_X1 _39934_ (.A(_13687_),
    .B1(_13688_),
    .B2(_13691_),
    .ZN(_13692_));
 NAND2_X1 _39935_ (.A1(_13675_),
    .A2(_11882_),
    .ZN(_13693_));
 OAI21_X1 _39936_ (.A(_11878_),
    .B1(_13689_),
    .B2(_13690_),
    .ZN(_13694_));
 AOI21_X1 _39937_ (.A(_13551_),
    .B1(_13693_),
    .B2(_13694_),
    .ZN(_13695_));
 OR2_X4 _39938_ (.A1(_13692_),
    .A2(_13695_),
    .ZN(_13696_));
 NAND2_X1 _39939_ (.A1(_13647_),
    .A2(_11891_),
    .ZN(_13697_));
 OAI21_X1 _39940_ (.A(_11888_),
    .B1(_13657_),
    .B2(_13658_),
    .ZN(_13698_));
 AOI21_X1 _39941_ (.A(_13632_),
    .B1(_13697_),
    .B2(_13698_),
    .ZN(_13699_));
 NAND2_X1 _39942_ (.A1(_13647_),
    .A2(_11899_),
    .ZN(_13700_));
 OAI21_X1 _39943_ (.A(_11896_),
    .B1(_13657_),
    .B2(_13658_),
    .ZN(_13701_));
 AOI21_X1 _39944_ (.A(_13651_),
    .B1(_13700_),
    .B2(_13701_),
    .ZN(_13702_));
 OR2_X4 _39945_ (.A1(_13699_),
    .A2(_13702_),
    .ZN(_13703_));
 BUF_X4 _39946_ (.A(_12640_),
    .Z(_13704_));
 MUX2_X2 _39947_ (.A(_13696_),
    .B(_13703_),
    .S(_13704_),
    .Z(\icache.data_mem_data_li [82]));
 NAND2_X1 _39948_ (.A1(_13675_),
    .A2(_11907_),
    .ZN(_13705_));
 OAI21_X1 _39949_ (.A(_11904_),
    .B1(_13689_),
    .B2(_13690_),
    .ZN(_13706_));
 AOI21_X1 _39950_ (.A(_13687_),
    .B1(_13705_),
    .B2(_13706_),
    .ZN(_13707_));
 BUF_X8 _39951_ (.A(_11709_),
    .Z(_13708_));
 NAND2_X1 _39952_ (.A1(_13675_),
    .A2(_11914_),
    .ZN(_13709_));
 OAI21_X1 _39953_ (.A(_11911_),
    .B1(_13689_),
    .B2(_13690_),
    .ZN(_13710_));
 AOI21_X1 _39954_ (.A(_13708_),
    .B1(_13709_),
    .B2(_13710_),
    .ZN(_13711_));
 OR2_X4 _39955_ (.A1(_13707_),
    .A2(_13711_),
    .ZN(_13712_));
 NAND2_X1 _39956_ (.A1(_13647_),
    .A2(_11924_),
    .ZN(_13713_));
 OAI21_X1 _39957_ (.A(_11921_),
    .B1(_13657_),
    .B2(_13658_),
    .ZN(_13714_));
 AOI21_X1 _39958_ (.A(_13632_),
    .B1(_13713_),
    .B2(_13714_),
    .ZN(_13715_));
 NAND2_X1 _39959_ (.A1(_13647_),
    .A2(_11932_),
    .ZN(_13716_));
 OAI21_X1 _39960_ (.A(_11929_),
    .B1(_13657_),
    .B2(_13658_),
    .ZN(_13717_));
 AOI21_X1 _39961_ (.A(_13651_),
    .B1(_13716_),
    .B2(_13717_),
    .ZN(_13718_));
 OR2_X4 _39962_ (.A1(_13715_),
    .A2(_13718_),
    .ZN(_13719_));
 MUX2_X2 _39963_ (.A(_13712_),
    .B(_13719_),
    .S(_13704_),
    .Z(\icache.data_mem_data_li [83]));
 BUF_X4 _39964_ (.A(_08490_),
    .Z(_13720_));
 NAND2_X1 _39965_ (.A1(_13720_),
    .A2(_11941_),
    .ZN(_13721_));
 OAI21_X1 _39966_ (.A(_11937_),
    .B1(_13657_),
    .B2(_13658_),
    .ZN(_13722_));
 AOI21_X1 _39967_ (.A(_13687_),
    .B1(_13721_),
    .B2(_13722_),
    .ZN(_13723_));
 NAND2_X1 _39968_ (.A1(_13675_),
    .A2(_11951_),
    .ZN(_13724_));
 OAI21_X1 _39969_ (.A(_11948_),
    .B1(_13689_),
    .B2(_13690_),
    .ZN(_13725_));
 AOI21_X1 _39970_ (.A(_13708_),
    .B1(_13724_),
    .B2(_13725_),
    .ZN(_13726_));
 OR2_X4 _39971_ (.A1(_13723_),
    .A2(_13726_),
    .ZN(_13727_));
 NAND2_X2 _39972_ (.A1(_13675_),
    .A2(_11959_),
    .ZN(_13728_));
 OAI21_X2 _39973_ (.A(_11956_),
    .B1(_13689_),
    .B2(_13690_),
    .ZN(_13729_));
 AOI21_X2 _39974_ (.A(_13632_),
    .B1(_13728_),
    .B2(_13729_),
    .ZN(_13730_));
 NAND2_X1 _39975_ (.A1(_13720_),
    .A2(_11966_),
    .ZN(_13731_));
 OAI21_X2 _39976_ (.A(_11963_),
    .B1(_13657_),
    .B2(_13658_),
    .ZN(_13732_));
 AOI21_X1 _39977_ (.A(_13651_),
    .B1(_13731_),
    .B2(_13732_),
    .ZN(_13733_));
 OR2_X4 _39978_ (.A1(_13730_),
    .A2(_13733_),
    .ZN(_13734_));
 MUX2_X2 _39979_ (.A(_13727_),
    .B(_13734_),
    .S(_13482_),
    .Z(\icache.data_mem_data_li [84]));
 NAND2_X1 _39980_ (.A1(_13675_),
    .A2(_11976_),
    .ZN(_13735_));
 OAI21_X1 _39981_ (.A(_11972_),
    .B1(_13689_),
    .B2(_13690_),
    .ZN(_13736_));
 AOI21_X1 _39982_ (.A(_13687_),
    .B1(_13735_),
    .B2(_13736_),
    .ZN(_13737_));
 NAND2_X1 _39983_ (.A1(_13675_),
    .A2(_11983_),
    .ZN(_13738_));
 OAI21_X1 _39984_ (.A(_11980_),
    .B1(_13689_),
    .B2(_13690_),
    .ZN(_13739_));
 AOI21_X1 _39985_ (.A(_13708_),
    .B1(_13738_),
    .B2(_13739_),
    .ZN(_13740_));
 OR2_X4 _39986_ (.A1(_13737_),
    .A2(_13740_),
    .ZN(_13741_));
 NAND2_X1 _39987_ (.A1(_13720_),
    .A2(_11991_),
    .ZN(_13742_));
 BUF_X4 _39988_ (.A(_12610_),
    .Z(_13743_));
 BUF_X4 _39989_ (.A(_12612_),
    .Z(_13744_));
 OAI21_X1 _39990_ (.A(_11988_),
    .B1(_13743_),
    .B2(_13744_),
    .ZN(_13745_));
 AOI21_X1 _39991_ (.A(_13632_),
    .B1(_13742_),
    .B2(_13745_),
    .ZN(_13746_));
 NAND2_X1 _39992_ (.A1(_13720_),
    .A2(_11999_),
    .ZN(_13747_));
 OAI21_X1 _39993_ (.A(_11995_),
    .B1(_13743_),
    .B2(_13744_),
    .ZN(_13748_));
 AOI21_X1 _39994_ (.A(_13651_),
    .B1(_13747_),
    .B2(_13748_),
    .ZN(_13749_));
 OR2_X4 _39995_ (.A1(_13746_),
    .A2(_13749_),
    .ZN(_13750_));
 MUX2_X2 _39996_ (.A(_13741_),
    .B(_13750_),
    .S(_13704_),
    .Z(\icache.data_mem_data_li [85]));
 NAND2_X1 _39997_ (.A1(_13720_),
    .A2(_12025_),
    .ZN(_13751_));
 OAI21_X1 _39998_ (.A(_12022_),
    .B1(_13743_),
    .B2(_13744_),
    .ZN(_13752_));
 AOI21_X1 _39999_ (.A(_13687_),
    .B1(_13751_),
    .B2(_13752_),
    .ZN(_13753_));
 BUF_X4 _40000_ (.A(_12973_),
    .Z(_13754_));
 NAND2_X1 _40001_ (.A1(_13754_),
    .A2(_12032_),
    .ZN(_13755_));
 OAI21_X1 _40002_ (.A(_12029_),
    .B1(_13689_),
    .B2(_13690_),
    .ZN(_13756_));
 AOI21_X1 _40003_ (.A(_13708_),
    .B1(_13755_),
    .B2(_13756_),
    .ZN(_13757_));
 OR2_X4 _40004_ (.A1(_13753_),
    .A2(_13757_),
    .ZN(_13758_));
 NAND2_X1 _40005_ (.A1(_13754_),
    .A2(_12008_),
    .ZN(_13759_));
 OAI21_X2 _40006_ (.A(_12005_),
    .B1(_13689_),
    .B2(_13690_),
    .ZN(_13760_));
 AOI21_X2 _40007_ (.A(_13632_),
    .B1(_13759_),
    .B2(_13760_),
    .ZN(_13761_));
 NAND2_X1 _40008_ (.A1(_13720_),
    .A2(_12017_),
    .ZN(_13762_));
 OAI21_X1 _40009_ (.A(_12014_),
    .B1(_13743_),
    .B2(_13744_),
    .ZN(_13763_));
 AOI21_X1 _40010_ (.A(_13651_),
    .B1(_13762_),
    .B2(_13763_),
    .ZN(_13764_));
 OR2_X4 _40011_ (.A1(_13761_),
    .A2(_13764_),
    .ZN(_13765_));
 MUX2_X2 _40012_ (.A(_13758_),
    .B(_13765_),
    .S(_13704_),
    .Z(\icache.data_mem_data_li [86]));
 NAND2_X1 _40013_ (.A1(_13754_),
    .A2(_12041_),
    .ZN(_13766_));
 BUF_X4 _40014_ (.A(_13342_),
    .Z(_13767_));
 BUF_X4 _40015_ (.A(_13344_),
    .Z(_13768_));
 OAI21_X1 _40016_ (.A(_12038_),
    .B1(_13767_),
    .B2(_13768_),
    .ZN(_13769_));
 AOI21_X1 _40017_ (.A(_13687_),
    .B1(_13766_),
    .B2(_13769_),
    .ZN(_13770_));
 NAND2_X1 _40018_ (.A1(_13754_),
    .A2(_12049_),
    .ZN(_13771_));
 OAI21_X1 _40019_ (.A(_12046_),
    .B1(_13767_),
    .B2(_13768_),
    .ZN(_13772_));
 AOI21_X1 _40020_ (.A(_13708_),
    .B1(_13771_),
    .B2(_13772_),
    .ZN(_13773_));
 OR2_X4 _40021_ (.A1(_13770_),
    .A2(_13773_),
    .ZN(_13774_));
 NAND2_X1 _40022_ (.A1(_13720_),
    .A2(_12057_),
    .ZN(_13775_));
 OAI21_X1 _40023_ (.A(_12054_),
    .B1(_13743_),
    .B2(_13744_),
    .ZN(_13776_));
 AOI21_X2 _40024_ (.A(_13632_),
    .B1(_13775_),
    .B2(_13776_),
    .ZN(_13777_));
 NAND2_X1 _40025_ (.A1(_13720_),
    .A2(_12065_),
    .ZN(_13778_));
 OAI21_X1 _40026_ (.A(_12062_),
    .B1(_13743_),
    .B2(_13744_),
    .ZN(_13779_));
 AOI21_X1 _40027_ (.A(_13651_),
    .B1(_13778_),
    .B2(_13779_),
    .ZN(_13780_));
 OR2_X4 _40028_ (.A1(_13777_),
    .A2(_13780_),
    .ZN(_13781_));
 MUX2_X2 _40029_ (.A(_13774_),
    .B(_13781_),
    .S(_13704_),
    .Z(\icache.data_mem_data_li [87]));
 NAND2_X1 _40030_ (.A1(_13720_),
    .A2(_12075_),
    .ZN(_13782_));
 OAI21_X1 _40031_ (.A(_12072_),
    .B1(_13743_),
    .B2(_13744_),
    .ZN(_13783_));
 AOI21_X1 _40032_ (.A(_13687_),
    .B1(_13782_),
    .B2(_13783_),
    .ZN(_13784_));
 NAND2_X1 _40033_ (.A1(_13754_),
    .A2(_12084_),
    .ZN(_13785_));
 OAI21_X1 _40034_ (.A(_12081_),
    .B1(_13767_),
    .B2(_13768_),
    .ZN(_13786_));
 AOI21_X1 _40035_ (.A(_13708_),
    .B1(_13785_),
    .B2(_13786_),
    .ZN(_13787_));
 OR2_X4 _40036_ (.A1(_13784_),
    .A2(_13787_),
    .ZN(_13788_));
 BUF_X8 _40037_ (.A(_13472_),
    .Z(_13789_));
 NAND2_X1 _40038_ (.A1(_13754_),
    .A2(_12092_),
    .ZN(_13790_));
 OAI21_X1 _40039_ (.A(_12089_),
    .B1(_13767_),
    .B2(_13768_),
    .ZN(_13791_));
 AOI21_X1 _40040_ (.A(_13789_),
    .B1(_13790_),
    .B2(_13791_),
    .ZN(_13792_));
 NAND2_X1 _40041_ (.A1(_13720_),
    .A2(_12099_),
    .ZN(_13793_));
 OAI21_X1 _40042_ (.A(_12096_),
    .B1(_13743_),
    .B2(_13744_),
    .ZN(_13794_));
 AOI21_X1 _40043_ (.A(_13651_),
    .B1(_13793_),
    .B2(_13794_),
    .ZN(_13795_));
 OR2_X4 _40044_ (.A1(_13792_),
    .A2(_13795_),
    .ZN(_13796_));
 MUX2_X2 _40045_ (.A(_13788_),
    .B(_13796_),
    .S(_13704_),
    .Z(\icache.data_mem_data_li [88]));
 BUF_X4 _40046_ (.A(_08490_),
    .Z(_13797_));
 NAND2_X1 _40047_ (.A1(_13797_),
    .A2(_12124_),
    .ZN(_13798_));
 OAI21_X2 _40048_ (.A(_12121_),
    .B1(_13743_),
    .B2(_13744_),
    .ZN(_13799_));
 AOI21_X2 _40049_ (.A(_13687_),
    .B1(_13798_),
    .B2(_13799_),
    .ZN(_13800_));
 NAND2_X1 _40050_ (.A1(_13754_),
    .A2(_12133_),
    .ZN(_13801_));
 OAI21_X1 _40051_ (.A(_12130_),
    .B1(_13767_),
    .B2(_13768_),
    .ZN(_13802_));
 AOI21_X1 _40052_ (.A(_13708_),
    .B1(_13801_),
    .B2(_13802_),
    .ZN(_13803_));
 OR2_X4 _40053_ (.A1(_13800_),
    .A2(_13803_),
    .ZN(_13804_));
 NAND2_X1 _40054_ (.A1(_13754_),
    .A2(_12107_),
    .ZN(_13805_));
 OAI21_X1 _40055_ (.A(_12104_),
    .B1(_13767_),
    .B2(_13768_),
    .ZN(_13806_));
 AOI21_X1 _40056_ (.A(_13789_),
    .B1(_13805_),
    .B2(_13806_),
    .ZN(_13807_));
 BUF_X8 _40057_ (.A(_13494_),
    .Z(_13808_));
 NAND2_X1 _40058_ (.A1(_13797_),
    .A2(_12115_),
    .ZN(_13809_));
 OAI21_X1 _40059_ (.A(_12111_),
    .B1(_13743_),
    .B2(_13744_),
    .ZN(_13810_));
 AOI21_X1 _40060_ (.A(_13808_),
    .B1(_13809_),
    .B2(_13810_),
    .ZN(_13811_));
 OR2_X4 _40061_ (.A1(_13807_),
    .A2(_13811_),
    .ZN(_13812_));
 MUX2_X2 _40062_ (.A(_13804_),
    .B(_13812_),
    .S(_13482_),
    .Z(\icache.data_mem_data_li [89]));
 NAND2_X1 _40063_ (.A1(_13797_),
    .A2(_12159_),
    .ZN(_13813_));
 BUF_X4 _40064_ (.A(_11269_),
    .Z(_13814_));
 BUF_X4 _40065_ (.A(_11271_),
    .Z(_13815_));
 OAI21_X1 _40066_ (.A(_12156_),
    .B1(_13814_),
    .B2(_13815_),
    .ZN(_13816_));
 AOI21_X1 _40067_ (.A(_13687_),
    .B1(_13813_),
    .B2(_13816_),
    .ZN(_13817_));
 NAND2_X1 _40068_ (.A1(_13754_),
    .A2(_12166_),
    .ZN(_13818_));
 OAI21_X2 _40069_ (.A(_12163_),
    .B1(_13767_),
    .B2(_13768_),
    .ZN(_13819_));
 AOI21_X1 _40070_ (.A(_13708_),
    .B1(_13818_),
    .B2(_13819_),
    .ZN(_13820_));
 OR2_X4 _40071_ (.A1(_13817_),
    .A2(_13820_),
    .ZN(_13821_));
 NAND2_X1 _40072_ (.A1(_13754_),
    .A2(_12142_),
    .ZN(_13822_));
 OAI21_X2 _40073_ (.A(_12139_),
    .B1(_13767_),
    .B2(_13768_),
    .ZN(_13823_));
 AOI21_X2 _40074_ (.A(_13789_),
    .B1(_13822_),
    .B2(_13823_),
    .ZN(_13824_));
 NAND2_X1 _40075_ (.A1(_13797_),
    .A2(_12151_),
    .ZN(_13825_));
 OAI21_X1 _40076_ (.A(_12147_),
    .B1(_13814_),
    .B2(_13815_),
    .ZN(_13826_));
 AOI21_X1 _40077_ (.A(_13808_),
    .B1(_13825_),
    .B2(_13826_),
    .ZN(_13827_));
 OR2_X4 _40078_ (.A1(_13824_),
    .A2(_13827_),
    .ZN(_13828_));
 MUX2_X2 _40079_ (.A(_13821_),
    .B(_13828_),
    .S(_13482_),
    .Z(\icache.data_mem_data_li [90]));
 BUF_X4 _40080_ (.A(_12973_),
    .Z(_13829_));
 NAND2_X1 _40081_ (.A1(_13829_),
    .A2(_12174_),
    .ZN(_13830_));
 OAI21_X1 _40082_ (.A(_12171_),
    .B1(_13767_),
    .B2(_13768_),
    .ZN(_13831_));
 AOI21_X1 _40083_ (.A(_13687_),
    .B1(_13830_),
    .B2(_13831_),
    .ZN(_13832_));
 NAND2_X1 _40084_ (.A1(_13829_),
    .A2(_12183_),
    .ZN(_13833_));
 OAI21_X1 _40085_ (.A(_12180_),
    .B1(_13767_),
    .B2(_13768_),
    .ZN(_13834_));
 AOI21_X1 _40086_ (.A(_13708_),
    .B1(_13833_),
    .B2(_13834_),
    .ZN(_13835_));
 OR2_X4 _40087_ (.A1(_13832_),
    .A2(_13835_),
    .ZN(_13836_));
 NAND2_X2 _40088_ (.A1(_13797_),
    .A2(_12191_),
    .ZN(_13837_));
 OAI21_X1 _40089_ (.A(_12188_),
    .B1(_13814_),
    .B2(_13815_),
    .ZN(_13838_));
 AOI21_X1 _40090_ (.A(_13789_),
    .B1(_13837_),
    .B2(_13838_),
    .ZN(_13839_));
 NAND2_X2 _40091_ (.A1(_13797_),
    .A2(_12199_),
    .ZN(_13840_));
 OAI21_X1 _40092_ (.A(_12195_),
    .B1(_13814_),
    .B2(_13815_),
    .ZN(_13841_));
 AOI21_X1 _40093_ (.A(_13808_),
    .B1(_13840_),
    .B2(_13841_),
    .ZN(_13842_));
 OR2_X4 _40094_ (.A1(_13839_),
    .A2(_13842_),
    .ZN(_13843_));
 MUX2_X2 _40095_ (.A(_13836_),
    .B(_13843_),
    .S(_13704_),
    .Z(\icache.data_mem_data_li [91]));
 BUF_X8 _40096_ (.A(_11665_),
    .Z(_13844_));
 NAND2_X1 _40097_ (.A1(_13829_),
    .A2(_12209_),
    .ZN(_13845_));
 BUF_X4 _40098_ (.A(_13342_),
    .Z(_13846_));
 BUF_X4 _40099_ (.A(_13344_),
    .Z(_13847_));
 OAI21_X1 _40100_ (.A(_12205_),
    .B1(_13846_),
    .B2(_13847_),
    .ZN(_13848_));
 AOI21_X1 _40101_ (.A(_13844_),
    .B1(_13845_),
    .B2(_13848_),
    .ZN(_13849_));
 NAND2_X1 _40102_ (.A1(_13829_),
    .A2(_12216_),
    .ZN(_13850_));
 OAI21_X1 _40103_ (.A(_12213_),
    .B1(_13846_),
    .B2(_13847_),
    .ZN(_13851_));
 AOI21_X1 _40104_ (.A(_13708_),
    .B1(_13850_),
    .B2(_13851_),
    .ZN(_13852_));
 OR2_X4 _40105_ (.A1(_13849_),
    .A2(_13852_),
    .ZN(_13853_));
 NAND2_X2 _40106_ (.A1(_13797_),
    .A2(_12225_),
    .ZN(_13854_));
 OAI21_X1 _40107_ (.A(_12222_),
    .B1(_13814_),
    .B2(_13815_),
    .ZN(_13855_));
 AOI21_X1 _40108_ (.A(_13789_),
    .B1(_13854_),
    .B2(_13855_),
    .ZN(_13856_));
 NAND2_X2 _40109_ (.A1(_13797_),
    .A2(_12232_),
    .ZN(_13857_));
 OAI21_X1 _40110_ (.A(_12229_),
    .B1(_13814_),
    .B2(_13815_),
    .ZN(_13858_));
 AOI21_X1 _40111_ (.A(_13808_),
    .B1(_13857_),
    .B2(_13858_),
    .ZN(_13859_));
 OR2_X4 _40112_ (.A1(_13856_),
    .A2(_13859_),
    .ZN(_13860_));
 MUX2_X2 _40113_ (.A(_13853_),
    .B(_13860_),
    .S(_13704_),
    .Z(\icache.data_mem_data_li [92]));
 NAND2_X2 _40114_ (.A1(_13797_),
    .A2(_12242_),
    .ZN(_13861_));
 OAI21_X1 _40115_ (.A(_12239_),
    .B1(_13814_),
    .B2(_13815_),
    .ZN(_13862_));
 AOI21_X1 _40116_ (.A(_13844_),
    .B1(_13861_),
    .B2(_13862_),
    .ZN(_13863_));
 BUF_X8 _40117_ (.A(_11709_),
    .Z(_13864_));
 NAND2_X2 _40118_ (.A1(_13829_),
    .A2(_12250_),
    .ZN(_13865_));
 OAI21_X2 _40119_ (.A(_12247_),
    .B1(_13846_),
    .B2(_13847_),
    .ZN(_13866_));
 AOI21_X2 _40120_ (.A(_13864_),
    .B1(_13865_),
    .B2(_13866_),
    .ZN(_13867_));
 OR2_X4 _40121_ (.A1(_13863_),
    .A2(_13867_),
    .ZN(_13868_));
 NAND2_X2 _40122_ (.A1(_13829_),
    .A2(_12258_),
    .ZN(_13869_));
 OAI21_X2 _40123_ (.A(_12255_),
    .B1(_13846_),
    .B2(_13847_),
    .ZN(_13870_));
 AOI21_X2 _40124_ (.A(_13789_),
    .B1(_13869_),
    .B2(_13870_),
    .ZN(_13871_));
 NAND2_X2 _40125_ (.A1(_13797_),
    .A2(_12266_),
    .ZN(_13872_));
 OAI21_X1 _40126_ (.A(_12263_),
    .B1(_13814_),
    .B2(_13815_),
    .ZN(_13873_));
 AOI21_X1 _40127_ (.A(_13808_),
    .B1(_13872_),
    .B2(_13873_),
    .ZN(_13874_));
 OR2_X4 _40128_ (.A1(_13871_),
    .A2(_13874_),
    .ZN(_13875_));
 MUX2_X2 _40129_ (.A(_13868_),
    .B(_13875_),
    .S(_13704_),
    .Z(\icache.data_mem_data_li [93]));
 NAND2_X1 _40130_ (.A1(_13829_),
    .A2(_12274_),
    .ZN(_13876_));
 OAI21_X1 _40131_ (.A(_12271_),
    .B1(_13846_),
    .B2(_13847_),
    .ZN(_13877_));
 AOI21_X1 _40132_ (.A(_13844_),
    .B1(_13876_),
    .B2(_13877_),
    .ZN(_13878_));
 NAND2_X1 _40133_ (.A1(_13829_),
    .A2(_12281_),
    .ZN(_13879_));
 OAI21_X1 _40134_ (.A(_12278_),
    .B1(_13846_),
    .B2(_13847_),
    .ZN(_13880_));
 AOI21_X1 _40135_ (.A(_13864_),
    .B1(_13879_),
    .B2(_13880_),
    .ZN(_13881_));
 OR2_X4 _40136_ (.A1(_13878_),
    .A2(_13881_),
    .ZN(_13882_));
 BUF_X4 _40137_ (.A(_08490_),
    .Z(_13883_));
 NAND2_X1 _40138_ (.A1(_13883_),
    .A2(_12289_),
    .ZN(_13884_));
 OAI21_X1 _40139_ (.A(_12286_),
    .B1(_13814_),
    .B2(_13815_),
    .ZN(_13885_));
 AOI21_X1 _40140_ (.A(_13789_),
    .B1(_13884_),
    .B2(_13885_),
    .ZN(_13886_));
 NAND2_X1 _40141_ (.A1(_13883_),
    .A2(_12300_),
    .ZN(_13887_));
 OAI21_X2 _40142_ (.A(_12295_),
    .B1(_13814_),
    .B2(_13815_),
    .ZN(_13888_));
 AOI21_X2 _40143_ (.A(_13808_),
    .B1(_13887_),
    .B2(_13888_),
    .ZN(_13889_));
 OR2_X4 _40144_ (.A1(_13886_),
    .A2(_13889_),
    .ZN(_13890_));
 MUX2_X2 _40145_ (.A(_13882_),
    .B(_13890_),
    .S(_13704_),
    .Z(\icache.data_mem_data_li [94]));
 NAND2_X1 _40146_ (.A1(_13829_),
    .A2(_12311_),
    .ZN(_13891_));
 OAI21_X1 _40147_ (.A(_12307_),
    .B1(_13846_),
    .B2(_13847_),
    .ZN(_13892_));
 AOI21_X1 _40148_ (.A(_13844_),
    .B1(_13891_),
    .B2(_13892_),
    .ZN(_13893_));
 NAND2_X2 _40149_ (.A1(_13829_),
    .A2(_12318_),
    .ZN(_13894_));
 OAI21_X2 _40150_ (.A(_12315_),
    .B1(_13846_),
    .B2(_13847_),
    .ZN(_13895_));
 AOI21_X2 _40151_ (.A(_13864_),
    .B1(_13894_),
    .B2(_13895_),
    .ZN(_13896_));
 OR2_X4 _40152_ (.A1(_13893_),
    .A2(_13896_),
    .ZN(_13897_));
 NAND2_X1 _40153_ (.A1(_13883_),
    .A2(_12326_),
    .ZN(_13898_));
 BUF_X4 _40154_ (.A(_11269_),
    .Z(_13899_));
 BUF_X4 _40155_ (.A(_11271_),
    .Z(_13900_));
 OAI21_X1 _40156_ (.A(_12323_),
    .B1(_13899_),
    .B2(_13900_),
    .ZN(_13901_));
 AOI21_X1 _40157_ (.A(_13789_),
    .B1(_13898_),
    .B2(_13901_),
    .ZN(_13902_));
 NAND2_X1 _40158_ (.A1(_13883_),
    .A2(_12333_),
    .ZN(_13903_));
 OAI21_X1 _40159_ (.A(_12330_),
    .B1(_13899_),
    .B2(_13900_),
    .ZN(_13904_));
 AOI21_X1 _40160_ (.A(_13808_),
    .B1(_13903_),
    .B2(_13904_),
    .ZN(_13905_));
 OR2_X4 _40161_ (.A1(_13902_),
    .A2(_13905_),
    .ZN(_13906_));
 MUX2_X2 _40162_ (.A(_13897_),
    .B(_13906_),
    .S(_13482_),
    .Z(\icache.data_mem_data_li [95]));
 BUF_X4 _40163_ (.A(_12973_),
    .Z(_13907_));
 NAND2_X1 _40164_ (.A1(_13907_),
    .A2(_12362_),
    .ZN(_13908_));
 OAI21_X1 _40165_ (.A(_12359_),
    .B1(_13846_),
    .B2(_13847_),
    .ZN(_13909_));
 AOI21_X1 _40166_ (.A(_13844_),
    .B1(_13908_),
    .B2(_13909_),
    .ZN(_13910_));
 NAND2_X1 _40167_ (.A1(_13907_),
    .A2(_12369_),
    .ZN(_13911_));
 OAI21_X1 _40168_ (.A(_12366_),
    .B1(_13846_),
    .B2(_13847_),
    .ZN(_13912_));
 AOI21_X1 _40169_ (.A(_13864_),
    .B1(_13911_),
    .B2(_13912_),
    .ZN(_13913_));
 OR2_X4 _40170_ (.A1(_13910_),
    .A2(_13913_),
    .ZN(_13914_));
 NAND2_X1 _40171_ (.A1(_13883_),
    .A2(_12344_),
    .ZN(_13915_));
 OAI21_X1 _40172_ (.A(_12340_),
    .B1(_13899_),
    .B2(_13900_),
    .ZN(_13916_));
 AOI21_X1 _40173_ (.A(_13789_),
    .B1(_13915_),
    .B2(_13916_),
    .ZN(_13917_));
 NAND2_X1 _40174_ (.A1(_13883_),
    .A2(_12352_),
    .ZN(_13918_));
 OAI21_X1 _40175_ (.A(_12348_),
    .B1(_13899_),
    .B2(_13900_),
    .ZN(_13919_));
 AOI21_X1 _40176_ (.A(_13808_),
    .B1(_13918_),
    .B2(_13919_),
    .ZN(_13920_));
 OR2_X4 _40177_ (.A1(_13917_),
    .A2(_13920_),
    .ZN(_13921_));
 BUF_X8 _40178_ (.A(_12640_),
    .Z(_13922_));
 MUX2_X2 _40179_ (.A(_13914_),
    .B(_13921_),
    .S(_13922_),
    .Z(\icache.data_mem_data_li [96]));
 NAND2_X1 _40180_ (.A1(_13883_),
    .A2(_12378_),
    .ZN(_13923_));
 OAI21_X1 _40181_ (.A(_12375_),
    .B1(_13899_),
    .B2(_13900_),
    .ZN(_13924_));
 AOI21_X1 _40182_ (.A(_13844_),
    .B1(_13923_),
    .B2(_13924_),
    .ZN(_13925_));
 NAND2_X1 _40183_ (.A1(_13907_),
    .A2(_12386_),
    .ZN(_13926_));
 BUF_X4 _40184_ (.A(_13342_),
    .Z(_13927_));
 BUF_X4 _40185_ (.A(_13344_),
    .Z(_13928_));
 OAI21_X2 _40186_ (.A(_12383_),
    .B1(_13927_),
    .B2(_13928_),
    .ZN(_13929_));
 AOI21_X2 _40187_ (.A(_13864_),
    .B1(_13926_),
    .B2(_13929_),
    .ZN(_13930_));
 OR2_X4 _40188_ (.A1(_13925_),
    .A2(_13930_),
    .ZN(_13931_));
 NAND2_X1 _40189_ (.A1(_13907_),
    .A2(_12394_),
    .ZN(_13932_));
 OAI21_X1 _40190_ (.A(_12391_),
    .B1(_13927_),
    .B2(_13928_),
    .ZN(_13933_));
 AOI21_X1 _40191_ (.A(_13789_),
    .B1(_13932_),
    .B2(_13933_),
    .ZN(_13934_));
 NAND2_X1 _40192_ (.A1(_13883_),
    .A2(_12401_),
    .ZN(_13935_));
 OAI21_X1 _40193_ (.A(_12398_),
    .B1(_13899_),
    .B2(_13900_),
    .ZN(_13936_));
 AOI21_X1 _40194_ (.A(_13808_),
    .B1(_13935_),
    .B2(_13936_),
    .ZN(_13937_));
 OR2_X4 _40195_ (.A1(_13934_),
    .A2(_13937_),
    .ZN(_13938_));
 MUX2_X2 _40196_ (.A(_13931_),
    .B(_13938_),
    .S(_13922_),
    .Z(\icache.data_mem_data_li [97]));
 NAND2_X1 _40197_ (.A1(_13907_),
    .A2(_12410_),
    .ZN(_13939_));
 OAI21_X1 _40198_ (.A(_12407_),
    .B1(_13927_),
    .B2(_13928_),
    .ZN(_13940_));
 AOI21_X1 _40199_ (.A(_13844_),
    .B1(_13939_),
    .B2(_13940_),
    .ZN(_13941_));
 NAND2_X1 _40200_ (.A1(_13907_),
    .A2(_12417_),
    .ZN(_13942_));
 OAI21_X1 _40201_ (.A(_12414_),
    .B1(_13927_),
    .B2(_13928_),
    .ZN(_13943_));
 AOI21_X1 _40202_ (.A(_13864_),
    .B1(_13942_),
    .B2(_13943_),
    .ZN(_13944_));
 OR2_X4 _40203_ (.A1(_13941_),
    .A2(_13944_),
    .ZN(_13945_));
 BUF_X8 _40204_ (.A(_13472_),
    .Z(_13946_));
 NAND2_X1 _40205_ (.A1(_13883_),
    .A2(_12428_),
    .ZN(_13947_));
 OAI21_X1 _40206_ (.A(_12425_),
    .B1(_13899_),
    .B2(_13900_),
    .ZN(_13948_));
 AOI21_X1 _40207_ (.A(_13946_),
    .B1(_13947_),
    .B2(_13948_),
    .ZN(_13949_));
 NAND2_X1 _40208_ (.A1(_13883_),
    .A2(_12435_),
    .ZN(_13950_));
 OAI21_X2 _40209_ (.A(_12432_),
    .B1(_13899_),
    .B2(_13900_),
    .ZN(_13951_));
 AOI21_X2 _40210_ (.A(_13808_),
    .B1(_13950_),
    .B2(_13951_),
    .ZN(_13952_));
 OR2_X4 _40211_ (.A1(_13949_),
    .A2(_13952_),
    .ZN(_13953_));
 MUX2_X2 _40212_ (.A(_13945_),
    .B(_13953_),
    .S(_13922_),
    .Z(\icache.data_mem_data_li [98]));
 NAND2_X1 _40213_ (.A1(_13907_),
    .A2(_12444_),
    .ZN(_13954_));
 OAI21_X1 _40214_ (.A(_12441_),
    .B1(_13927_),
    .B2(_13928_),
    .ZN(_13955_));
 AOI21_X1 _40215_ (.A(_13844_),
    .B1(_13954_),
    .B2(_13955_),
    .ZN(_13956_));
 NAND2_X1 _40216_ (.A1(_13907_),
    .A2(_12451_),
    .ZN(_13957_));
 OAI21_X1 _40217_ (.A(_12448_),
    .B1(_13927_),
    .B2(_13928_),
    .ZN(_13958_));
 AOI21_X1 _40218_ (.A(_13864_),
    .B1(_13957_),
    .B2(_13958_),
    .ZN(_13959_));
 OR2_X4 _40219_ (.A1(_13956_),
    .A2(_13959_),
    .ZN(_13960_));
 BUF_X4 _40220_ (.A(_08490_),
    .Z(_13961_));
 NAND2_X1 _40221_ (.A1(_13961_),
    .A2(_12459_),
    .ZN(_13962_));
 OAI21_X1 _40222_ (.A(_12456_),
    .B1(_13899_),
    .B2(_13900_),
    .ZN(_13963_));
 AOI21_X1 _40223_ (.A(_13946_),
    .B1(_13962_),
    .B2(_13963_),
    .ZN(_13964_));
 BUF_X8 _40224_ (.A(_13494_),
    .Z(_13965_));
 NAND2_X1 _40225_ (.A1(_13961_),
    .A2(_12469_),
    .ZN(_13966_));
 OAI21_X1 _40226_ (.A(_12466_),
    .B1(_13899_),
    .B2(_13900_),
    .ZN(_13967_));
 AOI21_X1 _40227_ (.A(_13965_),
    .B1(_13966_),
    .B2(_13967_),
    .ZN(_13968_));
 OR2_X4 _40228_ (.A1(_13964_),
    .A2(_13968_),
    .ZN(_13969_));
 MUX2_X2 _40229_ (.A(_13960_),
    .B(_13969_),
    .S(_13922_),
    .Z(\icache.data_mem_data_li [99]));
 NAND2_X1 _40230_ (.A1(_13961_),
    .A2(_12495_),
    .ZN(_13970_));
 BUF_X4 _40231_ (.A(_11269_),
    .Z(_13971_));
 BUF_X4 _40232_ (.A(_11271_),
    .Z(_13972_));
 OAI21_X1 _40233_ (.A(_12492_),
    .B1(_13971_),
    .B2(_13972_),
    .ZN(_13973_));
 AOI21_X1 _40234_ (.A(_13844_),
    .B1(_13970_),
    .B2(_13973_),
    .ZN(_13974_));
 NAND2_X1 _40235_ (.A1(_13907_),
    .A2(_12502_),
    .ZN(_13975_));
 OAI21_X1 _40236_ (.A(_12499_),
    .B1(_13927_),
    .B2(_13928_),
    .ZN(_13976_));
 AOI21_X1 _40237_ (.A(_13864_),
    .B1(_13975_),
    .B2(_13976_),
    .ZN(_13977_));
 OR2_X4 _40238_ (.A1(_13974_),
    .A2(_13977_),
    .ZN(_13978_));
 NAND2_X1 _40239_ (.A1(_13907_),
    .A2(_12479_),
    .ZN(_13979_));
 OAI21_X1 _40240_ (.A(_12475_),
    .B1(_13927_),
    .B2(_13928_),
    .ZN(_13980_));
 AOI21_X2 _40241_ (.A(_13946_),
    .B1(_13979_),
    .B2(_13980_),
    .ZN(_13981_));
 NAND2_X1 _40242_ (.A1(_13961_),
    .A2(_12487_),
    .ZN(_13982_));
 OAI21_X1 _40243_ (.A(_12484_),
    .B1(_13971_),
    .B2(_13972_),
    .ZN(_13983_));
 AOI21_X1 _40244_ (.A(_13965_),
    .B1(_13982_),
    .B2(_13983_),
    .ZN(_13984_));
 OR2_X4 _40245_ (.A1(_13981_),
    .A2(_13984_),
    .ZN(_13985_));
 MUX2_X2 _40246_ (.A(_13978_),
    .B(_13985_),
    .S(_13482_),
    .Z(\icache.data_mem_data_li [100]));
 NAND2_X1 _40247_ (.A1(_13961_),
    .A2(_12510_),
    .ZN(_13986_));
 OAI21_X1 _40248_ (.A(_12507_),
    .B1(_13971_),
    .B2(_13972_),
    .ZN(_13987_));
 AOI21_X1 _40249_ (.A(_13844_),
    .B1(_13986_),
    .B2(_13987_),
    .ZN(_13988_));
 BUF_X4 _40250_ (.A(_08489_),
    .Z(_13989_));
 NAND2_X1 _40251_ (.A1(_13989_),
    .A2(_12518_),
    .ZN(_13990_));
 OAI21_X1 _40252_ (.A(_12514_),
    .B1(_13927_),
    .B2(_13928_),
    .ZN(_13991_));
 AOI21_X1 _40253_ (.A(_13864_),
    .B1(_13990_),
    .B2(_13991_),
    .ZN(_13992_));
 OR2_X4 _40254_ (.A1(_13988_),
    .A2(_13992_),
    .ZN(_13993_));
 NAND2_X1 _40255_ (.A1(_13989_),
    .A2(_12528_),
    .ZN(_13994_));
 OAI21_X1 _40256_ (.A(_12525_),
    .B1(_13927_),
    .B2(_13928_),
    .ZN(_13995_));
 AOI21_X1 _40257_ (.A(_13946_),
    .B1(_13994_),
    .B2(_13995_),
    .ZN(_13996_));
 NAND2_X1 _40258_ (.A1(_13961_),
    .A2(_12535_),
    .ZN(_13997_));
 OAI21_X1 _40259_ (.A(_12532_),
    .B1(_13971_),
    .B2(_13972_),
    .ZN(_13998_));
 AOI21_X1 _40260_ (.A(_13965_),
    .B1(_13997_),
    .B2(_13998_),
    .ZN(_13999_));
 OR2_X4 _40261_ (.A1(_13996_),
    .A2(_13999_),
    .ZN(_14000_));
 MUX2_X2 _40262_ (.A(_13993_),
    .B(_14000_),
    .S(_13922_),
    .Z(\icache.data_mem_data_li [101]));
 BUF_X8 _40263_ (.A(_11665_),
    .Z(_14001_));
 NAND2_X1 _40264_ (.A1(_13961_),
    .A2(_12544_),
    .ZN(_14002_));
 OAI21_X1 _40265_ (.A(_12541_),
    .B1(_13971_),
    .B2(_13972_),
    .ZN(_14003_));
 AOI21_X1 _40266_ (.A(_14001_),
    .B1(_14002_),
    .B2(_14003_),
    .ZN(_14004_));
 NAND2_X1 _40267_ (.A1(_13989_),
    .A2(_12551_),
    .ZN(_14005_));
 BUF_X4 _40268_ (.A(_13342_),
    .Z(_14006_));
 BUF_X4 _40269_ (.A(_13344_),
    .Z(_14007_));
 OAI21_X2 _40270_ (.A(_12548_),
    .B1(_14006_),
    .B2(_14007_),
    .ZN(_14008_));
 AOI21_X1 _40271_ (.A(_13864_),
    .B1(_14005_),
    .B2(_14008_),
    .ZN(_14009_));
 OR2_X4 _40272_ (.A1(_14004_),
    .A2(_14009_),
    .ZN(_14010_));
 NAND2_X1 _40273_ (.A1(_13989_),
    .A2(_12560_),
    .ZN(_14011_));
 OAI21_X1 _40274_ (.A(_12557_),
    .B1(_14006_),
    .B2(_14007_),
    .ZN(_14012_));
 AOI21_X1 _40275_ (.A(_13946_),
    .B1(_14011_),
    .B2(_14012_),
    .ZN(_14013_));
 NAND2_X1 _40276_ (.A1(_13961_),
    .A2(_12567_),
    .ZN(_14014_));
 OAI21_X1 _40277_ (.A(_12564_),
    .B1(_13971_),
    .B2(_13972_),
    .ZN(_14015_));
 AOI21_X1 _40278_ (.A(_13965_),
    .B1(_14014_),
    .B2(_14015_),
    .ZN(_14016_));
 OR2_X4 _40279_ (.A1(_14013_),
    .A2(_14016_),
    .ZN(_14017_));
 MUX2_X2 _40280_ (.A(_14010_),
    .B(_14017_),
    .S(_13922_),
    .Z(\icache.data_mem_data_li [102]));
 NAND2_X1 _40281_ (.A1(_13989_),
    .A2(_12593_),
    .ZN(_14018_));
 OAI21_X1 _40282_ (.A(_12590_),
    .B1(_14006_),
    .B2(_14007_),
    .ZN(_14019_));
 AOI21_X1 _40283_ (.A(_14001_),
    .B1(_14018_),
    .B2(_14019_),
    .ZN(_14020_));
 BUF_X8 _40284_ (.A(_11709_),
    .Z(_14021_));
 NAND2_X1 _40285_ (.A1(_13989_),
    .A2(_12601_),
    .ZN(_14022_));
 OAI21_X1 _40286_ (.A(_12598_),
    .B1(_14006_),
    .B2(_14007_),
    .ZN(_14023_));
 AOI21_X1 _40287_ (.A(_14021_),
    .B1(_14022_),
    .B2(_14023_),
    .ZN(_14024_));
 OR2_X4 _40288_ (.A1(_14020_),
    .A2(_14024_),
    .ZN(_14025_));
 NAND2_X1 _40289_ (.A1(_13961_),
    .A2(_12577_),
    .ZN(_14026_));
 OAI21_X1 _40290_ (.A(_12573_),
    .B1(_13971_),
    .B2(_13972_),
    .ZN(_14027_));
 AOI21_X1 _40291_ (.A(_13946_),
    .B1(_14026_),
    .B2(_14027_),
    .ZN(_14028_));
 NAND2_X1 _40292_ (.A1(_13961_),
    .A2(_12585_),
    .ZN(_14029_));
 OAI21_X1 _40293_ (.A(_12581_),
    .B1(_13971_),
    .B2(_13972_),
    .ZN(_14030_));
 AOI21_X1 _40294_ (.A(_13965_),
    .B1(_14029_),
    .B2(_14030_),
    .ZN(_14031_));
 OR2_X4 _40295_ (.A1(_14028_),
    .A2(_14031_),
    .ZN(_14032_));
 MUX2_X2 _40296_ (.A(_14025_),
    .B(_14032_),
    .S(_13922_),
    .Z(\icache.data_mem_data_li [103]));
 NAND2_X1 _40297_ (.A1(_13989_),
    .A2(_12629_),
    .ZN(_14033_));
 OAI21_X1 _40298_ (.A(_12626_),
    .B1(_14006_),
    .B2(_14007_),
    .ZN(_14034_));
 AOI21_X1 _40299_ (.A(_14001_),
    .B1(_14033_),
    .B2(_14034_),
    .ZN(_14035_));
 NAND2_X1 _40300_ (.A1(_13989_),
    .A2(_12636_),
    .ZN(_14036_));
 OAI21_X1 _40301_ (.A(_12633_),
    .B1(_14006_),
    .B2(_14007_),
    .ZN(_14037_));
 AOI21_X1 _40302_ (.A(_14021_),
    .B1(_14036_),
    .B2(_14037_),
    .ZN(_14038_));
 OR2_X4 _40303_ (.A1(_14035_),
    .A2(_14038_),
    .ZN(_14039_));
 BUF_X4 _40304_ (.A(_08490_),
    .Z(_14040_));
 NAND2_X1 _40305_ (.A1(_14040_),
    .A2(_12609_),
    .ZN(_14041_));
 OAI21_X1 _40306_ (.A(_12606_),
    .B1(_13971_),
    .B2(_13972_),
    .ZN(_14042_));
 AOI21_X1 _40307_ (.A(_13946_),
    .B1(_14041_),
    .B2(_14042_),
    .ZN(_14043_));
 NAND2_X1 _40308_ (.A1(_14040_),
    .A2(_12621_),
    .ZN(_14044_));
 OAI21_X1 _40309_ (.A(_12617_),
    .B1(_13971_),
    .B2(_13972_),
    .ZN(_14045_));
 AOI21_X1 _40310_ (.A(_13965_),
    .B1(_14044_),
    .B2(_14045_),
    .ZN(_14046_));
 OR2_X4 _40311_ (.A1(_14043_),
    .A2(_14046_),
    .ZN(_14047_));
 BUF_X32 _40312_ (.A(_13481_),
    .Z(_14048_));
 MUX2_X2 _40313_ (.A(_14039_),
    .B(_14047_),
    .S(_14048_),
    .Z(\icache.data_mem_data_li [104]));
 NAND2_X1 _40314_ (.A1(_13989_),
    .A2(_12664_),
    .ZN(_14049_));
 OAI21_X1 _40315_ (.A(_12661_),
    .B1(_14006_),
    .B2(_14007_),
    .ZN(_14050_));
 AOI21_X1 _40316_ (.A(_14001_),
    .B1(_14049_),
    .B2(_14050_),
    .ZN(_14051_));
 NAND2_X1 _40317_ (.A1(_13989_),
    .A2(_12671_),
    .ZN(_14052_));
 OAI21_X1 _40318_ (.A(_12668_),
    .B1(_14006_),
    .B2(_14007_),
    .ZN(_14053_));
 AOI21_X1 _40319_ (.A(_14021_),
    .B1(_14052_),
    .B2(_14053_),
    .ZN(_14054_));
 OR2_X4 _40320_ (.A1(_14051_),
    .A2(_14054_),
    .ZN(_14055_));
 NAND2_X1 _40321_ (.A1(_14040_),
    .A2(_12648_),
    .ZN(_14056_));
 BUF_X4 _40322_ (.A(_11269_),
    .Z(_14057_));
 BUF_X4 _40323_ (.A(_11271_),
    .Z(_14058_));
 OAI21_X1 _40324_ (.A(_12644_),
    .B1(_14057_),
    .B2(_14058_),
    .ZN(_14059_));
 AOI21_X1 _40325_ (.A(_13946_),
    .B1(_14056_),
    .B2(_14059_),
    .ZN(_14060_));
 NAND2_X1 _40326_ (.A1(_14040_),
    .A2(_12656_),
    .ZN(_14061_));
 OAI21_X1 _40327_ (.A(_12653_),
    .B1(_14057_),
    .B2(_14058_),
    .ZN(_14062_));
 AOI21_X1 _40328_ (.A(_13965_),
    .B1(_14061_),
    .B2(_14062_),
    .ZN(_14063_));
 OR2_X4 _40329_ (.A1(_14060_),
    .A2(_14063_),
    .ZN(_14064_));
 MUX2_X2 _40330_ (.A(_14055_),
    .B(_14064_),
    .S(_13922_),
    .Z(\icache.data_mem_data_li [105]));
 BUF_X4 _40331_ (.A(_08489_),
    .Z(_14065_));
 NAND2_X1 _40332_ (.A1(_14065_),
    .A2(_12699_),
    .ZN(_14066_));
 OAI21_X1 _40333_ (.A(_12696_),
    .B1(_14006_),
    .B2(_14007_),
    .ZN(_14067_));
 AOI21_X1 _40334_ (.A(_14001_),
    .B1(_14066_),
    .B2(_14067_),
    .ZN(_14068_));
 NAND2_X1 _40335_ (.A1(_14065_),
    .A2(_12706_),
    .ZN(_14069_));
 OAI21_X1 _40336_ (.A(_12703_),
    .B1(_14006_),
    .B2(_14007_),
    .ZN(_14070_));
 AOI21_X1 _40337_ (.A(_14021_),
    .B1(_14069_),
    .B2(_14070_),
    .ZN(_14071_));
 OR2_X4 _40338_ (.A1(_14068_),
    .A2(_14071_),
    .ZN(_14072_));
 NAND2_X1 _40339_ (.A1(_14040_),
    .A2(_12681_),
    .ZN(_14073_));
 OAI21_X1 _40340_ (.A(_12677_),
    .B1(_14057_),
    .B2(_14058_),
    .ZN(_14074_));
 AOI21_X1 _40341_ (.A(_13946_),
    .B1(_14073_),
    .B2(_14074_),
    .ZN(_14075_));
 NAND2_X1 _40342_ (.A1(_14040_),
    .A2(_12691_),
    .ZN(_14076_));
 OAI21_X1 _40343_ (.A(_12688_),
    .B1(_14057_),
    .B2(_14058_),
    .ZN(_14077_));
 AOI21_X1 _40344_ (.A(_13965_),
    .B1(_14076_),
    .B2(_14077_),
    .ZN(_14078_));
 OR2_X4 _40345_ (.A1(_14075_),
    .A2(_14078_),
    .ZN(_14079_));
 MUX2_X2 _40346_ (.A(_14072_),
    .B(_14079_),
    .S(_13922_),
    .Z(\icache.data_mem_data_li [106]));
 NAND2_X1 _40347_ (.A1(_14065_),
    .A2(_12731_),
    .ZN(_14080_));
 BUF_X4 _40348_ (.A(_13342_),
    .Z(_14081_));
 BUF_X4 _40349_ (.A(_13344_),
    .Z(_14082_));
 OAI21_X1 _40350_ (.A(_12728_),
    .B1(_14081_),
    .B2(_14082_),
    .ZN(_14083_));
 AOI21_X1 _40351_ (.A(_14001_),
    .B1(_14080_),
    .B2(_14083_),
    .ZN(_14084_));
 NAND2_X1 _40352_ (.A1(_14065_),
    .A2(_12738_),
    .ZN(_14085_));
 OAI21_X1 _40353_ (.A(_12735_),
    .B1(_14081_),
    .B2(_14082_),
    .ZN(_14086_));
 AOI21_X1 _40354_ (.A(_14021_),
    .B1(_14085_),
    .B2(_14086_),
    .ZN(_14087_));
 OR2_X4 _40355_ (.A1(_14084_),
    .A2(_14087_),
    .ZN(_14088_));
 NAND2_X1 _40356_ (.A1(_14040_),
    .A2(_12714_),
    .ZN(_14089_));
 OAI21_X1 _40357_ (.A(_12711_),
    .B1(_14057_),
    .B2(_14058_),
    .ZN(_14090_));
 AOI21_X1 _40358_ (.A(_13946_),
    .B1(_14089_),
    .B2(_14090_),
    .ZN(_14091_));
 NAND2_X1 _40359_ (.A1(_14040_),
    .A2(_12723_),
    .ZN(_14092_));
 OAI21_X1 _40360_ (.A(_12719_),
    .B1(_14057_),
    .B2(_14058_),
    .ZN(_14093_));
 AOI21_X1 _40361_ (.A(_13965_),
    .B1(_14092_),
    .B2(_14093_),
    .ZN(_14094_));
 OR2_X4 _40362_ (.A1(_14091_),
    .A2(_14094_),
    .ZN(_14095_));
 MUX2_X2 _40363_ (.A(_14088_),
    .B(_14095_),
    .S(_13922_),
    .Z(\icache.data_mem_data_li [107]));
 NAND2_X1 _40364_ (.A1(_14040_),
    .A2(_12748_),
    .ZN(_14096_));
 OAI21_X1 _40365_ (.A(_12745_),
    .B1(_14057_),
    .B2(_14058_),
    .ZN(_14097_));
 AOI21_X1 _40366_ (.A(_14001_),
    .B1(_14096_),
    .B2(_14097_),
    .ZN(_14098_));
 NAND2_X1 _40367_ (.A1(_14065_),
    .A2(_12755_),
    .ZN(_14099_));
 OAI21_X1 _40368_ (.A(_12752_),
    .B1(_14081_),
    .B2(_14082_),
    .ZN(_14100_));
 AOI21_X1 _40369_ (.A(_14021_),
    .B1(_14099_),
    .B2(_14100_),
    .ZN(_14101_));
 OR2_X4 _40370_ (.A1(_14098_),
    .A2(_14101_),
    .ZN(_14102_));
 BUF_X8 _40371_ (.A(_13472_),
    .Z(_14103_));
 NAND2_X1 _40372_ (.A1(_14065_),
    .A2(_12763_),
    .ZN(_14104_));
 OAI21_X1 _40373_ (.A(_12760_),
    .B1(_14081_),
    .B2(_14082_),
    .ZN(_14105_));
 AOI21_X1 _40374_ (.A(_14103_),
    .B1(_14104_),
    .B2(_14105_),
    .ZN(_14106_));
 NAND2_X1 _40375_ (.A1(_14040_),
    .A2(_12770_),
    .ZN(_14107_));
 OAI21_X1 _40376_ (.A(_12767_),
    .B1(_14057_),
    .B2(_14058_),
    .ZN(_14108_));
 AOI21_X2 _40377_ (.A(_13965_),
    .B1(_14107_),
    .B2(_14108_),
    .ZN(_14109_));
 OR2_X4 _40378_ (.A1(_14106_),
    .A2(_14109_),
    .ZN(_14110_));
 BUF_X8 _40379_ (.A(_12640_),
    .Z(_14111_));
 MUX2_X2 _40380_ (.A(_14102_),
    .B(_14110_),
    .S(_14111_),
    .Z(\icache.data_mem_data_li [108]));
 BUF_X4 _40381_ (.A(_08490_),
    .Z(_14112_));
 NAND2_X1 _40382_ (.A1(_14112_),
    .A2(_12779_),
    .ZN(_14113_));
 OAI21_X1 _40383_ (.A(_12776_),
    .B1(_14057_),
    .B2(_14058_),
    .ZN(_14114_));
 AOI21_X1 _40384_ (.A(_14001_),
    .B1(_14113_),
    .B2(_14114_),
    .ZN(_14115_));
 NAND2_X1 _40385_ (.A1(_14065_),
    .A2(_12789_),
    .ZN(_14116_));
 OAI21_X1 _40386_ (.A(_12786_),
    .B1(_14081_),
    .B2(_14082_),
    .ZN(_14117_));
 AOI21_X1 _40387_ (.A(_14021_),
    .B1(_14116_),
    .B2(_14117_),
    .ZN(_14118_));
 OR2_X4 _40388_ (.A1(_14115_),
    .A2(_14118_),
    .ZN(_14119_));
 NAND2_X1 _40389_ (.A1(_14065_),
    .A2(_12797_),
    .ZN(_14120_));
 OAI21_X1 _40390_ (.A(_12794_),
    .B1(_14081_),
    .B2(_14082_),
    .ZN(_14121_));
 AOI21_X1 _40391_ (.A(_14103_),
    .B1(_14120_),
    .B2(_14121_),
    .ZN(_14122_));
 BUF_X8 _40392_ (.A(_13494_),
    .Z(_14123_));
 NAND2_X1 _40393_ (.A1(_14112_),
    .A2(_12804_),
    .ZN(_14124_));
 OAI21_X1 _40394_ (.A(_12801_),
    .B1(_14057_),
    .B2(_14058_),
    .ZN(_14125_));
 AOI21_X1 _40395_ (.A(_14123_),
    .B1(_14124_),
    .B2(_14125_),
    .ZN(_14126_));
 OR2_X4 _40396_ (.A1(_14122_),
    .A2(_14126_),
    .ZN(_14127_));
 MUX2_X2 _40397_ (.A(_14119_),
    .B(_14127_),
    .S(_14111_),
    .Z(\icache.data_mem_data_li [109]));
 NAND2_X1 _40398_ (.A1(_14112_),
    .A2(_12829_),
    .ZN(_14128_));
 BUF_X8 _40399_ (.A(_11269_),
    .Z(_14129_));
 BUF_X8 _40400_ (.A(_11271_),
    .Z(_14130_));
 OAI21_X1 _40401_ (.A(_12826_),
    .B1(_14129_),
    .B2(_14130_),
    .ZN(_14131_));
 AOI21_X1 _40402_ (.A(_14001_),
    .B1(_14128_),
    .B2(_14131_),
    .ZN(_14132_));
 NAND2_X1 _40403_ (.A1(_14065_),
    .A2(_12836_),
    .ZN(_14133_));
 OAI21_X1 _40404_ (.A(_12833_),
    .B1(_14081_),
    .B2(_14082_),
    .ZN(_14134_));
 AOI21_X1 _40405_ (.A(_14021_),
    .B1(_14133_),
    .B2(_14134_),
    .ZN(_14135_));
 OR2_X4 _40406_ (.A1(_14132_),
    .A2(_14135_),
    .ZN(_14136_));
 NAND2_X1 _40407_ (.A1(_14065_),
    .A2(_12814_),
    .ZN(_14137_));
 OAI21_X1 _40408_ (.A(_12811_),
    .B1(_14081_),
    .B2(_14082_),
    .ZN(_14138_));
 AOI21_X2 _40409_ (.A(_14103_),
    .B1(_14137_),
    .B2(_14138_),
    .ZN(_14139_));
 NAND2_X1 _40410_ (.A1(_14112_),
    .A2(_12821_),
    .ZN(_14140_));
 OAI21_X1 _40411_ (.A(_12818_),
    .B1(_14129_),
    .B2(_14130_),
    .ZN(_14141_));
 AOI21_X1 _40412_ (.A(_14123_),
    .B1(_14140_),
    .B2(_14141_),
    .ZN(_14142_));
 OR2_X4 _40413_ (.A1(_14139_),
    .A2(_14142_),
    .ZN(_14143_));
 MUX2_X2 _40414_ (.A(_14136_),
    .B(_14143_),
    .S(_14048_),
    .Z(\icache.data_mem_data_li [110]));
 BUF_X4 _40415_ (.A(_08489_),
    .Z(_14144_));
 NAND2_X1 _40416_ (.A1(_14144_),
    .A2(_12862_),
    .ZN(_14145_));
 OAI21_X1 _40417_ (.A(_12859_),
    .B1(_14081_),
    .B2(_14082_),
    .ZN(_14146_));
 AOI21_X1 _40418_ (.A(_14001_),
    .B1(_14145_),
    .B2(_14146_),
    .ZN(_14147_));
 NAND2_X1 _40419_ (.A1(_14144_),
    .A2(_12869_),
    .ZN(_14148_));
 OAI21_X1 _40420_ (.A(_12866_),
    .B1(_14081_),
    .B2(_14082_),
    .ZN(_14149_));
 AOI21_X1 _40421_ (.A(_14021_),
    .B1(_14148_),
    .B2(_14149_),
    .ZN(_14150_));
 OR2_X4 _40422_ (.A1(_14147_),
    .A2(_14150_),
    .ZN(_14151_));
 NAND2_X1 _40423_ (.A1(_14112_),
    .A2(_12845_),
    .ZN(_14152_));
 OAI21_X1 _40424_ (.A(_12842_),
    .B1(_14129_),
    .B2(_14130_),
    .ZN(_14153_));
 AOI21_X1 _40425_ (.A(_14103_),
    .B1(_14152_),
    .B2(_14153_),
    .ZN(_14154_));
 NAND2_X1 _40426_ (.A1(_14112_),
    .A2(_12852_),
    .ZN(_14155_));
 OAI21_X1 _40427_ (.A(_12849_),
    .B1(_14129_),
    .B2(_14130_),
    .ZN(_14156_));
 AOI21_X1 _40428_ (.A(_14123_),
    .B1(_14155_),
    .B2(_14156_),
    .ZN(_14157_));
 OR2_X4 _40429_ (.A1(_14154_),
    .A2(_14157_),
    .ZN(_14158_));
 MUX2_X2 _40430_ (.A(_14151_),
    .B(_14158_),
    .S(_14048_),
    .Z(\icache.data_mem_data_li [111]));
 BUF_X32 _40431_ (.A(_08447_),
    .Z(_14159_));
 BUF_X8 _40432_ (.A(_14159_),
    .Z(_14160_));
 NAND2_X1 _40433_ (.A1(_14112_),
    .A2(_12878_),
    .ZN(_14161_));
 OAI21_X2 _40434_ (.A(_12874_),
    .B1(_14129_),
    .B2(_14130_),
    .ZN(_14162_));
 AOI21_X2 _40435_ (.A(_14160_),
    .B1(_14161_),
    .B2(_14162_),
    .ZN(_14163_));
 NAND2_X1 _40436_ (.A1(_14144_),
    .A2(_12886_),
    .ZN(_14164_));
 BUF_X4 _40437_ (.A(_08483_),
    .Z(_14165_));
 BUF_X8 _40438_ (.A(_08487_),
    .Z(_14166_));
 OAI21_X2 _40439_ (.A(_12883_),
    .B1(_14165_),
    .B2(_14166_),
    .ZN(_14167_));
 AOI21_X1 _40440_ (.A(_14021_),
    .B1(_14164_),
    .B2(_14167_),
    .ZN(_14168_));
 OR2_X4 _40441_ (.A1(_14163_),
    .A2(_14168_),
    .ZN(_14169_));
 NAND2_X1 _40442_ (.A1(_14144_),
    .A2(_12895_),
    .ZN(_14170_));
 OAI21_X1 _40443_ (.A(_12892_),
    .B1(_14165_),
    .B2(_14166_),
    .ZN(_14171_));
 AOI21_X1 _40444_ (.A(_14103_),
    .B1(_14170_),
    .B2(_14171_),
    .ZN(_14172_));
 NAND2_X1 _40445_ (.A1(_14112_),
    .A2(_12902_),
    .ZN(_14173_));
 OAI21_X1 _40446_ (.A(_12899_),
    .B1(_14129_),
    .B2(_14130_),
    .ZN(_14174_));
 AOI21_X1 _40447_ (.A(_14123_),
    .B1(_14173_),
    .B2(_14174_),
    .ZN(_14175_));
 OR2_X4 _40448_ (.A1(_14172_),
    .A2(_14175_),
    .ZN(_14176_));
 MUX2_X2 _40449_ (.A(_14169_),
    .B(_14176_),
    .S(_14048_),
    .Z(\icache.data_mem_data_li [112]));
 NAND2_X1 _40450_ (.A1(_14112_),
    .A2(_12912_),
    .ZN(_14177_));
 OAI21_X1 _40451_ (.A(_12908_),
    .B1(_14129_),
    .B2(_14130_),
    .ZN(_14178_));
 AOI21_X1 _40452_ (.A(_14160_),
    .B1(_14177_),
    .B2(_14178_),
    .ZN(_14179_));
 BUF_X32 _40453_ (.A(_08446_),
    .Z(_14180_));
 BUF_X8 _40454_ (.A(_14180_),
    .Z(_14181_));
 NAND2_X1 _40455_ (.A1(_14144_),
    .A2(_12920_),
    .ZN(_14182_));
 OAI21_X1 _40456_ (.A(_12917_),
    .B1(_14165_),
    .B2(_14166_),
    .ZN(_14183_));
 AOI21_X1 _40457_ (.A(_14181_),
    .B1(_14182_),
    .B2(_14183_),
    .ZN(_14184_));
 OR2_X4 _40458_ (.A1(_14179_),
    .A2(_14184_),
    .ZN(_14185_));
 NAND2_X1 _40459_ (.A1(_14144_),
    .A2(_12928_),
    .ZN(_14186_));
 OAI21_X1 _40460_ (.A(_12925_),
    .B1(_14165_),
    .B2(_14166_),
    .ZN(_14187_));
 AOI21_X1 _40461_ (.A(_14103_),
    .B1(_14186_),
    .B2(_14187_),
    .ZN(_14188_));
 NAND2_X1 _40462_ (.A1(_14112_),
    .A2(_12936_),
    .ZN(_14189_));
 OAI21_X2 _40463_ (.A(_12933_),
    .B1(_14129_),
    .B2(_14130_),
    .ZN(_14190_));
 AOI21_X2 _40464_ (.A(_14123_),
    .B1(_14189_),
    .B2(_14190_),
    .ZN(_14191_));
 OR2_X4 _40465_ (.A1(_14188_),
    .A2(_14191_),
    .ZN(_14192_));
 MUX2_X2 _40466_ (.A(_14185_),
    .B(_14192_),
    .S(_14111_),
    .Z(\icache.data_mem_data_li [113]));
 NAND2_X1 _40467_ (.A1(_14144_),
    .A2(_12944_),
    .ZN(_14193_));
 OAI21_X1 _40468_ (.A(_12941_),
    .B1(_14165_),
    .B2(_14166_),
    .ZN(_14194_));
 AOI21_X1 _40469_ (.A(_14160_),
    .B1(_14193_),
    .B2(_14194_),
    .ZN(_14195_));
 NAND2_X1 _40470_ (.A1(_14144_),
    .A2(_12952_),
    .ZN(_14196_));
 OAI21_X1 _40471_ (.A(_12948_),
    .B1(_14165_),
    .B2(_14166_),
    .ZN(_14197_));
 AOI21_X1 _40472_ (.A(_14181_),
    .B1(_14196_),
    .B2(_14197_),
    .ZN(_14198_));
 OR2_X4 _40473_ (.A1(_14195_),
    .A2(_14198_),
    .ZN(_14199_));
 BUF_X4 _40474_ (.A(_08490_),
    .Z(_14200_));
 NAND2_X1 _40475_ (.A1(_14200_),
    .A2(_12960_),
    .ZN(_14201_));
 OAI21_X2 _40476_ (.A(_12957_),
    .B1(_14129_),
    .B2(_14130_),
    .ZN(_14202_));
 AOI21_X1 _40477_ (.A(_14103_),
    .B1(_14201_),
    .B2(_14202_),
    .ZN(_14203_));
 NAND2_X1 _40478_ (.A1(_14200_),
    .A2(_12969_),
    .ZN(_14204_));
 OAI21_X2 _40479_ (.A(_12966_),
    .B1(_14129_),
    .B2(_14130_),
    .ZN(_14205_));
 AOI21_X2 _40480_ (.A(_14123_),
    .B1(_14204_),
    .B2(_14205_),
    .ZN(_14206_));
 OR2_X4 _40481_ (.A1(_14203_),
    .A2(_14206_),
    .ZN(_14207_));
 MUX2_X2 _40482_ (.A(_14199_),
    .B(_14207_),
    .S(_14111_),
    .Z(\icache.data_mem_data_li [114]));
 NAND2_X1 _40483_ (.A1(_14144_),
    .A2(_12979_),
    .ZN(_14208_));
 OAI21_X1 _40484_ (.A(_12976_),
    .B1(_14165_),
    .B2(_14166_),
    .ZN(_14209_));
 AOI21_X1 _40485_ (.A(_14160_),
    .B1(_14208_),
    .B2(_14209_),
    .ZN(_14210_));
 NAND2_X1 _40486_ (.A1(_14144_),
    .A2(_12987_),
    .ZN(_14211_));
 OAI21_X1 _40487_ (.A(_12983_),
    .B1(_14165_),
    .B2(_14166_),
    .ZN(_14212_));
 AOI21_X1 _40488_ (.A(_14181_),
    .B1(_14211_),
    .B2(_14212_),
    .ZN(_14213_));
 OR2_X4 _40489_ (.A1(_14210_),
    .A2(_14213_),
    .ZN(_14214_));
 NAND2_X1 _40490_ (.A1(_14200_),
    .A2(_12996_),
    .ZN(_14215_));
 BUF_X4 _40491_ (.A(_11269_),
    .Z(_14216_));
 BUF_X4 _40492_ (.A(_11271_),
    .Z(_14217_));
 OAI21_X2 _40493_ (.A(_12992_),
    .B1(_14216_),
    .B2(_14217_),
    .ZN(_14218_));
 AOI21_X1 _40494_ (.A(_14103_),
    .B1(_14215_),
    .B2(_14218_),
    .ZN(_14219_));
 NAND2_X1 _40495_ (.A1(_14200_),
    .A2(_13003_),
    .ZN(_14220_));
 OAI21_X2 _40496_ (.A(_13000_),
    .B1(_14216_),
    .B2(_14217_),
    .ZN(_14221_));
 AOI21_X2 _40497_ (.A(_14123_),
    .B1(_14220_),
    .B2(_14221_),
    .ZN(_14222_));
 OR2_X4 _40498_ (.A1(_14219_),
    .A2(_14222_),
    .ZN(_14223_));
 MUX2_X2 _40499_ (.A(_14214_),
    .B(_14223_),
    .S(_14111_),
    .Z(\icache.data_mem_data_li [115]));
 NAND2_X1 _40500_ (.A1(_14200_),
    .A2(_13012_),
    .ZN(_14224_));
 OAI21_X2 _40501_ (.A(_13009_),
    .B1(_14216_),
    .B2(_14217_),
    .ZN(_14225_));
 AOI21_X2 _40502_ (.A(_14160_),
    .B1(_14224_),
    .B2(_14225_),
    .ZN(_14226_));
 BUF_X4 _40503_ (.A(_08489_),
    .Z(_14227_));
 NAND2_X1 _40504_ (.A1(_14227_),
    .A2(_13019_),
    .ZN(_14228_));
 OAI21_X2 _40505_ (.A(_13016_),
    .B1(_14165_),
    .B2(_14166_),
    .ZN(_14229_));
 AOI21_X1 _40506_ (.A(_14181_),
    .B1(_14228_),
    .B2(_14229_),
    .ZN(_14230_));
 OR2_X4 _40507_ (.A1(_14226_),
    .A2(_14230_),
    .ZN(_14231_));
 NAND2_X1 _40508_ (.A1(_14227_),
    .A2(_13029_),
    .ZN(_14232_));
 OAI21_X1 _40509_ (.A(_13026_),
    .B1(_14165_),
    .B2(_14166_),
    .ZN(_14233_));
 AOI21_X1 _40510_ (.A(_14103_),
    .B1(_14232_),
    .B2(_14233_),
    .ZN(_14234_));
 NAND2_X1 _40511_ (.A1(_14200_),
    .A2(_13036_),
    .ZN(_14235_));
 OAI21_X2 _40512_ (.A(_13033_),
    .B1(_14216_),
    .B2(_14217_),
    .ZN(_14236_));
 AOI21_X2 _40513_ (.A(_14123_),
    .B1(_14235_),
    .B2(_14236_),
    .ZN(_14237_));
 OR2_X4 _40514_ (.A1(_14234_),
    .A2(_14237_),
    .ZN(_14238_));
 MUX2_X2 _40515_ (.A(_14231_),
    .B(_14238_),
    .S(_14048_),
    .Z(\icache.data_mem_data_li [116]));
 NAND2_X1 _40516_ (.A1(_14227_),
    .A2(_13045_),
    .ZN(_14239_));
 BUF_X4 _40517_ (.A(_08483_),
    .Z(_14240_));
 BUF_X4 _40518_ (.A(_08487_),
    .Z(_14241_));
 OAI21_X1 _40519_ (.A(_13041_),
    .B1(_14240_),
    .B2(_14241_),
    .ZN(_14242_));
 AOI21_X1 _40520_ (.A(_14160_),
    .B1(_14239_),
    .B2(_14242_),
    .ZN(_14243_));
 NAND2_X1 _40521_ (.A1(_14227_),
    .A2(_13053_),
    .ZN(_14244_));
 OAI21_X1 _40522_ (.A(_13050_),
    .B1(_14240_),
    .B2(_14241_),
    .ZN(_14245_));
 AOI21_X1 _40523_ (.A(_14181_),
    .B1(_14244_),
    .B2(_14245_),
    .ZN(_14246_));
 OR2_X4 _40524_ (.A1(_14243_),
    .A2(_14246_),
    .ZN(_14247_));
 NAND2_X1 _40525_ (.A1(_14200_),
    .A2(_13062_),
    .ZN(_14248_));
 OAI21_X1 _40526_ (.A(_13058_),
    .B1(_14216_),
    .B2(_14217_),
    .ZN(_14249_));
 AOI21_X1 _40527_ (.A(_14103_),
    .B1(_14248_),
    .B2(_14249_),
    .ZN(_14250_));
 NAND2_X1 _40528_ (.A1(_14200_),
    .A2(_13069_),
    .ZN(_14251_));
 OAI21_X1 _40529_ (.A(_13066_),
    .B1(_14216_),
    .B2(_14217_),
    .ZN(_14252_));
 AOI21_X1 _40530_ (.A(_14123_),
    .B1(_14251_),
    .B2(_14252_),
    .ZN(_14253_));
 OR2_X4 _40531_ (.A1(_14250_),
    .A2(_14253_),
    .ZN(_14254_));
 MUX2_X2 _40532_ (.A(_14247_),
    .B(_14254_),
    .S(_14111_),
    .Z(\icache.data_mem_data_li [117]));
 NAND2_X1 _40533_ (.A1(_14200_),
    .A2(_13095_),
    .ZN(_14255_));
 OAI21_X1 _40534_ (.A(_13092_),
    .B1(_14216_),
    .B2(_14217_),
    .ZN(_14256_));
 AOI21_X1 _40535_ (.A(_14160_),
    .B1(_14255_),
    .B2(_14256_),
    .ZN(_14257_));
 NAND2_X1 _40536_ (.A1(_14227_),
    .A2(_13102_),
    .ZN(_14258_));
 OAI21_X1 _40537_ (.A(_13099_),
    .B1(_14240_),
    .B2(_14241_),
    .ZN(_14259_));
 AOI21_X1 _40538_ (.A(_14181_),
    .B1(_14258_),
    .B2(_14259_),
    .ZN(_14260_));
 OR2_X4 _40539_ (.A1(_14257_),
    .A2(_14260_),
    .ZN(_14261_));
 BUF_X8 _40540_ (.A(_13472_),
    .Z(_14262_));
 NAND2_X1 _40541_ (.A1(_14227_),
    .A2(_13078_),
    .ZN(_14263_));
 OAI21_X1 _40542_ (.A(_13074_),
    .B1(_14240_),
    .B2(_14241_),
    .ZN(_14264_));
 AOI21_X1 _40543_ (.A(_14262_),
    .B1(_14263_),
    .B2(_14264_),
    .ZN(_14265_));
 NAND2_X1 _40544_ (.A1(_14200_),
    .A2(_13086_),
    .ZN(_14266_));
 OAI21_X2 _40545_ (.A(_13083_),
    .B1(_14216_),
    .B2(_14217_),
    .ZN(_14267_));
 AOI21_X2 _40546_ (.A(_14123_),
    .B1(_14266_),
    .B2(_14267_),
    .ZN(_14268_));
 OR2_X4 _40547_ (.A1(_14265_),
    .A2(_14268_),
    .ZN(_14269_));
 MUX2_X2 _40548_ (.A(_14261_),
    .B(_14269_),
    .S(_14111_),
    .Z(\icache.data_mem_data_li [118]));
 NAND2_X1 _40549_ (.A1(_14227_),
    .A2(_13110_),
    .ZN(_14270_));
 OAI21_X1 _40550_ (.A(_13107_),
    .B1(_14240_),
    .B2(_14241_),
    .ZN(_14271_));
 AOI21_X1 _40551_ (.A(_14160_),
    .B1(_14270_),
    .B2(_14271_),
    .ZN(_14272_));
 NAND2_X1 _40552_ (.A1(_14227_),
    .A2(_13117_),
    .ZN(_14273_));
 OAI21_X1 _40553_ (.A(_13114_),
    .B1(_14240_),
    .B2(_14241_),
    .ZN(_14274_));
 AOI21_X1 _40554_ (.A(_14181_),
    .B1(_14273_),
    .B2(_14274_),
    .ZN(_14275_));
 OR2_X4 _40555_ (.A1(_14272_),
    .A2(_14275_),
    .ZN(_14276_));
 BUF_X4 _40556_ (.A(_08490_),
    .Z(_14277_));
 NAND2_X1 _40557_ (.A1(_14277_),
    .A2(_13125_),
    .ZN(_14278_));
 OAI21_X1 _40558_ (.A(_13122_),
    .B1(_14216_),
    .B2(_14217_),
    .ZN(_14279_));
 AOI21_X1 _40559_ (.A(_14262_),
    .B1(_14278_),
    .B2(_14279_),
    .ZN(_14280_));
 BUF_X8 _40560_ (.A(_13494_),
    .Z(_14281_));
 NAND2_X1 _40561_ (.A1(_14277_),
    .A2(_13134_),
    .ZN(_14282_));
 OAI21_X1 _40562_ (.A(_13131_),
    .B1(_14216_),
    .B2(_14217_),
    .ZN(_14283_));
 AOI21_X1 _40563_ (.A(_14281_),
    .B1(_14282_),
    .B2(_14283_),
    .ZN(_14284_));
 OR2_X4 _40564_ (.A1(_14280_),
    .A2(_14284_),
    .ZN(_14285_));
 MUX2_X2 _40565_ (.A(_14276_),
    .B(_14285_),
    .S(_14111_),
    .Z(\icache.data_mem_data_li [119]));
 NAND2_X1 _40566_ (.A1(_14277_),
    .A2(_13143_),
    .ZN(_14286_));
 BUF_X8 _40567_ (.A(_11269_),
    .Z(_14287_));
 BUF_X8 _40568_ (.A(_11271_),
    .Z(_14288_));
 OAI21_X2 _40569_ (.A(_13140_),
    .B1(_14287_),
    .B2(_14288_),
    .ZN(_14289_));
 AOI21_X2 _40570_ (.A(_14160_),
    .B1(_14286_),
    .B2(_14289_),
    .ZN(_14290_));
 NAND2_X1 _40571_ (.A1(_14227_),
    .A2(_13152_),
    .ZN(_14291_));
 OAI21_X1 _40572_ (.A(_13149_),
    .B1(_14240_),
    .B2(_14241_),
    .ZN(_14292_));
 AOI21_X1 _40573_ (.A(_14181_),
    .B1(_14291_),
    .B2(_14292_),
    .ZN(_14293_));
 OR2_X4 _40574_ (.A1(_14290_),
    .A2(_14293_),
    .ZN(_14294_));
 NAND2_X1 _40575_ (.A1(_14227_),
    .A2(_13160_),
    .ZN(_14295_));
 OAI21_X1 _40576_ (.A(_13157_),
    .B1(_14240_),
    .B2(_14241_),
    .ZN(_14296_));
 AOI21_X1 _40577_ (.A(_14262_),
    .B1(_14295_),
    .B2(_14296_),
    .ZN(_14297_));
 NAND2_X1 _40578_ (.A1(_14277_),
    .A2(_13167_),
    .ZN(_14298_));
 OAI21_X1 _40579_ (.A(_13164_),
    .B1(_14287_),
    .B2(_14288_),
    .ZN(_14299_));
 AOI21_X1 _40580_ (.A(_14281_),
    .B1(_14298_),
    .B2(_14299_),
    .ZN(_14300_));
 OR2_X4 _40581_ (.A1(_14297_),
    .A2(_14300_),
    .ZN(_14301_));
 MUX2_X2 _40582_ (.A(_14294_),
    .B(_14301_),
    .S(_14111_),
    .Z(\icache.data_mem_data_li [120]));
 NAND2_X1 _40583_ (.A1(_14277_),
    .A2(_13195_),
    .ZN(_14302_));
 OAI21_X2 _40584_ (.A(_13192_),
    .B1(_14287_),
    .B2(_14288_),
    .ZN(_14303_));
 AOI21_X1 _40585_ (.A(_14160_),
    .B1(_14302_),
    .B2(_14303_),
    .ZN(_14304_));
 BUF_X4 _40586_ (.A(_08489_),
    .Z(_14305_));
 NAND2_X1 _40587_ (.A1(_14305_),
    .A2(_13202_),
    .ZN(_14306_));
 OAI21_X1 _40588_ (.A(_13199_),
    .B1(_14240_),
    .B2(_14241_),
    .ZN(_14307_));
 AOI21_X1 _40589_ (.A(_14181_),
    .B1(_14306_),
    .B2(_14307_),
    .ZN(_14308_));
 OR2_X4 _40590_ (.A1(_14304_),
    .A2(_14308_),
    .ZN(_14309_));
 NAND2_X1 _40591_ (.A1(_14305_),
    .A2(_13177_),
    .ZN(_14310_));
 OAI21_X1 _40592_ (.A(_13174_),
    .B1(_14240_),
    .B2(_14241_),
    .ZN(_14311_));
 AOI21_X1 _40593_ (.A(_14262_),
    .B1(_14310_),
    .B2(_14311_),
    .ZN(_14312_));
 NAND2_X1 _40594_ (.A1(_14277_),
    .A2(_13187_),
    .ZN(_14313_));
 OAI21_X1 _40595_ (.A(_13184_),
    .B1(_14287_),
    .B2(_14288_),
    .ZN(_14314_));
 AOI21_X1 _40596_ (.A(_14281_),
    .B1(_14313_),
    .B2(_14314_),
    .ZN(_14315_));
 OR2_X4 _40597_ (.A1(_14312_),
    .A2(_14315_),
    .ZN(_14316_));
 MUX2_X2 _40598_ (.A(_14309_),
    .B(_14316_),
    .S(_14048_),
    .Z(\icache.data_mem_data_li [121]));
 BUF_X8 _40599_ (.A(_14159_),
    .Z(_14317_));
 NAND2_X1 _40600_ (.A1(_14277_),
    .A2(_13227_),
    .ZN(_14318_));
 OAI21_X1 _40601_ (.A(_13224_),
    .B1(_14287_),
    .B2(_14288_),
    .ZN(_14319_));
 AOI21_X1 _40602_ (.A(_14317_),
    .B1(_14318_),
    .B2(_14319_),
    .ZN(_14320_));
 NAND2_X1 _40603_ (.A1(_14305_),
    .A2(_13234_),
    .ZN(_14321_));
 BUF_X4 _40604_ (.A(_08483_),
    .Z(_14322_));
 BUF_X4 _40605_ (.A(_08487_),
    .Z(_14323_));
 OAI21_X1 _40606_ (.A(_13231_),
    .B1(_14322_),
    .B2(_14323_),
    .ZN(_14324_));
 AOI21_X1 _40607_ (.A(_14181_),
    .B1(_14321_),
    .B2(_14324_),
    .ZN(_14325_));
 OR2_X4 _40608_ (.A1(_14320_),
    .A2(_14325_),
    .ZN(_14326_));
 NAND2_X1 _40609_ (.A1(_14305_),
    .A2(_13210_),
    .ZN(_14327_));
 OAI21_X2 _40610_ (.A(_13207_),
    .B1(_14322_),
    .B2(_14323_),
    .ZN(_14328_));
 AOI21_X2 _40611_ (.A(_14262_),
    .B1(_14327_),
    .B2(_14328_),
    .ZN(_14329_));
 NAND2_X1 _40612_ (.A1(_14277_),
    .A2(_13218_),
    .ZN(_14330_));
 OAI21_X2 _40613_ (.A(_13214_),
    .B1(_14287_),
    .B2(_14288_),
    .ZN(_14331_));
 AOI21_X1 _40614_ (.A(_14281_),
    .B1(_14330_),
    .B2(_14331_),
    .ZN(_14332_));
 OR2_X4 _40615_ (.A1(_14329_),
    .A2(_14332_),
    .ZN(_14333_));
 MUX2_X2 _40616_ (.A(_14326_),
    .B(_14333_),
    .S(_14048_),
    .Z(\icache.data_mem_data_li [122]));
 NAND2_X1 _40617_ (.A1(_14305_),
    .A2(_13242_),
    .ZN(_14334_));
 OAI21_X1 _40618_ (.A(_13239_),
    .B1(_14322_),
    .B2(_14323_),
    .ZN(_14335_));
 AOI21_X1 _40619_ (.A(_14317_),
    .B1(_14334_),
    .B2(_14335_),
    .ZN(_14336_));
 BUF_X8 _40620_ (.A(_14180_),
    .Z(_14337_));
 NAND2_X1 _40621_ (.A1(_14305_),
    .A2(_13250_),
    .ZN(_14338_));
 OAI21_X1 _40622_ (.A(_13246_),
    .B1(_14322_),
    .B2(_14323_),
    .ZN(_14339_));
 AOI21_X1 _40623_ (.A(_14337_),
    .B1(_14338_),
    .B2(_14339_),
    .ZN(_14340_));
 OR2_X4 _40624_ (.A1(_14336_),
    .A2(_14340_),
    .ZN(_14341_));
 NAND2_X1 _40625_ (.A1(_14277_),
    .A2(_13260_),
    .ZN(_14342_));
 OAI21_X2 _40626_ (.A(_13256_),
    .B1(_14287_),
    .B2(_14288_),
    .ZN(_14343_));
 AOI21_X2 _40627_ (.A(_14262_),
    .B1(_14342_),
    .B2(_14343_),
    .ZN(_14344_));
 NAND2_X1 _40628_ (.A1(_14277_),
    .A2(_13268_),
    .ZN(_14345_));
 OAI21_X2 _40629_ (.A(_13265_),
    .B1(_14287_),
    .B2(_14288_),
    .ZN(_14346_));
 AOI21_X1 _40630_ (.A(_14281_),
    .B1(_14345_),
    .B2(_14346_),
    .ZN(_14347_));
 OR2_X4 _40631_ (.A1(_14344_),
    .A2(_14347_),
    .ZN(_14348_));
 MUX2_X2 _40632_ (.A(_14341_),
    .B(_14348_),
    .S(_14111_),
    .Z(\icache.data_mem_data_li [123]));
 NAND2_X1 _40633_ (.A1(_14305_),
    .A2(_13276_),
    .ZN(_14349_));
 OAI21_X1 _40634_ (.A(_13273_),
    .B1(_14322_),
    .B2(_14323_),
    .ZN(_14350_));
 AOI21_X1 _40635_ (.A(_14317_),
    .B1(_14349_),
    .B2(_14350_),
    .ZN(_14351_));
 NAND2_X1 _40636_ (.A1(_14305_),
    .A2(_13283_),
    .ZN(_14352_));
 OAI21_X1 _40637_ (.A(_13280_),
    .B1(_14322_),
    .B2(_14323_),
    .ZN(_14353_));
 AOI21_X1 _40638_ (.A(_14337_),
    .B1(_14352_),
    .B2(_14353_),
    .ZN(_14354_));
 OR2_X4 _40639_ (.A1(_14351_),
    .A2(_14354_),
    .ZN(_14355_));
 NAND2_X1 _40640_ (.A1(_11259_),
    .A2(_13291_),
    .ZN(_14356_));
 OAI21_X1 _40641_ (.A(_13288_),
    .B1(_14287_),
    .B2(_14288_),
    .ZN(_14357_));
 AOI21_X1 _40642_ (.A(_14262_),
    .B1(_14356_),
    .B2(_14357_),
    .ZN(_14358_));
 NAND2_X1 _40643_ (.A1(_11259_),
    .A2(_13301_),
    .ZN(_14359_));
 OAI21_X1 _40644_ (.A(_13298_),
    .B1(_14287_),
    .B2(_14288_),
    .ZN(_14360_));
 AOI21_X1 _40645_ (.A(_14281_),
    .B1(_14359_),
    .B2(_14360_),
    .ZN(_14361_));
 OR2_X4 _40646_ (.A1(_14358_),
    .A2(_14361_),
    .ZN(_14362_));
 BUF_X32 _40647_ (.A(_12640_),
    .Z(_14363_));
 MUX2_X2 _40648_ (.A(_14355_),
    .B(_14362_),
    .S(_14363_),
    .Z(\icache.data_mem_data_li [124]));
 NAND2_X1 _40649_ (.A1(_11259_),
    .A2(_13309_),
    .ZN(_14364_));
 OAI21_X2 _40650_ (.A(_13306_),
    .B1(_11270_),
    .B2(_11272_),
    .ZN(_14365_));
 AOI21_X1 _40651_ (.A(_14317_),
    .B1(_14364_),
    .B2(_14365_),
    .ZN(_14366_));
 NAND2_X1 _40652_ (.A1(_14305_),
    .A2(_13317_),
    .ZN(_14367_));
 OAI21_X1 _40653_ (.A(_13314_),
    .B1(_14322_),
    .B2(_14323_),
    .ZN(_14368_));
 AOI21_X1 _40654_ (.A(_14337_),
    .B1(_14367_),
    .B2(_14368_),
    .ZN(_14369_));
 OR2_X4 _40655_ (.A1(_14366_),
    .A2(_14369_),
    .ZN(_14370_));
 NAND2_X1 _40656_ (.A1(_14305_),
    .A2(_13325_),
    .ZN(_14371_));
 OAI21_X2 _40657_ (.A(_13322_),
    .B1(_14322_),
    .B2(_14323_),
    .ZN(_14372_));
 AOI21_X1 _40658_ (.A(_14262_),
    .B1(_14371_),
    .B2(_14372_),
    .ZN(_14373_));
 NAND2_X1 _40659_ (.A1(_11259_),
    .A2(_13332_),
    .ZN(_14374_));
 OAI21_X2 _40660_ (.A(_13329_),
    .B1(_11270_),
    .B2(_11272_),
    .ZN(_14375_));
 AOI21_X1 _40661_ (.A(_14281_),
    .B1(_14374_),
    .B2(_14375_),
    .ZN(_14376_));
 OR2_X4 _40662_ (.A1(_14373_),
    .A2(_14376_),
    .ZN(_14377_));
 MUX2_X2 _40663_ (.A(_14370_),
    .B(_14377_),
    .S(_14363_),
    .Z(\icache.data_mem_data_li [125]));
 NAND2_X1 _40664_ (.A1(_11413_),
    .A2(_13341_),
    .ZN(_14378_));
 OAI21_X1 _40665_ (.A(_13338_),
    .B1(_14322_),
    .B2(_14323_),
    .ZN(_14379_));
 AOI21_X1 _40666_ (.A(_14317_),
    .B1(_14378_),
    .B2(_14379_),
    .ZN(_14380_));
 NAND2_X1 _40667_ (.A1(_11413_),
    .A2(_13352_),
    .ZN(_14381_));
 OAI21_X1 _40668_ (.A(_13349_),
    .B1(_14322_),
    .B2(_14323_),
    .ZN(_14382_));
 AOI21_X1 _40669_ (.A(_14337_),
    .B1(_14381_),
    .B2(_14382_),
    .ZN(_14383_));
 OR2_X4 _40670_ (.A1(_14380_),
    .A2(_14383_),
    .ZN(_14384_));
 NAND2_X1 _40671_ (.A1(_11259_),
    .A2(_13360_),
    .ZN(_14385_));
 OAI21_X2 _40672_ (.A(_13357_),
    .B1(_11270_),
    .B2(_11272_),
    .ZN(_14386_));
 AOI21_X2 _40673_ (.A(_14262_),
    .B1(_14385_),
    .B2(_14386_),
    .ZN(_14387_));
 NAND2_X1 _40674_ (.A1(_11259_),
    .A2(_13367_),
    .ZN(_14388_));
 OAI21_X1 _40675_ (.A(_13364_),
    .B1(_11270_),
    .B2(_11272_),
    .ZN(_14389_));
 AOI21_X1 _40676_ (.A(_14281_),
    .B1(_14388_),
    .B2(_14389_),
    .ZN(_14390_));
 OR2_X4 _40677_ (.A1(_14387_),
    .A2(_14390_),
    .ZN(_14391_));
 MUX2_X2 _40678_ (.A(_14384_),
    .B(_14391_),
    .S(_14363_),
    .Z(\icache.data_mem_data_li [126]));
 NAND2_X1 _40679_ (.A1(_11413_),
    .A2(_13375_),
    .ZN(_14392_));
 OAI21_X1 _40680_ (.A(_13372_),
    .B1(_11251_),
    .B2(_11253_),
    .ZN(_14393_));
 AOI21_X1 _40681_ (.A(_14317_),
    .B1(_14392_),
    .B2(_14393_),
    .ZN(_14394_));
 NAND2_X1 _40682_ (.A1(_11413_),
    .A2(_13383_),
    .ZN(_14395_));
 OAI21_X1 _40683_ (.A(_13380_),
    .B1(_11251_),
    .B2(_11253_),
    .ZN(_14396_));
 AOI21_X1 _40684_ (.A(_14337_),
    .B1(_14395_),
    .B2(_14396_),
    .ZN(_14397_));
 OR2_X4 _40685_ (.A1(_14394_),
    .A2(_14397_),
    .ZN(_14398_));
 NAND2_X1 _40686_ (.A1(_11259_),
    .A2(_13391_),
    .ZN(_14399_));
 OAI21_X1 _40687_ (.A(_13388_),
    .B1(_11270_),
    .B2(_11272_),
    .ZN(_14400_));
 AOI21_X1 _40688_ (.A(_14262_),
    .B1(_14399_),
    .B2(_14400_),
    .ZN(_14401_));
 NAND2_X1 _40689_ (.A1(_11259_),
    .A2(_13398_),
    .ZN(_14402_));
 OAI21_X2 _40690_ (.A(_13395_),
    .B1(_11270_),
    .B2(_11272_),
    .ZN(_14403_));
 AOI21_X1 _40691_ (.A(_14281_),
    .B1(_14402_),
    .B2(_14403_),
    .ZN(_14404_));
 OR2_X4 _40692_ (.A1(_14401_),
    .A2(_14404_),
    .ZN(_14405_));
 MUX2_X2 _40693_ (.A(_14398_),
    .B(_14405_),
    .S(_14048_),
    .Z(\icache.data_mem_data_li [127]));
 AOI21_X1 _40694_ (.A(_14317_),
    .B1(_11286_),
    .B2(_11289_),
    .ZN(_14406_));
 AOI21_X1 _40695_ (.A(_14337_),
    .B1(_11279_),
    .B2(_11282_),
    .ZN(_14407_));
 OR2_X1 _40696_ (.A1(_14406_),
    .A2(_14407_),
    .ZN(_14408_));
 BUF_X8 _40697_ (.A(_13472_),
    .Z(_14409_));
 AOI21_X1 _40698_ (.A(_14409_),
    .B1(_11262_),
    .B2(_11273_),
    .ZN(_14410_));
 AOI21_X1 _40699_ (.A(_14281_),
    .B1(_11247_),
    .B2(_11255_),
    .ZN(_14411_));
 OR2_X1 _40700_ (.A1(_14410_),
    .A2(_14411_),
    .ZN(_14412_));
 MUX2_X2 _40701_ (.A(_14408_),
    .B(_14412_),
    .S(_14363_),
    .Z(\icache.data_mem_data_li [128]));
 AOI21_X1 _40702_ (.A(_14317_),
    .B1(_11322_),
    .B2(_11325_),
    .ZN(_14413_));
 AOI21_X1 _40703_ (.A(_14337_),
    .B1(_11315_),
    .B2(_11318_),
    .ZN(_14414_));
 OR2_X2 _40704_ (.A1(_14413_),
    .A2(_14414_),
    .ZN(_14415_));
 AOI21_X1 _40705_ (.A(_14409_),
    .B1(_11305_),
    .B2(_11308_),
    .ZN(_14416_));
 BUF_X8 _40706_ (.A(_13494_),
    .Z(_14417_));
 AOI21_X1 _40707_ (.A(_14417_),
    .B1(_11296_),
    .B2(_11299_),
    .ZN(_14418_));
 OR2_X2 _40708_ (.A1(_14416_),
    .A2(_14418_),
    .ZN(_14419_));
 MUX2_X2 _40709_ (.A(_14415_),
    .B(_14419_),
    .S(_14048_),
    .Z(\icache.data_mem_data_li [129]));
 AOI21_X1 _40710_ (.A(_14317_),
    .B1(_11341_),
    .B2(_11344_),
    .ZN(_14420_));
 AOI21_X1 _40711_ (.A(_14337_),
    .B1(_11332_),
    .B2(_11337_),
    .ZN(_14421_));
 OR2_X1 _40712_ (.A1(_14420_),
    .A2(_14421_),
    .ZN(_14422_));
 AOI21_X1 _40713_ (.A(_14409_),
    .B1(_11357_),
    .B2(_11361_),
    .ZN(_14423_));
 AOI21_X1 _40714_ (.A(_14417_),
    .B1(_11350_),
    .B2(_11353_),
    .ZN(_14424_));
 OR2_X1 _40715_ (.A1(_14423_),
    .A2(_14424_),
    .ZN(_14425_));
 MUX2_X2 _40716_ (.A(_14422_),
    .B(_14425_),
    .S(_14363_),
    .Z(\icache.data_mem_data_li [130]));
 AOI21_X1 _40717_ (.A(_14317_),
    .B1(_11375_),
    .B2(_11378_),
    .ZN(_14426_));
 AOI21_X1 _40718_ (.A(_14337_),
    .B1(_11366_),
    .B2(_11369_),
    .ZN(_14427_));
 OR2_X1 _40719_ (.A1(_14426_),
    .A2(_14427_),
    .ZN(_14428_));
 AOI21_X1 _40720_ (.A(_14409_),
    .B1(_11390_),
    .B2(_11393_),
    .ZN(_14429_));
 AOI21_X1 _40721_ (.A(_14417_),
    .B1(_11383_),
    .B2(_11386_),
    .ZN(_14430_));
 OR2_X1 _40722_ (.A1(_14429_),
    .A2(_14430_),
    .ZN(_14431_));
 MUX2_X2 _40723_ (.A(_14428_),
    .B(_14431_),
    .S(_14363_),
    .Z(\icache.data_mem_data_li [131]));
 BUF_X8 _40724_ (.A(_14159_),
    .Z(_14432_));
 AOI21_X1 _40725_ (.A(_14432_),
    .B1(_11407_),
    .B2(_11410_),
    .ZN(_14433_));
 AOI21_X1 _40726_ (.A(_14337_),
    .B1(_11398_),
    .B2(_11402_),
    .ZN(_14434_));
 OR2_X1 _40727_ (.A1(_14433_),
    .A2(_14434_),
    .ZN(_14435_));
 AOI21_X1 _40728_ (.A(_14409_),
    .B1(_11424_),
    .B2(_11427_),
    .ZN(_14436_));
 AOI21_X1 _40729_ (.A(_14417_),
    .B1(_11417_),
    .B2(_11420_),
    .ZN(_14437_));
 OR2_X1 _40730_ (.A1(_14436_),
    .A2(_14437_),
    .ZN(_14438_));
 MUX2_X2 _40731_ (.A(_14435_),
    .B(_14438_),
    .S(_14363_),
    .Z(\icache.data_mem_data_li [132]));
 AOI21_X1 _40732_ (.A(_14432_),
    .B1(_11458_),
    .B2(_11461_),
    .ZN(_14439_));
 BUF_X16 _40733_ (.A(_14180_),
    .Z(_14440_));
 AOI21_X1 _40734_ (.A(_14440_),
    .B1(_11451_),
    .B2(_11454_),
    .ZN(_14441_));
 OR2_X2 _40735_ (.A1(_14439_),
    .A2(_14441_),
    .ZN(_14442_));
 AOI21_X1 _40736_ (.A(_14409_),
    .B1(_11442_),
    .B2(_11445_),
    .ZN(_14443_));
 AOI21_X1 _40737_ (.A(_14417_),
    .B1(_11432_),
    .B2(_11438_),
    .ZN(_14444_));
 OR2_X2 _40738_ (.A1(_14443_),
    .A2(_14444_),
    .ZN(_14445_));
 MUX2_X2 _40739_ (.A(_14442_),
    .B(_14445_),
    .S(_14048_),
    .Z(\icache.data_mem_data_li [133]));
 AOI21_X1 _40740_ (.A(_14432_),
    .B1(_11491_),
    .B2(_11494_),
    .ZN(_14446_));
 AOI21_X1 _40741_ (.A(_14440_),
    .B1(_11484_),
    .B2(_11487_),
    .ZN(_14447_));
 OR2_X4 _40742_ (.A1(_14446_),
    .A2(_14447_),
    .ZN(_14448_));
 AOI21_X1 _40743_ (.A(_14409_),
    .B1(_11476_),
    .B2(_11479_),
    .ZN(_14449_));
 AOI21_X1 _40744_ (.A(_14417_),
    .B1(_11466_),
    .B2(_11470_),
    .ZN(_14450_));
 OR2_X4 _40745_ (.A1(_14449_),
    .A2(_14450_),
    .ZN(_14451_));
 BUF_X8 _40746_ (.A(_13481_),
    .Z(_14452_));
 MUX2_X2 _40747_ (.A(_14448_),
    .B(_14451_),
    .S(_14452_),
    .Z(\icache.data_mem_data_li [134]));
 AOI21_X1 _40748_ (.A(_14432_),
    .B1(_11524_),
    .B2(_11527_),
    .ZN(_14453_));
 AOI21_X1 _40749_ (.A(_14440_),
    .B1(_11517_),
    .B2(_11520_),
    .ZN(_14454_));
 OR2_X1 _40750_ (.A1(_14453_),
    .A2(_14454_),
    .ZN(_14455_));
 AOI21_X1 _40751_ (.A(_14409_),
    .B1(_11506_),
    .B2(_11512_),
    .ZN(_14456_));
 AOI21_X1 _40752_ (.A(_14417_),
    .B1(_11499_),
    .B2(_11502_),
    .ZN(_14457_));
 OR2_X1 _40753_ (.A1(_14456_),
    .A2(_14457_),
    .ZN(_14458_));
 MUX2_X2 _40754_ (.A(_14455_),
    .B(_14458_),
    .S(_14363_),
    .Z(\icache.data_mem_data_li [135]));
 AOI21_X1 _40755_ (.A(_14432_),
    .B1(_11557_),
    .B2(_11560_),
    .ZN(_14459_));
 AOI21_X1 _40756_ (.A(_14440_),
    .B1(_11550_),
    .B2(_11553_),
    .ZN(_14460_));
 OR2_X1 _40757_ (.A1(_14459_),
    .A2(_14460_),
    .ZN(_14461_));
 AOI21_X1 _40758_ (.A(_14409_),
    .B1(_11540_),
    .B2(_11543_),
    .ZN(_14462_));
 AOI21_X1 _40759_ (.A(_14417_),
    .B1(_11532_),
    .B2(_11536_),
    .ZN(_14463_));
 OR2_X1 _40760_ (.A1(_14462_),
    .A2(_14463_),
    .ZN(_14464_));
 MUX2_X2 _40761_ (.A(_14461_),
    .B(_14464_),
    .S(_14452_),
    .Z(\icache.data_mem_data_li [136]));
 AOI21_X1 _40762_ (.A(_14432_),
    .B1(_11592_),
    .B2(_11595_),
    .ZN(_14465_));
 AOI21_X1 _40763_ (.A(_14440_),
    .B1(_11584_),
    .B2(_11587_),
    .ZN(_14466_));
 OR2_X2 _40764_ (.A1(_14465_),
    .A2(_14466_),
    .ZN(_14467_));
 AOI21_X1 _40765_ (.A(_14409_),
    .B1(_11575_),
    .B2(_11579_),
    .ZN(_14468_));
 AOI21_X1 _40766_ (.A(_14417_),
    .B1(_11567_),
    .B2(_11570_),
    .ZN(_14469_));
 OR2_X2 _40767_ (.A1(_14468_),
    .A2(_14469_),
    .ZN(_14470_));
 MUX2_X2 _40768_ (.A(_14467_),
    .B(_14470_),
    .S(_14363_),
    .Z(\icache.data_mem_data_li [137]));
 AOI21_X1 _40769_ (.A(_14432_),
    .B1(_11608_),
    .B2(_11611_),
    .ZN(_14471_));
 AOI21_X1 _40770_ (.A(_14440_),
    .B1(_11600_),
    .B2(_11604_),
    .ZN(_14472_));
 OR2_X1 _40771_ (.A1(_14471_),
    .A2(_14472_),
    .ZN(_14473_));
 BUF_X8 _40772_ (.A(_13472_),
    .Z(_14474_));
 AOI21_X1 _40773_ (.A(_14474_),
    .B1(_11625_),
    .B2(_11628_),
    .ZN(_14475_));
 AOI21_X1 _40774_ (.A(_14417_),
    .B1(_11616_),
    .B2(_11621_),
    .ZN(_14476_));
 OR2_X1 _40775_ (.A1(_14475_),
    .A2(_14476_),
    .ZN(_14477_));
 MUX2_X2 _40776_ (.A(_14473_),
    .B(_14477_),
    .S(_14452_),
    .Z(\icache.data_mem_data_li [138]));
 AOI21_X1 _40777_ (.A(_14432_),
    .B1(_11659_),
    .B2(_11662_),
    .ZN(_14478_));
 AOI21_X1 _40778_ (.A(_14440_),
    .B1(_11652_),
    .B2(_11655_),
    .ZN(_14479_));
 OR2_X2 _40779_ (.A1(_14478_),
    .A2(_14479_),
    .ZN(_14480_));
 AOI21_X1 _40780_ (.A(_14474_),
    .B1(_11642_),
    .B2(_11647_),
    .ZN(_14481_));
 BUF_X8 _40781_ (.A(_13494_),
    .Z(_14482_));
 AOI21_X1 _40782_ (.A(_14482_),
    .B1(_11633_),
    .B2(_11636_),
    .ZN(_14483_));
 OR2_X1 _40783_ (.A1(_14481_),
    .A2(_14483_),
    .ZN(_14484_));
 MUX2_X2 _40784_ (.A(_14480_),
    .B(_14484_),
    .S(_14363_),
    .Z(\icache.data_mem_data_li [139]));
 AOI21_X1 _40785_ (.A(_14432_),
    .B1(_11696_),
    .B2(_11699_),
    .ZN(_14485_));
 AOI21_X1 _40786_ (.A(_14440_),
    .B1(_11689_),
    .B2(_11692_),
    .ZN(_14486_));
 OR2_X2 _40787_ (.A1(_14485_),
    .A2(_14486_),
    .ZN(_14487_));
 AOI21_X1 _40788_ (.A(_14474_),
    .B1(_11677_),
    .B2(_11684_),
    .ZN(_14488_));
 AOI21_X1 _40789_ (.A(_14482_),
    .B1(_11669_),
    .B2(_11673_),
    .ZN(_14489_));
 OR2_X2 _40790_ (.A1(_14488_),
    .A2(_14489_),
    .ZN(_14490_));
 MUX2_X2 _40791_ (.A(_14487_),
    .B(_14490_),
    .S(_14452_),
    .Z(\icache.data_mem_data_li [140]));
 AOI21_X1 _40792_ (.A(_14432_),
    .B1(_11730_),
    .B2(_11733_),
    .ZN(_14491_));
 AOI21_X1 _40793_ (.A(_14440_),
    .B1(_11723_),
    .B2(_11726_),
    .ZN(_14492_));
 OR2_X2 _40794_ (.A1(_14491_),
    .A2(_14492_),
    .ZN(_14493_));
 AOI21_X2 _40795_ (.A(_14474_),
    .B1(_11714_),
    .B2(_11717_),
    .ZN(_14494_));
 AOI21_X1 _40796_ (.A(_14482_),
    .B1(_11704_),
    .B2(_11707_),
    .ZN(_14495_));
 OR2_X4 _40797_ (.A1(_14494_),
    .A2(_14495_),
    .ZN(_14496_));
 MUX2_X2 _40798_ (.A(_14493_),
    .B(_14496_),
    .S(_14452_),
    .Z(\icache.data_mem_data_li [141]));
 BUF_X8 _40799_ (.A(_14159_),
    .Z(_14497_));
 AOI21_X1 _40800_ (.A(_14497_),
    .B1(_11746_),
    .B2(_11750_),
    .ZN(_14498_));
 AOI21_X1 _40801_ (.A(_14440_),
    .B1(_11738_),
    .B2(_11741_),
    .ZN(_14499_));
 OR2_X4 _40802_ (.A1(_14498_),
    .A2(_14499_),
    .ZN(_14500_));
 AOI21_X1 _40803_ (.A(_14474_),
    .B1(_11763_),
    .B2(_11766_),
    .ZN(_14501_));
 AOI21_X1 _40804_ (.A(_14482_),
    .B1(_11756_),
    .B2(_11759_),
    .ZN(_14502_));
 OR2_X4 _40805_ (.A1(_14501_),
    .A2(_14502_),
    .ZN(_14503_));
 BUF_X8 _40806_ (.A(_12640_),
    .Z(_14504_));
 MUX2_X2 _40807_ (.A(_14500_),
    .B(_14503_),
    .S(_14504_),
    .Z(\icache.data_mem_data_li [142]));
 AOI21_X1 _40808_ (.A(_14497_),
    .B1(_11797_),
    .B2(_11800_),
    .ZN(_14505_));
 BUF_X8 _40809_ (.A(_14180_),
    .Z(_14506_));
 AOI21_X1 _40810_ (.A(_14506_),
    .B1(_11790_),
    .B2(_11793_),
    .ZN(_14507_));
 OR2_X4 _40811_ (.A1(_14505_),
    .A2(_14507_),
    .ZN(_14508_));
 AOI21_X1 _40812_ (.A(_14474_),
    .B1(_11782_),
    .B2(_11785_),
    .ZN(_14509_));
 AOI21_X1 _40813_ (.A(_14482_),
    .B1(_11772_),
    .B2(_11778_),
    .ZN(_14510_));
 OR2_X4 _40814_ (.A1(_14509_),
    .A2(_14510_),
    .ZN(_14511_));
 MUX2_X2 _40815_ (.A(_14508_),
    .B(_14511_),
    .S(_14452_),
    .Z(\icache.data_mem_data_li [143]));
 AOI21_X1 _40816_ (.A(_14497_),
    .B1(_11829_),
    .B2(_11832_),
    .ZN(_14512_));
 AOI21_X1 _40817_ (.A(_14506_),
    .B1(_11822_),
    .B2(_11825_),
    .ZN(_14513_));
 OR2_X4 _40818_ (.A1(_14512_),
    .A2(_14513_),
    .ZN(_14514_));
 AOI21_X1 _40819_ (.A(_14474_),
    .B1(_11814_),
    .B2(_11817_),
    .ZN(_14515_));
 AOI21_X1 _40820_ (.A(_14482_),
    .B1(_11805_),
    .B2(_11808_),
    .ZN(_14516_));
 OR2_X4 _40821_ (.A1(_14515_),
    .A2(_14516_),
    .ZN(_14517_));
 MUX2_X2 _40822_ (.A(_14514_),
    .B(_14517_),
    .S(_14504_),
    .Z(\icache.data_mem_data_li [144]));
 AOI21_X1 _40823_ (.A(_14497_),
    .B1(_11864_),
    .B2(_11867_),
    .ZN(_14518_));
 AOI21_X1 _40824_ (.A(_14506_),
    .B1(_11857_),
    .B2(_11860_),
    .ZN(_14519_));
 OR2_X4 _40825_ (.A1(_14518_),
    .A2(_14519_),
    .ZN(_14520_));
 AOI21_X1 _40826_ (.A(_14474_),
    .B1(_11846_),
    .B2(_11852_),
    .ZN(_14521_));
 AOI21_X1 _40827_ (.A(_14482_),
    .B1(_11839_),
    .B2(_11842_),
    .ZN(_14522_));
 OR2_X4 _40828_ (.A1(_14521_),
    .A2(_14522_),
    .ZN(_14523_));
 MUX2_X2 _40829_ (.A(_14520_),
    .B(_14523_),
    .S(_14452_),
    .Z(\icache.data_mem_data_li [145]));
 AOI21_X1 _40830_ (.A(_14497_),
    .B1(_11879_),
    .B2(_11883_),
    .ZN(_14524_));
 AOI21_X1 _40831_ (.A(_14506_),
    .B1(_11872_),
    .B2(_11875_),
    .ZN(_14525_));
 OR2_X4 _40832_ (.A1(_14524_),
    .A2(_14525_),
    .ZN(_14526_));
 AOI21_X1 _40833_ (.A(_14474_),
    .B1(_11897_),
    .B2(_11900_),
    .ZN(_14527_));
 AOI21_X1 _40834_ (.A(_14482_),
    .B1(_11889_),
    .B2(_11892_),
    .ZN(_14528_));
 OR2_X4 _40835_ (.A1(_14527_),
    .A2(_14528_),
    .ZN(_14529_));
 MUX2_X2 _40836_ (.A(_14526_),
    .B(_14529_),
    .S(_14504_),
    .Z(\icache.data_mem_data_li [146]));
 AOI21_X1 _40837_ (.A(_14497_),
    .B1(_11912_),
    .B2(_11915_),
    .ZN(_14530_));
 AOI21_X1 _40838_ (.A(_14506_),
    .B1(_11905_),
    .B2(_11908_),
    .ZN(_14531_));
 OR2_X4 _40839_ (.A1(_14530_),
    .A2(_14531_),
    .ZN(_14532_));
 AOI21_X1 _40840_ (.A(_14474_),
    .B1(_11930_),
    .B2(_11933_),
    .ZN(_14533_));
 AOI21_X1 _40841_ (.A(_14482_),
    .B1(_11922_),
    .B2(_11925_),
    .ZN(_14534_));
 OR2_X4 _40842_ (.A1(_14533_),
    .A2(_14534_),
    .ZN(_14535_));
 MUX2_X2 _40843_ (.A(_14532_),
    .B(_14535_),
    .S(_14504_),
    .Z(\icache.data_mem_data_li [147]));
 AOI21_X1 _40844_ (.A(_14497_),
    .B1(_11964_),
    .B2(_11967_),
    .ZN(_14536_));
 AOI21_X1 _40845_ (.A(_14506_),
    .B1(_11957_),
    .B2(_11960_),
    .ZN(_14537_));
 OR2_X4 _40846_ (.A1(_14536_),
    .A2(_14537_),
    .ZN(_14538_));
 BUF_X8 _40847_ (.A(_13472_),
    .Z(_14539_));
 AOI21_X1 _40848_ (.A(_14539_),
    .B1(_11949_),
    .B2(_11952_),
    .ZN(_14540_));
 AOI21_X1 _40849_ (.A(_14482_),
    .B1(_11938_),
    .B2(_11944_),
    .ZN(_14541_));
 OR2_X4 _40850_ (.A1(_14540_),
    .A2(_14541_),
    .ZN(_14542_));
 MUX2_X2 _40851_ (.A(_14538_),
    .B(_14542_),
    .S(_14504_),
    .Z(\icache.data_mem_data_li [148]));
 AOI21_X1 _40852_ (.A(_14497_),
    .B1(_11981_),
    .B2(_11984_),
    .ZN(_14543_));
 AOI21_X1 _40853_ (.A(_14506_),
    .B1(_11973_),
    .B2(_11977_),
    .ZN(_14544_));
 OR2_X4 _40854_ (.A1(_14543_),
    .A2(_14544_),
    .ZN(_14545_));
 AOI21_X1 _40855_ (.A(_14539_),
    .B1(_11996_),
    .B2(_12000_),
    .ZN(_14546_));
 BUF_X8 _40856_ (.A(_13494_),
    .Z(_14547_));
 AOI21_X1 _40857_ (.A(_14547_),
    .B1(_11989_),
    .B2(_11992_),
    .ZN(_14548_));
 OR2_X4 _40858_ (.A1(_14546_),
    .A2(_14548_),
    .ZN(_14549_));
 MUX2_X2 _40859_ (.A(_14545_),
    .B(_14549_),
    .S(_14504_),
    .Z(\icache.data_mem_data_li [149]));
 AOI21_X1 _40860_ (.A(_14497_),
    .B1(_12015_),
    .B2(_12018_),
    .ZN(_14550_));
 AOI21_X1 _40861_ (.A(_14506_),
    .B1(_12006_),
    .B2(_12011_),
    .ZN(_14551_));
 OR2_X4 _40862_ (.A1(_14550_),
    .A2(_14551_),
    .ZN(_14552_));
 AOI21_X1 _40863_ (.A(_14539_),
    .B1(_12030_),
    .B2(_12033_),
    .ZN(_14553_));
 AOI21_X1 _40864_ (.A(_14547_),
    .B1(_12023_),
    .B2(_12026_),
    .ZN(_14554_));
 OR2_X4 _40865_ (.A1(_14553_),
    .A2(_14554_),
    .ZN(_14555_));
 MUX2_X2 _40866_ (.A(_14552_),
    .B(_14555_),
    .S(_14452_),
    .Z(\icache.data_mem_data_li [150]));
 AOI21_X1 _40867_ (.A(_14497_),
    .B1(_12047_),
    .B2(_12050_),
    .ZN(_14556_));
 AOI21_X1 _40868_ (.A(_14506_),
    .B1(_12039_),
    .B2(_12042_),
    .ZN(_14557_));
 OR2_X4 _40869_ (.A1(_14556_),
    .A2(_14557_),
    .ZN(_14558_));
 AOI21_X1 _40870_ (.A(_14539_),
    .B1(_12063_),
    .B2(_12066_),
    .ZN(_14559_));
 AOI21_X1 _40871_ (.A(_14547_),
    .B1(_12055_),
    .B2(_12058_),
    .ZN(_14560_));
 OR2_X4 _40872_ (.A1(_14559_),
    .A2(_14560_),
    .ZN(_14561_));
 MUX2_X2 _40873_ (.A(_14558_),
    .B(_14561_),
    .S(_14504_),
    .Z(\icache.data_mem_data_li [151]));
 BUF_X8 _40874_ (.A(_14159_),
    .Z(_14562_));
 AOI21_X1 _40875_ (.A(_14562_),
    .B1(_12097_),
    .B2(_12100_),
    .ZN(_14563_));
 AOI21_X1 _40876_ (.A(_14506_),
    .B1(_12090_),
    .B2(_12093_),
    .ZN(_14564_));
 OR2_X4 _40877_ (.A1(_14563_),
    .A2(_14564_),
    .ZN(_14565_));
 AOI21_X1 _40878_ (.A(_14539_),
    .B1(_12082_),
    .B2(_12085_),
    .ZN(_14566_));
 AOI21_X1 _40879_ (.A(_14547_),
    .B1(_12073_),
    .B2(_12076_),
    .ZN(_14567_));
 OR2_X4 _40880_ (.A1(_14566_),
    .A2(_14567_),
    .ZN(_14568_));
 MUX2_X2 _40881_ (.A(_14565_),
    .B(_14568_),
    .S(_14452_),
    .Z(\icache.data_mem_data_li [152]));
 AOI21_X1 _40882_ (.A(_14562_),
    .B1(_12112_),
    .B2(_12116_),
    .ZN(_14569_));
 BUF_X8 _40883_ (.A(_14180_),
    .Z(_14570_));
 AOI21_X1 _40884_ (.A(_14570_),
    .B1(_12105_),
    .B2(_12108_),
    .ZN(_14571_));
 OR2_X4 _40885_ (.A1(_14569_),
    .A2(_14571_),
    .ZN(_14572_));
 AOI21_X1 _40886_ (.A(_14539_),
    .B1(_12131_),
    .B2(_12134_),
    .ZN(_14573_));
 AOI21_X1 _40887_ (.A(_14547_),
    .B1(_12122_),
    .B2(_12127_),
    .ZN(_14574_));
 OR2_X2 _40888_ (.A1(_14573_),
    .A2(_14574_),
    .ZN(_14575_));
 MUX2_X2 _40889_ (.A(_14572_),
    .B(_14575_),
    .S(_14504_),
    .Z(\icache.data_mem_data_li [153]));
 AOI21_X1 _40890_ (.A(_14562_),
    .B1(_12148_),
    .B2(_12152_),
    .ZN(_14576_));
 AOI21_X1 _40891_ (.A(_14570_),
    .B1(_12140_),
    .B2(_12143_),
    .ZN(_14577_));
 OR2_X4 _40892_ (.A1(_14576_),
    .A2(_14577_),
    .ZN(_14578_));
 AOI21_X1 _40893_ (.A(_14539_),
    .B1(_12164_),
    .B2(_12167_),
    .ZN(_14579_));
 AOI21_X1 _40894_ (.A(_14547_),
    .B1(_12157_),
    .B2(_12160_),
    .ZN(_14580_));
 OR2_X2 _40895_ (.A1(_14579_),
    .A2(_14580_),
    .ZN(_14581_));
 MUX2_X2 _40896_ (.A(_14578_),
    .B(_14581_),
    .S(_14504_),
    .Z(\icache.data_mem_data_li [154]));
 AOI21_X1 _40897_ (.A(_14562_),
    .B1(_12181_),
    .B2(_12184_),
    .ZN(_14582_));
 AOI21_X1 _40898_ (.A(_14570_),
    .B1(_12172_),
    .B2(_12177_),
    .ZN(_14583_));
 OR2_X4 _40899_ (.A1(_14582_),
    .A2(_14583_),
    .ZN(_14584_));
 AOI21_X1 _40900_ (.A(_14539_),
    .B1(_12196_),
    .B2(_12200_),
    .ZN(_14585_));
 AOI21_X1 _40901_ (.A(_14547_),
    .B1(_12189_),
    .B2(_12192_),
    .ZN(_14586_));
 OR2_X2 _40902_ (.A1(_14585_),
    .A2(_14586_),
    .ZN(_14587_));
 MUX2_X2 _40903_ (.A(_14584_),
    .B(_14587_),
    .S(_14504_),
    .Z(\icache.data_mem_data_li [155]));
 AOI21_X1 _40904_ (.A(_14562_),
    .B1(_12214_),
    .B2(_12217_),
    .ZN(_14588_));
 AOI21_X1 _40905_ (.A(_14570_),
    .B1(_12206_),
    .B2(_12210_),
    .ZN(_14589_));
 OR2_X2 _40906_ (.A1(_14588_),
    .A2(_14589_),
    .ZN(_14590_));
 AOI21_X1 _40907_ (.A(_14539_),
    .B1(_12230_),
    .B2(_12233_),
    .ZN(_14591_));
 AOI21_X1 _40908_ (.A(_14547_),
    .B1(_12223_),
    .B2(_12226_),
    .ZN(_14592_));
 OR2_X2 _40909_ (.A1(_14591_),
    .A2(_14592_),
    .ZN(_14593_));
 BUF_X8 _40910_ (.A(_12640_),
    .Z(_14594_));
 MUX2_X2 _40911_ (.A(_14590_),
    .B(_14593_),
    .S(_14594_),
    .Z(\icache.data_mem_data_li [156]));
 AOI21_X1 _40912_ (.A(_14562_),
    .B1(_12264_),
    .B2(_12267_),
    .ZN(_14595_));
 AOI21_X1 _40913_ (.A(_14570_),
    .B1(_12256_),
    .B2(_12259_),
    .ZN(_14596_));
 OR2_X1 _40914_ (.A1(_14595_),
    .A2(_14596_),
    .ZN(_14597_));
 AOI21_X1 _40915_ (.A(_14539_),
    .B1(_12248_),
    .B2(_12251_),
    .ZN(_14598_));
 AOI21_X1 _40916_ (.A(_14547_),
    .B1(_12240_),
    .B2(_12243_),
    .ZN(_14599_));
 OR2_X1 _40917_ (.A1(_14598_),
    .A2(_14599_),
    .ZN(_14600_));
 MUX2_X2 _40918_ (.A(_14597_),
    .B(_14600_),
    .S(_14452_),
    .Z(\icache.data_mem_data_li [157]));
 AOI21_X1 _40919_ (.A(_14562_),
    .B1(_12279_),
    .B2(_12282_),
    .ZN(_14601_));
 AOI21_X1 _40920_ (.A(_14570_),
    .B1(_12272_),
    .B2(_12275_),
    .ZN(_14602_));
 OR2_X2 _40921_ (.A1(_14601_),
    .A2(_14602_),
    .ZN(_14603_));
 BUF_X8 _40922_ (.A(_13472_),
    .Z(_14604_));
 AOI21_X1 _40923_ (.A(_14604_),
    .B1(_12296_),
    .B2(_12301_),
    .ZN(_14605_));
 AOI21_X1 _40924_ (.A(_14547_),
    .B1(_12287_),
    .B2(_12292_),
    .ZN(_14606_));
 OR2_X2 _40925_ (.A1(_14605_),
    .A2(_14606_),
    .ZN(_14607_));
 MUX2_X2 _40926_ (.A(_14603_),
    .B(_14607_),
    .S(_14594_),
    .Z(\icache.data_mem_data_li [158]));
 AOI21_X1 _40927_ (.A(_14562_),
    .B1(_12316_),
    .B2(_12319_),
    .ZN(_14608_));
 AOI21_X1 _40928_ (.A(_14570_),
    .B1(_12308_),
    .B2(_12312_),
    .ZN(_14609_));
 OR2_X2 _40929_ (.A1(_14608_),
    .A2(_14609_),
    .ZN(_14610_));
 AOI21_X1 _40930_ (.A(_14604_),
    .B1(_12331_),
    .B2(_12334_),
    .ZN(_14611_));
 BUF_X8 _40931_ (.A(_13494_),
    .Z(_14612_));
 AOI21_X1 _40932_ (.A(_14612_),
    .B1(_12324_),
    .B2(_12327_),
    .ZN(_14613_));
 OR2_X1 _40933_ (.A1(_14611_),
    .A2(_14613_),
    .ZN(_14614_));
 BUF_X8 _40934_ (.A(_13481_),
    .Z(_14615_));
 MUX2_X2 _40935_ (.A(_14610_),
    .B(_14614_),
    .S(_14615_),
    .Z(\icache.data_mem_data_li [159]));
 AOI21_X1 _40936_ (.A(_14562_),
    .B1(_12367_),
    .B2(_12370_),
    .ZN(_14616_));
 AOI21_X1 _40937_ (.A(_14570_),
    .B1(_12360_),
    .B2(_12363_),
    .ZN(_14617_));
 OR2_X1 _40938_ (.A1(_14616_),
    .A2(_14617_),
    .ZN(_14618_));
 AOI21_X1 _40939_ (.A(_14604_),
    .B1(_12349_),
    .B2(_12355_),
    .ZN(_14619_));
 AOI21_X1 _40940_ (.A(_14612_),
    .B1(_12341_),
    .B2(_12345_),
    .ZN(_14620_));
 OR2_X1 _40941_ (.A1(_14619_),
    .A2(_14620_),
    .ZN(_14621_));
 MUX2_X2 _40942_ (.A(_14618_),
    .B(_14621_),
    .S(_14594_),
    .Z(\icache.data_mem_data_li [160]));
 AOI21_X1 _40943_ (.A(_14562_),
    .B1(_12399_),
    .B2(_12402_),
    .ZN(_14622_));
 AOI21_X1 _40944_ (.A(_14570_),
    .B1(_12392_),
    .B2(_12395_),
    .ZN(_14623_));
 OR2_X2 _40945_ (.A1(_14622_),
    .A2(_14623_),
    .ZN(_14624_));
 AOI21_X1 _40946_ (.A(_14604_),
    .B1(_12384_),
    .B2(_12387_),
    .ZN(_14625_));
 AOI21_X1 _40947_ (.A(_14612_),
    .B1(_12376_),
    .B2(_12379_),
    .ZN(_14626_));
 OR2_X2 _40948_ (.A1(_14625_),
    .A2(_14626_),
    .ZN(_14627_));
 MUX2_X2 _40949_ (.A(_14624_),
    .B(_14627_),
    .S(_14615_),
    .Z(\icache.data_mem_data_li [161]));
 BUF_X8 _40950_ (.A(_14159_),
    .Z(_14628_));
 AOI21_X1 _40951_ (.A(_14628_),
    .B1(_12415_),
    .B2(_12418_),
    .ZN(_14629_));
 AOI21_X1 _40952_ (.A(_14570_),
    .B1(_12408_),
    .B2(_12411_),
    .ZN(_14630_));
 OR2_X2 _40953_ (.A1(_14629_),
    .A2(_14630_),
    .ZN(_14631_));
 AOI21_X1 _40954_ (.A(_14604_),
    .B1(_12433_),
    .B2(_12436_),
    .ZN(_14632_));
 AOI21_X1 _40955_ (.A(_14612_),
    .B1(_12426_),
    .B2(_12429_),
    .ZN(_14633_));
 OR2_X2 _40956_ (.A1(_14632_),
    .A2(_14633_),
    .ZN(_14634_));
 MUX2_X2 _40957_ (.A(_14631_),
    .B(_14634_),
    .S(_14594_),
    .Z(\icache.data_mem_data_li [162]));
 AOI21_X1 _40958_ (.A(_14628_),
    .B1(_12449_),
    .B2(_12452_),
    .ZN(_14635_));
 BUF_X8 _40959_ (.A(_14180_),
    .Z(_14636_));
 AOI21_X1 _40960_ (.A(_14636_),
    .B1(_12442_),
    .B2(_12445_),
    .ZN(_14637_));
 OR2_X2 _40961_ (.A1(_14635_),
    .A2(_14637_),
    .ZN(_14638_));
 AOI21_X1 _40962_ (.A(_14604_),
    .B1(_12467_),
    .B2(_12470_),
    .ZN(_14639_));
 AOI21_X1 _40963_ (.A(_14612_),
    .B1(_12457_),
    .B2(_12462_),
    .ZN(_14640_));
 OR2_X1 _40964_ (.A1(_14639_),
    .A2(_14640_),
    .ZN(_14641_));
 MUX2_X2 _40965_ (.A(_14638_),
    .B(_14641_),
    .S(_14594_),
    .Z(\icache.data_mem_data_li [163]));
 AOI21_X1 _40966_ (.A(_14628_),
    .B1(_12485_),
    .B2(_12488_),
    .ZN(_14642_));
 AOI21_X1 _40967_ (.A(_14636_),
    .B1(_12476_),
    .B2(_12480_),
    .ZN(_14643_));
 OR2_X1 _40968_ (.A1(_14642_),
    .A2(_14643_),
    .ZN(_14644_));
 AOI21_X1 _40969_ (.A(_14604_),
    .B1(_12500_),
    .B2(_12503_),
    .ZN(_14645_));
 AOI21_X1 _40970_ (.A(_14612_),
    .B1(_12493_),
    .B2(_12496_),
    .ZN(_14646_));
 OR2_X1 _40971_ (.A1(_14645_),
    .A2(_14646_),
    .ZN(_14647_));
 MUX2_X2 _40972_ (.A(_14644_),
    .B(_14647_),
    .S(_14594_),
    .Z(\icache.data_mem_data_li [164]));
 AOI21_X1 _40973_ (.A(_14628_),
    .B1(_12533_),
    .B2(_12536_),
    .ZN(_14648_));
 AOI21_X1 _40974_ (.A(_14636_),
    .B1(_12526_),
    .B2(_12529_),
    .ZN(_14649_));
 OR2_X1 _40975_ (.A1(_14648_),
    .A2(_14649_),
    .ZN(_14650_));
 AOI21_X1 _40976_ (.A(_14604_),
    .B1(_12515_),
    .B2(_12521_),
    .ZN(_14651_));
 AOI21_X1 _40977_ (.A(_14612_),
    .B1(_12508_),
    .B2(_12511_),
    .ZN(_14652_));
 OR2_X1 _40978_ (.A1(_14651_),
    .A2(_14652_),
    .ZN(_14653_));
 MUX2_X2 _40979_ (.A(_14650_),
    .B(_14653_),
    .S(_14615_),
    .Z(\icache.data_mem_data_li [165]));
 AOI21_X1 _40980_ (.A(_14628_),
    .B1(_12565_),
    .B2(_12568_),
    .ZN(_14654_));
 AOI21_X1 _40981_ (.A(_14636_),
    .B1(_12558_),
    .B2(_12561_),
    .ZN(_14655_));
 OR2_X1 _40982_ (.A1(_14654_),
    .A2(_14655_),
    .ZN(_14656_));
 AOI21_X1 _40983_ (.A(_14604_),
    .B1(_12549_),
    .B2(_12552_),
    .ZN(_14657_));
 AOI21_X1 _40984_ (.A(_14612_),
    .B1(_12542_),
    .B2(_12545_),
    .ZN(_14658_));
 OR2_X1 _40985_ (.A1(_14657_),
    .A2(_14658_),
    .ZN(_14659_));
 MUX2_X2 _40986_ (.A(_14656_),
    .B(_14659_),
    .S(_14615_),
    .Z(\icache.data_mem_data_li [166]));
 AOI21_X1 _40987_ (.A(_14628_),
    .B1(_12599_),
    .B2(_12602_),
    .ZN(_14660_));
 AOI21_X1 _40988_ (.A(_14636_),
    .B1(_12591_),
    .B2(_12594_),
    .ZN(_14661_));
 OR2_X1 _40989_ (.A1(_14660_),
    .A2(_14661_),
    .ZN(_14662_));
 AOI21_X1 _40990_ (.A(_14604_),
    .B1(_12582_),
    .B2(_12586_),
    .ZN(_14663_));
 AOI21_X1 _40991_ (.A(_14612_),
    .B1(_12574_),
    .B2(_12578_),
    .ZN(_14664_));
 OR2_X1 _40992_ (.A1(_14663_),
    .A2(_14664_),
    .ZN(_14665_));
 MUX2_X2 _40993_ (.A(_14662_),
    .B(_14665_),
    .S(_14594_),
    .Z(\icache.data_mem_data_li [167]));
 AOI21_X1 _40994_ (.A(_14628_),
    .B1(_12634_),
    .B2(_12637_),
    .ZN(_14666_));
 AOI21_X1 _40995_ (.A(_14636_),
    .B1(_12627_),
    .B2(_12630_),
    .ZN(_14667_));
 OR2_X1 _40996_ (.A1(_14666_),
    .A2(_14667_),
    .ZN(_14668_));
 BUF_X4 _40997_ (.A(_11239_),
    .Z(_14669_));
 AOI21_X1 _40998_ (.A(_14669_),
    .B1(_12618_),
    .B2(_12622_),
    .ZN(_14670_));
 AOI21_X1 _40999_ (.A(_14612_),
    .B1(_12607_),
    .B2(_12614_),
    .ZN(_14671_));
 OR2_X1 _41000_ (.A1(_14670_),
    .A2(_14671_),
    .ZN(_14672_));
 MUX2_X2 _41001_ (.A(_14668_),
    .B(_14672_),
    .S(_14615_),
    .Z(\icache.data_mem_data_li [168]));
 AOI21_X1 _41002_ (.A(_14628_),
    .B1(_12669_),
    .B2(_12672_),
    .ZN(_14673_));
 AOI21_X1 _41003_ (.A(_14636_),
    .B1(_12662_),
    .B2(_12665_),
    .ZN(_14674_));
 OR2_X1 _41004_ (.A1(_14673_),
    .A2(_14674_),
    .ZN(_14675_));
 AOI21_X1 _41005_ (.A(_14669_),
    .B1(_12654_),
    .B2(_12657_),
    .ZN(_14676_));
 BUF_X8 _41006_ (.A(_11257_),
    .Z(_14677_));
 AOI21_X1 _41007_ (.A(_14677_),
    .B1(_12645_),
    .B2(_12649_),
    .ZN(_14678_));
 OR2_X1 _41008_ (.A1(_14676_),
    .A2(_14678_),
    .ZN(_14679_));
 MUX2_X2 _41009_ (.A(_14675_),
    .B(_14679_),
    .S(_14594_),
    .Z(\icache.data_mem_data_li [169]));
 AOI21_X1 _41010_ (.A(_14628_),
    .B1(_12689_),
    .B2(_12692_),
    .ZN(_14680_));
 AOI21_X1 _41011_ (.A(_14636_),
    .B1(_12678_),
    .B2(_12684_),
    .ZN(_14681_));
 OR2_X1 _41012_ (.A1(_14680_),
    .A2(_14681_),
    .ZN(_14682_));
 AOI21_X1 _41013_ (.A(_14669_),
    .B1(_12704_),
    .B2(_12707_),
    .ZN(_14683_));
 AOI21_X1 _41014_ (.A(_14677_),
    .B1(_12697_),
    .B2(_12700_),
    .ZN(_14684_));
 OR2_X1 _41015_ (.A1(_14683_),
    .A2(_14684_),
    .ZN(_14685_));
 MUX2_X2 _41016_ (.A(_14682_),
    .B(_14685_),
    .S(_14615_),
    .Z(\icache.data_mem_data_li [170]));
 AOI21_X1 _41017_ (.A(_14628_),
    .B1(_12736_),
    .B2(_12739_),
    .ZN(_14686_));
 AOI21_X1 _41018_ (.A(_14636_),
    .B1(_12729_),
    .B2(_12732_),
    .ZN(_14687_));
 OR2_X1 _41019_ (.A1(_14686_),
    .A2(_14687_),
    .ZN(_14688_));
 AOI21_X1 _41020_ (.A(_14669_),
    .B1(_12720_),
    .B2(_12724_),
    .ZN(_14689_));
 AOI21_X1 _41021_ (.A(_14677_),
    .B1(_12712_),
    .B2(_12715_),
    .ZN(_14690_));
 OR2_X1 _41022_ (.A1(_14689_),
    .A2(_14690_),
    .ZN(_14691_));
 MUX2_X2 _41023_ (.A(_14688_),
    .B(_14691_),
    .S(_14594_),
    .Z(\icache.data_mem_data_li [171]));
 BUF_X8 _41024_ (.A(_14159_),
    .Z(_14692_));
 AOI21_X1 _41025_ (.A(_14692_),
    .B1(_12768_),
    .B2(_12771_),
    .ZN(_14693_));
 AOI21_X1 _41026_ (.A(_14636_),
    .B1(_12761_),
    .B2(_12764_),
    .ZN(_14694_));
 OR2_X1 _41027_ (.A1(_14693_),
    .A2(_14694_),
    .ZN(_14695_));
 AOI21_X1 _41028_ (.A(_14669_),
    .B1(_12753_),
    .B2(_12756_),
    .ZN(_14696_));
 AOI21_X1 _41029_ (.A(_14677_),
    .B1(_12746_),
    .B2(_12749_),
    .ZN(_14697_));
 OR2_X1 _41030_ (.A1(_14696_),
    .A2(_14697_),
    .ZN(_14698_));
 MUX2_X2 _41031_ (.A(_14695_),
    .B(_14698_),
    .S(_14615_),
    .Z(\icache.data_mem_data_li [172]));
 AOI21_X1 _41032_ (.A(_14692_),
    .B1(_12802_),
    .B2(_12805_),
    .ZN(_14699_));
 BUF_X8 _41033_ (.A(_14180_),
    .Z(_14700_));
 AOI21_X1 _41034_ (.A(_14700_),
    .B1(_12795_),
    .B2(_12798_),
    .ZN(_14701_));
 OR2_X1 _41035_ (.A1(_14699_),
    .A2(_14701_),
    .ZN(_14702_));
 AOI21_X1 _41036_ (.A(_14669_),
    .B1(_12787_),
    .B2(_12790_),
    .ZN(_14703_));
 AOI21_X1 _41037_ (.A(_14677_),
    .B1(_12777_),
    .B2(_12782_),
    .ZN(_14704_));
 OR2_X1 _41038_ (.A1(_14703_),
    .A2(_14704_),
    .ZN(_14705_));
 MUX2_X2 _41039_ (.A(_14702_),
    .B(_14705_),
    .S(_14615_),
    .Z(\icache.data_mem_data_li [173]));
 AOI21_X1 _41040_ (.A(_14692_),
    .B1(_12819_),
    .B2(_12822_),
    .ZN(_14706_));
 AOI21_X1 _41041_ (.A(_14700_),
    .B1(_12812_),
    .B2(_12815_),
    .ZN(_14707_));
 OR2_X4 _41042_ (.A1(_14706_),
    .A2(_14707_),
    .ZN(_14708_));
 AOI21_X1 _41043_ (.A(_14669_),
    .B1(_12834_),
    .B2(_12837_),
    .ZN(_14709_));
 AOI21_X1 _41044_ (.A(_14677_),
    .B1(_12827_),
    .B2(_12830_),
    .ZN(_14710_));
 OR2_X2 _41045_ (.A1(_14709_),
    .A2(_14710_),
    .ZN(_14711_));
 MUX2_X2 _41046_ (.A(_14708_),
    .B(_14711_),
    .S(_14594_),
    .Z(\icache.data_mem_data_li [174]));
 AOI21_X1 _41047_ (.A(_14692_),
    .B1(_12867_),
    .B2(_12870_),
    .ZN(_14712_));
 AOI21_X1 _41048_ (.A(_14700_),
    .B1(_12860_),
    .B2(_12863_),
    .ZN(_14713_));
 OR2_X1 _41049_ (.A1(_14712_),
    .A2(_14713_),
    .ZN(_14714_));
 AOI21_X1 _41050_ (.A(_14669_),
    .B1(_12850_),
    .B2(_12855_),
    .ZN(_14715_));
 AOI21_X1 _41051_ (.A(_14677_),
    .B1(_12843_),
    .B2(_12846_),
    .ZN(_14716_));
 OR2_X1 _41052_ (.A1(_14715_),
    .A2(_14716_),
    .ZN(_14717_));
 MUX2_X2 _41053_ (.A(_14714_),
    .B(_14717_),
    .S(_14615_),
    .Z(\icache.data_mem_data_li [175]));
 AOI21_X1 _41054_ (.A(_14692_),
    .B1(_12900_),
    .B2(_12903_),
    .ZN(_14718_));
 AOI21_X1 _41055_ (.A(_14700_),
    .B1(_12893_),
    .B2(_12896_),
    .ZN(_14719_));
 OR2_X1 _41056_ (.A1(_14718_),
    .A2(_14719_),
    .ZN(_14720_));
 AOI21_X1 _41057_ (.A(_14669_),
    .B1(_12884_),
    .B2(_12887_),
    .ZN(_14721_));
 AOI21_X1 _41058_ (.A(_14677_),
    .B1(_12875_),
    .B2(_12879_),
    .ZN(_14722_));
 OR2_X1 _41059_ (.A1(_14721_),
    .A2(_14722_),
    .ZN(_14723_));
 BUF_X8 _41060_ (.A(_12640_),
    .Z(_14724_));
 MUX2_X2 _41061_ (.A(_14720_),
    .B(_14723_),
    .S(_14724_),
    .Z(\icache.data_mem_data_li [176]));
 AOI21_X1 _41062_ (.A(_14692_),
    .B1(_12934_),
    .B2(_12937_),
    .ZN(_14725_));
 AOI21_X1 _41063_ (.A(_14700_),
    .B1(_12926_),
    .B2(_12929_),
    .ZN(_14726_));
 OR2_X1 _41064_ (.A1(_14725_),
    .A2(_14726_),
    .ZN(_14727_));
 AOI21_X1 _41065_ (.A(_14669_),
    .B1(_12918_),
    .B2(_12921_),
    .ZN(_14728_));
 AOI21_X1 _41066_ (.A(_14677_),
    .B1(_12909_),
    .B2(_12913_),
    .ZN(_14729_));
 OR2_X1 _41067_ (.A1(_14728_),
    .A2(_14729_),
    .ZN(_14730_));
 MUX2_X2 _41068_ (.A(_14727_),
    .B(_14730_),
    .S(_14615_),
    .Z(\icache.data_mem_data_li [177]));
 AOI21_X1 _41069_ (.A(_14692_),
    .B1(_12949_),
    .B2(_12953_),
    .ZN(_14731_));
 AOI21_X1 _41070_ (.A(_14700_),
    .B1(_12942_),
    .B2(_12945_),
    .ZN(_14732_));
 OR2_X1 _41071_ (.A1(_14731_),
    .A2(_14732_),
    .ZN(_14733_));
 BUF_X8 _41072_ (.A(_11239_),
    .Z(_14734_));
 AOI21_X1 _41073_ (.A(_14734_),
    .B1(_12967_),
    .B2(_12970_),
    .ZN(_14735_));
 AOI21_X1 _41074_ (.A(_14677_),
    .B1(_12958_),
    .B2(_12963_),
    .ZN(_14736_));
 OR2_X1 _41075_ (.A1(_14735_),
    .A2(_14736_),
    .ZN(_14737_));
 MUX2_X2 _41076_ (.A(_14733_),
    .B(_14737_),
    .S(_14724_),
    .Z(\icache.data_mem_data_li [178]));
 AOI21_X1 _41077_ (.A(_14692_),
    .B1(_12984_),
    .B2(_12988_),
    .ZN(_14738_));
 AOI21_X1 _41078_ (.A(_14700_),
    .B1(_12977_),
    .B2(_12980_),
    .ZN(_14739_));
 OR2_X2 _41079_ (.A1(_14738_),
    .A2(_14739_),
    .ZN(_14740_));
 AOI21_X1 _41080_ (.A(_14734_),
    .B1(_13001_),
    .B2(_13004_),
    .ZN(_14741_));
 BUF_X8 _41081_ (.A(_11257_),
    .Z(_14742_));
 AOI21_X1 _41082_ (.A(_14742_),
    .B1(_12993_),
    .B2(_12997_),
    .ZN(_14743_));
 OR2_X1 _41083_ (.A1(_14741_),
    .A2(_14743_),
    .ZN(_14744_));
 MUX2_X2 _41084_ (.A(_14740_),
    .B(_14744_),
    .S(_14724_),
    .Z(\icache.data_mem_data_li [179]));
 AOI21_X1 _41085_ (.A(_14692_),
    .B1(_13034_),
    .B2(_13037_),
    .ZN(_14745_));
 AOI21_X1 _41086_ (.A(_14700_),
    .B1(_13027_),
    .B2(_13030_),
    .ZN(_14746_));
 OR2_X1 _41087_ (.A1(_14745_),
    .A2(_14746_),
    .ZN(_14747_));
 AOI21_X1 _41088_ (.A(_14734_),
    .B1(_13017_),
    .B2(_13022_),
    .ZN(_14748_));
 AOI21_X1 _41089_ (.A(_14742_),
    .B1(_13010_),
    .B2(_13013_),
    .ZN(_14749_));
 OR2_X1 _41090_ (.A1(_14748_),
    .A2(_14749_),
    .ZN(_14750_));
 MUX2_X2 _41091_ (.A(_14747_),
    .B(_14750_),
    .S(_14724_),
    .Z(\icache.data_mem_data_li [180]));
 AOI21_X1 _41092_ (.A(_14692_),
    .B1(_13051_),
    .B2(_13054_),
    .ZN(_14751_));
 AOI21_X1 _41093_ (.A(_14700_),
    .B1(_13042_),
    .B2(_13046_),
    .ZN(_14752_));
 OR2_X2 _41094_ (.A1(_14751_),
    .A2(_14752_),
    .ZN(_14753_));
 AOI21_X1 _41095_ (.A(_14734_),
    .B1(_13067_),
    .B2(_13070_),
    .ZN(_14754_));
 AOI21_X1 _41096_ (.A(_14742_),
    .B1(_13059_),
    .B2(_13063_),
    .ZN(_14755_));
 OR2_X1 _41097_ (.A1(_14754_),
    .A2(_14755_),
    .ZN(_14756_));
 MUX2_X2 _41098_ (.A(_14753_),
    .B(_14756_),
    .S(_14724_),
    .Z(\icache.data_mem_data_li [181]));
 BUF_X8 _41099_ (.A(_14159_),
    .Z(_14757_));
 AOI21_X1 _41100_ (.A(_14757_),
    .B1(_13084_),
    .B2(_13087_),
    .ZN(_14758_));
 AOI21_X1 _41101_ (.A(_14700_),
    .B1(_13075_),
    .B2(_13079_),
    .ZN(_14759_));
 OR2_X4 _41102_ (.A1(_14758_),
    .A2(_14759_),
    .ZN(_14760_));
 AOI21_X1 _41103_ (.A(_14734_),
    .B1(_13100_),
    .B2(_13103_),
    .ZN(_14761_));
 AOI21_X1 _41104_ (.A(_14742_),
    .B1(_13093_),
    .B2(_13096_),
    .ZN(_14762_));
 OR2_X4 _41105_ (.A1(_14761_),
    .A2(_14762_),
    .ZN(_14763_));
 BUF_X8 _41106_ (.A(_13481_),
    .Z(_14764_));
 MUX2_X2 _41107_ (.A(_14760_),
    .B(_14763_),
    .S(_14764_),
    .Z(\icache.data_mem_data_li [182]));
 AOI21_X1 _41108_ (.A(_14757_),
    .B1(_13115_),
    .B2(_13118_),
    .ZN(_14765_));
 BUF_X8 _41109_ (.A(_14180_),
    .Z(_14766_));
 AOI21_X1 _41110_ (.A(_14766_),
    .B1(_13108_),
    .B2(_13111_),
    .ZN(_14767_));
 OR2_X1 _41111_ (.A1(_14765_),
    .A2(_14767_),
    .ZN(_14768_));
 AOI21_X1 _41112_ (.A(_14734_),
    .B1(_13132_),
    .B2(_13135_),
    .ZN(_14769_));
 AOI21_X1 _41113_ (.A(_14742_),
    .B1(_13123_),
    .B2(_13128_),
    .ZN(_14770_));
 OR2_X1 _41114_ (.A1(_14769_),
    .A2(_14770_),
    .ZN(_14771_));
 MUX2_X2 _41115_ (.A(_14768_),
    .B(_14771_),
    .S(_14724_),
    .Z(\icache.data_mem_data_li [183]));
 AOI21_X1 _41116_ (.A(_14757_),
    .B1(_13165_),
    .B2(_13168_),
    .ZN(_14772_));
 AOI21_X1 _41117_ (.A(_14766_),
    .B1(_13158_),
    .B2(_13161_),
    .ZN(_14773_));
 OR2_X2 _41118_ (.A1(_14772_),
    .A2(_14773_),
    .ZN(_14774_));
 AOI21_X1 _41119_ (.A(_14734_),
    .B1(_13150_),
    .B2(_13153_),
    .ZN(_14775_));
 AOI21_X1 _41120_ (.A(_14742_),
    .B1(_13141_),
    .B2(_13144_),
    .ZN(_14776_));
 OR2_X2 _41121_ (.A1(_14775_),
    .A2(_14776_),
    .ZN(_14777_));
 MUX2_X2 _41122_ (.A(_14774_),
    .B(_14777_),
    .S(_14764_),
    .Z(\icache.data_mem_data_li [184]));
 AOI21_X1 _41123_ (.A(_14757_),
    .B1(_13185_),
    .B2(_13188_),
    .ZN(_14778_));
 AOI21_X1 _41124_ (.A(_14766_),
    .B1(_13175_),
    .B2(_13180_),
    .ZN(_14779_));
 OR2_X1 _41125_ (.A1(_14778_),
    .A2(_14779_),
    .ZN(_14780_));
 AOI21_X1 _41126_ (.A(_14734_),
    .B1(_13200_),
    .B2(_13203_),
    .ZN(_14781_));
 AOI21_X1 _41127_ (.A(_14742_),
    .B1(_13193_),
    .B2(_13196_),
    .ZN(_14782_));
 OR2_X1 _41128_ (.A1(_14781_),
    .A2(_14782_),
    .ZN(_14783_));
 MUX2_X2 _41129_ (.A(_14780_),
    .B(_14783_),
    .S(_14724_),
    .Z(\icache.data_mem_data_li [185]));
 AOI21_X1 _41130_ (.A(_14757_),
    .B1(_13215_),
    .B2(_13219_),
    .ZN(_14784_));
 AOI21_X1 _41131_ (.A(_14766_),
    .B1(_13208_),
    .B2(_13211_),
    .ZN(_14785_));
 OR2_X1 _41132_ (.A1(_14784_),
    .A2(_14785_),
    .ZN(_14786_));
 AOI21_X1 _41133_ (.A(_14734_),
    .B1(_13232_),
    .B2(_13235_),
    .ZN(_14787_));
 AOI21_X1 _41134_ (.A(_14742_),
    .B1(_13225_),
    .B2(_13228_),
    .ZN(_14788_));
 OR2_X1 _41135_ (.A1(_14787_),
    .A2(_14788_),
    .ZN(_14789_));
 MUX2_X2 _41136_ (.A(_14786_),
    .B(_14789_),
    .S(_14724_),
    .Z(\icache.data_mem_data_li [186]));
 AOI21_X1 _41137_ (.A(_14757_),
    .B1(_13247_),
    .B2(_13251_),
    .ZN(_14790_));
 AOI21_X1 _41138_ (.A(_14766_),
    .B1(_13240_),
    .B2(_13243_),
    .ZN(_14791_));
 OR2_X1 _41139_ (.A1(_14790_),
    .A2(_14791_),
    .ZN(_14792_));
 AOI21_X1 _41140_ (.A(_14734_),
    .B1(_13266_),
    .B2(_13269_),
    .ZN(_14793_));
 AOI21_X1 _41141_ (.A(_14742_),
    .B1(_13257_),
    .B2(_13261_),
    .ZN(_14794_));
 OR2_X1 _41142_ (.A1(_14793_),
    .A2(_14794_),
    .ZN(_14795_));
 MUX2_X2 _41143_ (.A(_14792_),
    .B(_14795_),
    .S(_14724_),
    .Z(\icache.data_mem_data_li [187]));
 AOI21_X1 _41144_ (.A(_14757_),
    .B1(_13281_),
    .B2(_13284_),
    .ZN(_14796_));
 AOI21_X1 _41145_ (.A(_14766_),
    .B1(_13274_),
    .B2(_13277_),
    .ZN(_14797_));
 OR2_X1 _41146_ (.A1(_14796_),
    .A2(_14797_),
    .ZN(_14798_));
 BUF_X8 _41147_ (.A(_11239_),
    .Z(_14799_));
 AOI21_X1 _41148_ (.A(_14799_),
    .B1(_13299_),
    .B2(_13302_),
    .ZN(_14800_));
 AOI21_X1 _41149_ (.A(_14742_),
    .B1(_13289_),
    .B2(_13294_),
    .ZN(_14801_));
 OR2_X1 _41150_ (.A1(_14800_),
    .A2(_14801_),
    .ZN(_14802_));
 MUX2_X2 _41151_ (.A(_14798_),
    .B(_14802_),
    .S(_14724_),
    .Z(\icache.data_mem_data_li [188]));
 AOI21_X1 _41152_ (.A(_14757_),
    .B1(_13330_),
    .B2(_13333_),
    .ZN(_14803_));
 AOI21_X1 _41153_ (.A(_14766_),
    .B1(_13323_),
    .B2(_13326_),
    .ZN(_14804_));
 OR2_X1 _41154_ (.A1(_14803_),
    .A2(_14804_),
    .ZN(_14805_));
 AOI21_X1 _41155_ (.A(_14799_),
    .B1(_13315_),
    .B2(_13318_),
    .ZN(_14806_));
 BUF_X8 _41156_ (.A(_11257_),
    .Z(_14807_));
 AOI21_X1 _41157_ (.A(_14807_),
    .B1(_13307_),
    .B2(_13310_),
    .ZN(_14808_));
 OR2_X1 _41158_ (.A1(_14806_),
    .A2(_14808_),
    .ZN(_14809_));
 MUX2_X2 _41159_ (.A(_14805_),
    .B(_14809_),
    .S(_14764_),
    .Z(\icache.data_mem_data_li [189]));
 AOI21_X1 _41160_ (.A(_14757_),
    .B1(_13350_),
    .B2(_13353_),
    .ZN(_14810_));
 AOI21_X1 _41161_ (.A(_14766_),
    .B1(_13339_),
    .B2(_13346_),
    .ZN(_14811_));
 OR2_X2 _41162_ (.A1(_14810_),
    .A2(_14811_),
    .ZN(_14812_));
 AOI21_X1 _41163_ (.A(_14799_),
    .B1(_13365_),
    .B2(_13368_),
    .ZN(_14813_));
 AOI21_X1 _41164_ (.A(_14807_),
    .B1(_13358_),
    .B2(_13361_),
    .ZN(_14814_));
 OR2_X2 _41165_ (.A1(_14813_),
    .A2(_14814_),
    .ZN(_14815_));
 BUF_X32 _41166_ (.A(_08431_),
    .Z(_14816_));
 BUF_X4 _41167_ (.A(_14816_),
    .Z(_14817_));
 MUX2_X2 _41168_ (.A(_14812_),
    .B(_14815_),
    .S(_14817_),
    .Z(\icache.data_mem_data_li [190]));
 AOI21_X1 _41169_ (.A(_14757_),
    .B1(_13381_),
    .B2(_13384_),
    .ZN(_14818_));
 AOI21_X1 _41170_ (.A(_14766_),
    .B1(_13373_),
    .B2(_13376_),
    .ZN(_14819_));
 OR2_X2 _41171_ (.A1(_14818_),
    .A2(_14819_),
    .ZN(_14820_));
 AOI21_X1 _41172_ (.A(_14799_),
    .B1(_13396_),
    .B2(_13399_),
    .ZN(_14821_));
 AOI21_X1 _41173_ (.A(_14807_),
    .B1(_13389_),
    .B2(_13392_),
    .ZN(_14822_));
 OR2_X2 _41174_ (.A1(_14821_),
    .A2(_14822_),
    .ZN(_14823_));
 MUX2_X2 _41175_ (.A(_14820_),
    .B(_14823_),
    .S(_14764_),
    .Z(\icache.data_mem_data_li [191]));
 BUF_X8 _41176_ (.A(_14159_),
    .Z(_14824_));
 AOI21_X2 _41177_ (.A(_14824_),
    .B1(_13405_),
    .B2(_13406_),
    .ZN(_14825_));
 AOI21_X1 _41178_ (.A(_14766_),
    .B1(_13402_),
    .B2(_13403_),
    .ZN(_14826_));
 OR2_X2 _41179_ (.A1(_14825_),
    .A2(_14826_),
    .ZN(_14827_));
 AOI21_X1 _41180_ (.A(_14799_),
    .B1(_13413_),
    .B2(_13414_),
    .ZN(_14828_));
 AOI21_X1 _41181_ (.A(_14807_),
    .B1(_13410_),
    .B2(_13411_),
    .ZN(_14829_));
 OR2_X4 _41182_ (.A1(_14828_),
    .A2(_14829_),
    .ZN(_14830_));
 MUX2_X2 _41183_ (.A(_14827_),
    .B(_14830_),
    .S(_14817_),
    .Z(\icache.data_mem_data_li [192]));
 AOI21_X1 _41184_ (.A(_14824_),
    .B1(_13429_),
    .B2(_13430_),
    .ZN(_14831_));
 BUF_X8 _41185_ (.A(_14180_),
    .Z(_14832_));
 AOI21_X2 _41186_ (.A(_14832_),
    .B1(_13426_),
    .B2(_13427_),
    .ZN(_14833_));
 OR2_X4 _41187_ (.A1(_14831_),
    .A2(_14833_),
    .ZN(_14834_));
 AOI21_X1 _41188_ (.A(_14799_),
    .B1(_13422_),
    .B2(_13423_),
    .ZN(_14835_));
 AOI21_X1 _41189_ (.A(_14807_),
    .B1(_13417_),
    .B2(_13420_),
    .ZN(_14836_));
 OR2_X4 _41190_ (.A1(_14835_),
    .A2(_14836_),
    .ZN(_14837_));
 MUX2_X2 _41191_ (.A(_14834_),
    .B(_14837_),
    .S(_14764_),
    .Z(\icache.data_mem_data_li [193]));
 AOI21_X1 _41192_ (.A(_14824_),
    .B1(_13437_),
    .B2(_13438_),
    .ZN(_14838_));
 AOI21_X1 _41193_ (.A(_14832_),
    .B1(_13434_),
    .B2(_13435_),
    .ZN(_14839_));
 OR2_X4 _41194_ (.A1(_14838_),
    .A2(_14839_),
    .ZN(_14840_));
 AOI21_X1 _41195_ (.A(_14799_),
    .B1(_13444_),
    .B2(_13445_),
    .ZN(_14841_));
 AOI21_X2 _41196_ (.A(_14807_),
    .B1(_13441_),
    .B2(_13442_),
    .ZN(_14842_));
 OR2_X4 _41197_ (.A1(_14841_),
    .A2(_14842_),
    .ZN(_14843_));
 MUX2_X2 _41198_ (.A(_14840_),
    .B(_14843_),
    .S(_14817_),
    .Z(\icache.data_mem_data_li [194]));
 AOI21_X1 _41199_ (.A(_14824_),
    .B1(_13453_),
    .B2(_13454_),
    .ZN(_14844_));
 AOI21_X1 _41200_ (.A(_14832_),
    .B1(_13448_),
    .B2(_13451_),
    .ZN(_14845_));
 OR2_X4 _41201_ (.A1(_14844_),
    .A2(_14845_),
    .ZN(_14846_));
 AOI21_X1 _41202_ (.A(_14799_),
    .B1(_13460_),
    .B2(_13461_),
    .ZN(_14847_));
 AOI21_X2 _41203_ (.A(_14807_),
    .B1(_13457_),
    .B2(_13458_),
    .ZN(_14848_));
 OR2_X4 _41204_ (.A1(_14847_),
    .A2(_14848_),
    .ZN(_14849_));
 MUX2_X2 _41205_ (.A(_14846_),
    .B(_14849_),
    .S(_14817_),
    .Z(\icache.data_mem_data_li [195]));
 AOI21_X1 _41206_ (.A(_14824_),
    .B1(_13477_),
    .B2(_13478_),
    .ZN(_14850_));
 AOI21_X2 _41207_ (.A(_14832_),
    .B1(_13474_),
    .B2(_13475_),
    .ZN(_14851_));
 OR2_X4 _41208_ (.A1(_14850_),
    .A2(_14851_),
    .ZN(_14852_));
 AOI21_X1 _41209_ (.A(_14799_),
    .B1(_13468_),
    .B2(_13469_),
    .ZN(_14853_));
 AOI21_X1 _41210_ (.A(_14807_),
    .B1(_13465_),
    .B2(_13466_),
    .ZN(_14854_));
 OR2_X4 _41211_ (.A1(_14853_),
    .A2(_14854_),
    .ZN(_14855_));
 MUX2_X2 _41212_ (.A(_14852_),
    .B(_14855_),
    .S(_14817_),
    .Z(\icache.data_mem_data_li [196]));
 AOI21_X1 _41213_ (.A(_14824_),
    .B1(_13496_),
    .B2(_13497_),
    .ZN(_14856_));
 AOI21_X1 _41214_ (.A(_14832_),
    .B1(_13491_),
    .B2(_13492_),
    .ZN(_14857_));
 OR2_X4 _41215_ (.A1(_14856_),
    .A2(_14857_),
    .ZN(_14858_));
 AOI21_X1 _41216_ (.A(_14799_),
    .B1(_13487_),
    .B2(_13488_),
    .ZN(_14859_));
 AOI21_X1 _41217_ (.A(_14807_),
    .B1(_13484_),
    .B2(_13485_),
    .ZN(_14860_));
 OR2_X4 _41218_ (.A1(_14859_),
    .A2(_14860_),
    .ZN(_14861_));
 MUX2_X2 _41219_ (.A(_14858_),
    .B(_14861_),
    .S(_14764_),
    .Z(\icache.data_mem_data_li [197]));
 AOI21_X1 _41220_ (.A(_14824_),
    .B1(_13512_),
    .B2(_13513_),
    .ZN(_14862_));
 AOI21_X1 _41221_ (.A(_14832_),
    .B1(_13509_),
    .B2(_13510_),
    .ZN(_14863_));
 OR2_X4 _41222_ (.A1(_14862_),
    .A2(_14863_),
    .ZN(_14864_));
 BUF_X8 _41223_ (.A(_11239_),
    .Z(_14865_));
 AOI21_X1 _41224_ (.A(_14865_),
    .B1(_13505_),
    .B2(_13506_),
    .ZN(_14866_));
 AOI21_X1 _41225_ (.A(_14807_),
    .B1(_13500_),
    .B2(_13503_),
    .ZN(_14867_));
 OR2_X4 _41226_ (.A1(_14866_),
    .A2(_14867_),
    .ZN(_14868_));
 MUX2_X2 _41227_ (.A(_14864_),
    .B(_14868_),
    .S(_14764_),
    .Z(\icache.data_mem_data_li [198]));
 AOI21_X1 _41228_ (.A(_14824_),
    .B1(_13520_),
    .B2(_13521_),
    .ZN(_14869_));
 AOI21_X1 _41229_ (.A(_14832_),
    .B1(_13517_),
    .B2(_13518_),
    .ZN(_14870_));
 OR2_X4 _41230_ (.A1(_14869_),
    .A2(_14870_),
    .ZN(_14871_));
 AOI21_X1 _41231_ (.A(_14865_),
    .B1(_13527_),
    .B2(_13528_),
    .ZN(_14872_));
 BUF_X8 _41232_ (.A(_11257_),
    .Z(_14873_));
 AOI21_X1 _41233_ (.A(_14873_),
    .B1(_13524_),
    .B2(_13525_),
    .ZN(_14874_));
 OR2_X4 _41234_ (.A1(_14872_),
    .A2(_14874_),
    .ZN(_14875_));
 MUX2_X2 _41235_ (.A(_14871_),
    .B(_14875_),
    .S(_14817_),
    .Z(\icache.data_mem_data_li [199]));
 AOI21_X1 _41236_ (.A(_14824_),
    .B1(_13537_),
    .B2(_13538_),
    .ZN(_14876_));
 AOI21_X1 _41237_ (.A(_14832_),
    .B1(_13532_),
    .B2(_13535_),
    .ZN(_14877_));
 OR2_X4 _41238_ (.A1(_14876_),
    .A2(_14877_),
    .ZN(_14878_));
 AOI21_X1 _41239_ (.A(_14865_),
    .B1(_13544_),
    .B2(_13545_),
    .ZN(_14879_));
 AOI21_X1 _41240_ (.A(_14873_),
    .B1(_13541_),
    .B2(_13542_),
    .ZN(_14880_));
 OR2_X4 _41241_ (.A1(_14879_),
    .A2(_14880_),
    .ZN(_14881_));
 MUX2_X2 _41242_ (.A(_14878_),
    .B(_14881_),
    .S(_14764_),
    .Z(\icache.data_mem_data_li [200]));
 AOI21_X1 _41243_ (.A(_14824_),
    .B1(_13552_),
    .B2(_13553_),
    .ZN(_14882_));
 AOI21_X1 _41244_ (.A(_14832_),
    .B1(_13548_),
    .B2(_13549_),
    .ZN(_14883_));
 OR2_X4 _41245_ (.A1(_14882_),
    .A2(_14883_),
    .ZN(_14884_));
 AOI21_X1 _41246_ (.A(_14865_),
    .B1(_13559_),
    .B2(_13560_),
    .ZN(_14885_));
 AOI21_X1 _41247_ (.A(_14873_),
    .B1(_13556_),
    .B2(_13557_),
    .ZN(_14886_));
 OR2_X4 _41248_ (.A1(_14885_),
    .A2(_14886_),
    .ZN(_14887_));
 MUX2_X2 _41249_ (.A(_14884_),
    .B(_14887_),
    .S(_14817_),
    .Z(\icache.data_mem_data_li [201]));
 BUF_X8 _41250_ (.A(_14159_),
    .Z(_14888_));
 AOI21_X2 _41251_ (.A(_14888_),
    .B1(_13566_),
    .B2(_13567_),
    .ZN(_14889_));
 AOI21_X1 _41252_ (.A(_14832_),
    .B1(_13563_),
    .B2(_13564_),
    .ZN(_14890_));
 OR2_X4 _41253_ (.A1(_14889_),
    .A2(_14890_),
    .ZN(_14891_));
 AOI21_X1 _41254_ (.A(_14865_),
    .B1(_13574_),
    .B2(_13575_),
    .ZN(_14892_));
 AOI21_X1 _41255_ (.A(_14873_),
    .B1(_13571_),
    .B2(_13572_),
    .ZN(_14893_));
 OR2_X4 _41256_ (.A1(_14892_),
    .A2(_14893_),
    .ZN(_14894_));
 MUX2_X2 _41257_ (.A(_14891_),
    .B(_14894_),
    .S(_14817_),
    .Z(\icache.data_mem_data_li [202]));
 AOI21_X1 _41258_ (.A(_14888_),
    .B1(_13581_),
    .B2(_13582_),
    .ZN(_14895_));
 BUF_X8 _41259_ (.A(_14180_),
    .Z(_14896_));
 AOI21_X1 _41260_ (.A(_14896_),
    .B1(_13578_),
    .B2(_13579_),
    .ZN(_14897_));
 OR2_X4 _41261_ (.A1(_14895_),
    .A2(_14897_),
    .ZN(_14898_));
 AOI21_X1 _41262_ (.A(_14865_),
    .B1(_13590_),
    .B2(_13591_),
    .ZN(_14899_));
 AOI21_X1 _41263_ (.A(_14873_),
    .B1(_13585_),
    .B2(_13588_),
    .ZN(_14900_));
 OR2_X4 _41264_ (.A1(_14899_),
    .A2(_14900_),
    .ZN(_14901_));
 MUX2_X2 _41265_ (.A(_14898_),
    .B(_14901_),
    .S(_14817_),
    .Z(\icache.data_mem_data_li [203]));
 AOI21_X1 _41266_ (.A(_14888_),
    .B1(_13605_),
    .B2(_13606_),
    .ZN(_14902_));
 AOI21_X1 _41267_ (.A(_14896_),
    .B1(_13602_),
    .B2(_13603_),
    .ZN(_14903_));
 OR2_X4 _41268_ (.A1(_14902_),
    .A2(_14903_),
    .ZN(_14904_));
 AOI21_X1 _41269_ (.A(_14865_),
    .B1(_13598_),
    .B2(_13599_),
    .ZN(_14905_));
 AOI21_X1 _41270_ (.A(_14873_),
    .B1(_13594_),
    .B2(_13595_),
    .ZN(_14906_));
 OR2_X4 _41271_ (.A1(_14905_),
    .A2(_14906_),
    .ZN(_14907_));
 MUX2_X2 _41272_ (.A(_14904_),
    .B(_14907_),
    .S(_14764_),
    .Z(\icache.data_mem_data_li [204]));
 AOI21_X1 _41273_ (.A(_14888_),
    .B1(_13621_),
    .B2(_13622_),
    .ZN(_14908_));
 AOI21_X1 _41274_ (.A(_14896_),
    .B1(_13618_),
    .B2(_13619_),
    .ZN(_14909_));
 OR2_X4 _41275_ (.A1(_14908_),
    .A2(_14909_),
    .ZN(_14910_));
 AOI21_X1 _41276_ (.A(_14865_),
    .B1(_13612_),
    .B2(_13615_),
    .ZN(_14911_));
 AOI21_X1 _41277_ (.A(_14873_),
    .B1(_13609_),
    .B2(_13610_),
    .ZN(_14912_));
 OR2_X4 _41278_ (.A1(_14911_),
    .A2(_14912_),
    .ZN(_14913_));
 MUX2_X2 _41279_ (.A(_14910_),
    .B(_14913_),
    .S(_14764_),
    .Z(\icache.data_mem_data_li [205]));
 AOI21_X1 _41280_ (.A(_14888_),
    .B1(_13636_),
    .B2(_13637_),
    .ZN(_14914_));
 AOI21_X1 _41281_ (.A(_14896_),
    .B1(_13633_),
    .B2(_13634_),
    .ZN(_14915_));
 OR2_X4 _41282_ (.A1(_14914_),
    .A2(_14915_),
    .ZN(_14916_));
 AOI21_X1 _41283_ (.A(_14865_),
    .B1(_13628_),
    .B2(_13629_),
    .ZN(_14917_));
 AOI21_X1 _41284_ (.A(_14873_),
    .B1(_13625_),
    .B2(_13626_),
    .ZN(_14918_));
 OR2_X4 _41285_ (.A1(_14917_),
    .A2(_14918_),
    .ZN(_14919_));
 MUX2_X2 _41286_ (.A(_14916_),
    .B(_14919_),
    .S(_14817_),
    .Z(\icache.data_mem_data_li [206]));
 AOI21_X1 _41287_ (.A(_14888_),
    .B1(_13643_),
    .B2(_13644_),
    .ZN(_14920_));
 AOI21_X1 _41288_ (.A(_14896_),
    .B1(_13640_),
    .B2(_13641_),
    .ZN(_14921_));
 OR2_X4 _41289_ (.A1(_14920_),
    .A2(_14921_),
    .ZN(_14922_));
 AOI21_X1 _41290_ (.A(_14865_),
    .B1(_13652_),
    .B2(_13653_),
    .ZN(_14923_));
 AOI21_X1 _41291_ (.A(_14873_),
    .B1(_13648_),
    .B2(_13649_),
    .ZN(_14924_));
 OR2_X4 _41292_ (.A1(_14923_),
    .A2(_14924_),
    .ZN(_14925_));
 BUF_X8 _41293_ (.A(_13481_),
    .Z(_14926_));
 MUX2_X2 _41294_ (.A(_14922_),
    .B(_14925_),
    .S(_14926_),
    .Z(\icache.data_mem_data_li [207]));
 AOI21_X1 _41295_ (.A(_14888_),
    .B1(_13668_),
    .B2(_13669_),
    .ZN(_14927_));
 AOI21_X1 _41296_ (.A(_14896_),
    .B1(_13665_),
    .B2(_13666_),
    .ZN(_14928_));
 OR2_X4 _41297_ (.A1(_14927_),
    .A2(_14928_),
    .ZN(_14929_));
 BUF_X8 _41298_ (.A(_11239_),
    .Z(_14930_));
 AOI21_X1 _41299_ (.A(_14930_),
    .B1(_13661_),
    .B2(_13662_),
    .ZN(_14931_));
 AOI21_X1 _41300_ (.A(_14873_),
    .B1(_13656_),
    .B2(_13659_),
    .ZN(_14932_));
 OR2_X4 _41301_ (.A1(_14931_),
    .A2(_14932_),
    .ZN(_14933_));
 BUF_X4 _41302_ (.A(_14816_),
    .Z(_14934_));
 MUX2_X2 _41303_ (.A(_14929_),
    .B(_14933_),
    .S(_14934_),
    .Z(\icache.data_mem_data_li [208]));
 AOI21_X1 _41304_ (.A(_14888_),
    .B1(_13683_),
    .B2(_13684_),
    .ZN(_14935_));
 AOI21_X1 _41305_ (.A(_14896_),
    .B1(_13680_),
    .B2(_13681_),
    .ZN(_14936_));
 OR2_X4 _41306_ (.A1(_14935_),
    .A2(_14936_),
    .ZN(_14937_));
 AOI21_X1 _41307_ (.A(_14930_),
    .B1(_13676_),
    .B2(_13677_),
    .ZN(_14938_));
 BUF_X8 _41308_ (.A(_11257_),
    .Z(_14939_));
 AOI21_X1 _41309_ (.A(_14939_),
    .B1(_13672_),
    .B2(_13673_),
    .ZN(_14940_));
 OR2_X4 _41310_ (.A1(_14938_),
    .A2(_14940_),
    .ZN(_14941_));
 MUX2_X2 _41311_ (.A(_14937_),
    .B(_14941_),
    .S(_14926_),
    .Z(\icache.data_mem_data_li [209]));
 AOI21_X1 _41312_ (.A(_14888_),
    .B1(_13693_),
    .B2(_13694_),
    .ZN(_14942_));
 AOI21_X1 _41313_ (.A(_14896_),
    .B1(_13688_),
    .B2(_13691_),
    .ZN(_14943_));
 OR2_X4 _41314_ (.A1(_14942_),
    .A2(_14943_),
    .ZN(_14944_));
 AOI21_X1 _41315_ (.A(_14930_),
    .B1(_13700_),
    .B2(_13701_),
    .ZN(_14945_));
 AOI21_X1 _41316_ (.A(_14939_),
    .B1(_13697_),
    .B2(_13698_),
    .ZN(_14946_));
 OR2_X4 _41317_ (.A1(_14945_),
    .A2(_14946_),
    .ZN(_14947_));
 MUX2_X2 _41318_ (.A(_14944_),
    .B(_14947_),
    .S(_14934_),
    .Z(\icache.data_mem_data_li [210]));
 AOI21_X1 _41319_ (.A(_14888_),
    .B1(_13709_),
    .B2(_13710_),
    .ZN(_14948_));
 AOI21_X1 _41320_ (.A(_14896_),
    .B1(_13705_),
    .B2(_13706_),
    .ZN(_14949_));
 OR2_X4 _41321_ (.A1(_14948_),
    .A2(_14949_),
    .ZN(_14950_));
 AOI21_X1 _41322_ (.A(_14930_),
    .B1(_13716_),
    .B2(_13717_),
    .ZN(_14951_));
 AOI21_X1 _41323_ (.A(_14939_),
    .B1(_13713_),
    .B2(_13714_),
    .ZN(_14952_));
 OR2_X4 _41324_ (.A1(_14951_),
    .A2(_14952_),
    .ZN(_14953_));
 MUX2_X2 _41325_ (.A(_14950_),
    .B(_14953_),
    .S(_14934_),
    .Z(\icache.data_mem_data_li [211]));
 BUF_X8 _41326_ (.A(_08447_),
    .Z(_14954_));
 AOI21_X1 _41327_ (.A(_14954_),
    .B1(_13731_),
    .B2(_13732_),
    .ZN(_14955_));
 AOI21_X2 _41328_ (.A(_14896_),
    .B1(_13728_),
    .B2(_13729_),
    .ZN(_14956_));
 OR2_X4 _41329_ (.A1(_14955_),
    .A2(_14956_),
    .ZN(_14957_));
 AOI21_X1 _41330_ (.A(_14930_),
    .B1(_13724_),
    .B2(_13725_),
    .ZN(_14958_));
 AOI21_X1 _41331_ (.A(_14939_),
    .B1(_13721_),
    .B2(_13722_),
    .ZN(_14959_));
 OR2_X4 _41332_ (.A1(_14958_),
    .A2(_14959_),
    .ZN(_14960_));
 MUX2_X2 _41333_ (.A(_14957_),
    .B(_14960_),
    .S(_14934_),
    .Z(\icache.data_mem_data_li [212]));
 AOI21_X1 _41334_ (.A(_14954_),
    .B1(_13738_),
    .B2(_13739_),
    .ZN(_14961_));
 BUF_X8 _41335_ (.A(_08446_),
    .Z(_14962_));
 AOI21_X1 _41336_ (.A(_14962_),
    .B1(_13735_),
    .B2(_13736_),
    .ZN(_14963_));
 OR2_X4 _41337_ (.A1(_14961_),
    .A2(_14963_),
    .ZN(_14964_));
 AOI21_X1 _41338_ (.A(_14930_),
    .B1(_13747_),
    .B2(_13748_),
    .ZN(_14965_));
 AOI21_X1 _41339_ (.A(_14939_),
    .B1(_13742_),
    .B2(_13745_),
    .ZN(_14966_));
 OR2_X4 _41340_ (.A1(_14965_),
    .A2(_14966_),
    .ZN(_14967_));
 MUX2_X2 _41341_ (.A(_14964_),
    .B(_14967_),
    .S(_14934_),
    .Z(\icache.data_mem_data_li [213]));
 AOI21_X1 _41342_ (.A(_14954_),
    .B1(_13762_),
    .B2(_13763_),
    .ZN(_14968_));
 AOI21_X1 _41343_ (.A(_14962_),
    .B1(_13759_),
    .B2(_13760_),
    .ZN(_14969_));
 OR2_X4 _41344_ (.A1(_14968_),
    .A2(_14969_),
    .ZN(_14970_));
 AOI21_X1 _41345_ (.A(_14930_),
    .B1(_13755_),
    .B2(_13756_),
    .ZN(_14971_));
 AOI21_X1 _41346_ (.A(_14939_),
    .B1(_13751_),
    .B2(_13752_),
    .ZN(_14972_));
 OR2_X4 _41347_ (.A1(_14971_),
    .A2(_14972_),
    .ZN(_14973_));
 MUX2_X2 _41348_ (.A(_14970_),
    .B(_14973_),
    .S(_14926_),
    .Z(\icache.data_mem_data_li [214]));
 AOI21_X1 _41349_ (.A(_14954_),
    .B1(_13771_),
    .B2(_13772_),
    .ZN(_14974_));
 AOI21_X1 _41350_ (.A(_14962_),
    .B1(_13766_),
    .B2(_13769_),
    .ZN(_14975_));
 OR2_X4 _41351_ (.A1(_14974_),
    .A2(_14975_),
    .ZN(_14976_));
 AOI21_X1 _41352_ (.A(_14930_),
    .B1(_13778_),
    .B2(_13779_),
    .ZN(_14977_));
 AOI21_X1 _41353_ (.A(_14939_),
    .B1(_13775_),
    .B2(_13776_),
    .ZN(_14978_));
 OR2_X4 _41354_ (.A1(_14977_),
    .A2(_14978_),
    .ZN(_14979_));
 MUX2_X2 _41355_ (.A(_14976_),
    .B(_14979_),
    .S(_14934_),
    .Z(\icache.data_mem_data_li [215]));
 AOI21_X1 _41356_ (.A(_14954_),
    .B1(_13793_),
    .B2(_13794_),
    .ZN(_14980_));
 AOI21_X1 _41357_ (.A(_14962_),
    .B1(_13790_),
    .B2(_13791_),
    .ZN(_14981_));
 OR2_X4 _41358_ (.A1(_14980_),
    .A2(_14981_),
    .ZN(_14982_));
 AOI21_X1 _41359_ (.A(_14930_),
    .B1(_13785_),
    .B2(_13786_),
    .ZN(_14983_));
 AOI21_X1 _41360_ (.A(_14939_),
    .B1(_13782_),
    .B2(_13783_),
    .ZN(_14984_));
 OR2_X4 _41361_ (.A1(_14983_),
    .A2(_14984_),
    .ZN(_14985_));
 MUX2_X2 _41362_ (.A(_14982_),
    .B(_14985_),
    .S(_14926_),
    .Z(\icache.data_mem_data_li [216]));
 AOI21_X1 _41363_ (.A(_14954_),
    .B1(_13809_),
    .B2(_13810_),
    .ZN(_14986_));
 AOI21_X1 _41364_ (.A(_14962_),
    .B1(_13805_),
    .B2(_13806_),
    .ZN(_14987_));
 OR2_X4 _41365_ (.A1(_14986_),
    .A2(_14987_),
    .ZN(_14988_));
 AOI21_X1 _41366_ (.A(_14930_),
    .B1(_13801_),
    .B2(_13802_),
    .ZN(_14989_));
 AOI21_X1 _41367_ (.A(_14939_),
    .B1(_13798_),
    .B2(_13799_),
    .ZN(_14990_));
 OR2_X4 _41368_ (.A1(_14989_),
    .A2(_14990_),
    .ZN(_14991_));
 MUX2_X2 _41369_ (.A(_14988_),
    .B(_14991_),
    .S(_14934_),
    .Z(\icache.data_mem_data_li [217]));
 AOI21_X1 _41370_ (.A(_14954_),
    .B1(_13825_),
    .B2(_13826_),
    .ZN(_14992_));
 AOI21_X1 _41371_ (.A(_14962_),
    .B1(_13822_),
    .B2(_13823_),
    .ZN(_14993_));
 OR2_X4 _41372_ (.A1(_14992_),
    .A2(_14993_),
    .ZN(_14994_));
 BUF_X8 _41373_ (.A(_11239_),
    .Z(_14995_));
 AOI21_X1 _41374_ (.A(_14995_),
    .B1(_13818_),
    .B2(_13819_),
    .ZN(_14996_));
 AOI21_X1 _41375_ (.A(_14939_),
    .B1(_13813_),
    .B2(_13816_),
    .ZN(_14997_));
 OR2_X2 _41376_ (.A1(_14996_),
    .A2(_14997_),
    .ZN(_14998_));
 MUX2_X2 _41377_ (.A(_14994_),
    .B(_14998_),
    .S(_14934_),
    .Z(\icache.data_mem_data_li [218]));
 AOI21_X1 _41378_ (.A(_14954_),
    .B1(_13833_),
    .B2(_13834_),
    .ZN(_14999_));
 AOI21_X1 _41379_ (.A(_14962_),
    .B1(_13830_),
    .B2(_13831_),
    .ZN(_15000_));
 OR2_X4 _41380_ (.A1(_14999_),
    .A2(_15000_),
    .ZN(_15001_));
 AOI21_X1 _41381_ (.A(_14995_),
    .B1(_13840_),
    .B2(_13841_),
    .ZN(_15002_));
 BUF_X8 _41382_ (.A(_11257_),
    .Z(_15003_));
 AOI21_X1 _41383_ (.A(_15003_),
    .B1(_13837_),
    .B2(_13838_),
    .ZN(_15004_));
 OR2_X1 _41384_ (.A1(_15002_),
    .A2(_15004_),
    .ZN(_15005_));
 MUX2_X2 _41385_ (.A(_15001_),
    .B(_15005_),
    .S(_14934_),
    .Z(\icache.data_mem_data_li [219]));
 AOI21_X1 _41386_ (.A(_14954_),
    .B1(_13850_),
    .B2(_13851_),
    .ZN(_15006_));
 AOI21_X1 _41387_ (.A(_14962_),
    .B1(_13845_),
    .B2(_13848_),
    .ZN(_15007_));
 OR2_X2 _41388_ (.A1(_15006_),
    .A2(_15007_),
    .ZN(_15008_));
 AOI21_X1 _41389_ (.A(_14995_),
    .B1(_13857_),
    .B2(_13858_),
    .ZN(_15009_));
 AOI21_X1 _41390_ (.A(_15003_),
    .B1(_13854_),
    .B2(_13855_),
    .ZN(_15010_));
 OR2_X1 _41391_ (.A1(_15009_),
    .A2(_15010_),
    .ZN(_15011_));
 MUX2_X2 _41392_ (.A(_15008_),
    .B(_15011_),
    .S(_14934_),
    .Z(\icache.data_mem_data_li [220]));
 AOI21_X1 _41393_ (.A(_14954_),
    .B1(_13872_),
    .B2(_13873_),
    .ZN(_15012_));
 AOI21_X1 _41394_ (.A(_14962_),
    .B1(_13869_),
    .B2(_13870_),
    .ZN(_15013_));
 OR2_X1 _41395_ (.A1(_15012_),
    .A2(_15013_),
    .ZN(_15014_));
 AOI21_X1 _41396_ (.A(_14995_),
    .B1(_13865_),
    .B2(_13866_),
    .ZN(_15015_));
 AOI21_X1 _41397_ (.A(_15003_),
    .B1(_13861_),
    .B2(_13862_),
    .ZN(_15016_));
 OR2_X1 _41398_ (.A1(_15015_),
    .A2(_15016_),
    .ZN(_15017_));
 MUX2_X2 _41399_ (.A(_15014_),
    .B(_15017_),
    .S(_14926_),
    .Z(\icache.data_mem_data_li [221]));
 BUF_X8 _41400_ (.A(_08447_),
    .Z(_15018_));
 AOI21_X1 _41401_ (.A(_15018_),
    .B1(_13879_),
    .B2(_13880_),
    .ZN(_15019_));
 AOI21_X1 _41402_ (.A(_14962_),
    .B1(_13876_),
    .B2(_13877_),
    .ZN(_15020_));
 OR2_X2 _41403_ (.A1(_15019_),
    .A2(_15020_),
    .ZN(_15021_));
 AOI21_X1 _41404_ (.A(_14995_),
    .B1(_13887_),
    .B2(_13888_),
    .ZN(_15022_));
 AOI21_X1 _41405_ (.A(_15003_),
    .B1(_13884_),
    .B2(_13885_),
    .ZN(_15023_));
 OR2_X1 _41406_ (.A1(_15022_),
    .A2(_15023_),
    .ZN(_15024_));
 BUF_X4 _41407_ (.A(_14816_),
    .Z(_15025_));
 MUX2_X2 _41408_ (.A(_15021_),
    .B(_15024_),
    .S(_15025_),
    .Z(\icache.data_mem_data_li [222]));
 AOI21_X1 _41409_ (.A(_15018_),
    .B1(_13894_),
    .B2(_13895_),
    .ZN(_15026_));
 BUF_X8 _41410_ (.A(_08446_),
    .Z(_15027_));
 AOI21_X1 _41411_ (.A(_15027_),
    .B1(_13891_),
    .B2(_13892_),
    .ZN(_15028_));
 OR2_X1 _41412_ (.A1(_15026_),
    .A2(_15028_),
    .ZN(_15029_));
 AOI21_X1 _41413_ (.A(_14995_),
    .B1(_13903_),
    .B2(_13904_),
    .ZN(_15030_));
 AOI21_X1 _41414_ (.A(_15003_),
    .B1(_13898_),
    .B2(_13901_),
    .ZN(_15031_));
 OR2_X1 _41415_ (.A1(_15030_),
    .A2(_15031_),
    .ZN(_15032_));
 MUX2_X2 _41416_ (.A(_15029_),
    .B(_15032_),
    .S(_14926_),
    .Z(\icache.data_mem_data_li [223]));
 AOI21_X1 _41417_ (.A(_15018_),
    .B1(_13911_),
    .B2(_13912_),
    .ZN(_15033_));
 AOI21_X1 _41418_ (.A(_15027_),
    .B1(_13908_),
    .B2(_13909_),
    .ZN(_15034_));
 OR2_X1 _41419_ (.A1(_15033_),
    .A2(_15034_),
    .ZN(_15035_));
 AOI21_X1 _41420_ (.A(_14995_),
    .B1(_13918_),
    .B2(_13919_),
    .ZN(_15036_));
 AOI21_X1 _41421_ (.A(_15003_),
    .B1(_13915_),
    .B2(_13916_),
    .ZN(_15037_));
 OR2_X1 _41422_ (.A1(_15036_),
    .A2(_15037_),
    .ZN(_15038_));
 MUX2_X2 _41423_ (.A(_15035_),
    .B(_15038_),
    .S(_15025_),
    .Z(\icache.data_mem_data_li [224]));
 AOI21_X1 _41424_ (.A(_15018_),
    .B1(_13935_),
    .B2(_13936_),
    .ZN(_15039_));
 AOI21_X1 _41425_ (.A(_15027_),
    .B1(_13932_),
    .B2(_13933_),
    .ZN(_15040_));
 OR2_X1 _41426_ (.A1(_15039_),
    .A2(_15040_),
    .ZN(_15041_));
 AOI21_X1 _41427_ (.A(_14995_),
    .B1(_13926_),
    .B2(_13929_),
    .ZN(_15042_));
 AOI21_X1 _41428_ (.A(_15003_),
    .B1(_13923_),
    .B2(_13924_),
    .ZN(_15043_));
 OR2_X1 _41429_ (.A1(_15042_),
    .A2(_15043_),
    .ZN(_15044_));
 MUX2_X2 _41430_ (.A(_15041_),
    .B(_15044_),
    .S(_14926_),
    .Z(\icache.data_mem_data_li [225]));
 AOI21_X1 _41431_ (.A(_15018_),
    .B1(_13942_),
    .B2(_13943_),
    .ZN(_15045_));
 AOI21_X1 _41432_ (.A(_15027_),
    .B1(_13939_),
    .B2(_13940_),
    .ZN(_15046_));
 OR2_X2 _41433_ (.A1(_15045_),
    .A2(_15046_),
    .ZN(_15047_));
 AOI21_X1 _41434_ (.A(_14995_),
    .B1(_13950_),
    .B2(_13951_),
    .ZN(_15048_));
 AOI21_X1 _41435_ (.A(_15003_),
    .B1(_13947_),
    .B2(_13948_),
    .ZN(_15049_));
 OR2_X2 _41436_ (.A1(_15048_),
    .A2(_15049_),
    .ZN(_15050_));
 MUX2_X2 _41437_ (.A(_15047_),
    .B(_15050_),
    .S(_15025_),
    .Z(\icache.data_mem_data_li [226]));
 AOI21_X1 _41438_ (.A(_15018_),
    .B1(_13957_),
    .B2(_13958_),
    .ZN(_15051_));
 AOI21_X1 _41439_ (.A(_15027_),
    .B1(_13954_),
    .B2(_13955_),
    .ZN(_15052_));
 OR2_X1 _41440_ (.A1(_15051_),
    .A2(_15052_),
    .ZN(_15053_));
 AOI21_X1 _41441_ (.A(_14995_),
    .B1(_13966_),
    .B2(_13967_),
    .ZN(_15054_));
 AOI21_X1 _41442_ (.A(_15003_),
    .B1(_13962_),
    .B2(_13963_),
    .ZN(_15055_));
 OR2_X2 _41443_ (.A1(_15054_),
    .A2(_15055_),
    .ZN(_15056_));
 MUX2_X2 _41444_ (.A(_15053_),
    .B(_15056_),
    .S(_15025_),
    .Z(\icache.data_mem_data_li [227]));
 AOI21_X1 _41445_ (.A(_15018_),
    .B1(_13982_),
    .B2(_13983_),
    .ZN(_15057_));
 AOI21_X1 _41446_ (.A(_15027_),
    .B1(_13979_),
    .B2(_13980_),
    .ZN(_15058_));
 OR2_X2 _41447_ (.A1(_15057_),
    .A2(_15058_),
    .ZN(_15059_));
 BUF_X4 _41448_ (.A(_11239_),
    .Z(_15060_));
 AOI21_X1 _41449_ (.A(_15060_),
    .B1(_13975_),
    .B2(_13976_),
    .ZN(_15061_));
 AOI21_X1 _41450_ (.A(_15003_),
    .B1(_13970_),
    .B2(_13973_),
    .ZN(_15062_));
 OR2_X2 _41451_ (.A1(_15061_),
    .A2(_15062_),
    .ZN(_15063_));
 MUX2_X2 _41452_ (.A(_15059_),
    .B(_15063_),
    .S(_15025_),
    .Z(\icache.data_mem_data_li [228]));
 AOI21_X1 _41453_ (.A(_15018_),
    .B1(_13997_),
    .B2(_13998_),
    .ZN(_15064_));
 AOI21_X1 _41454_ (.A(_15027_),
    .B1(_13994_),
    .B2(_13995_),
    .ZN(_15065_));
 OR2_X2 _41455_ (.A1(_15064_),
    .A2(_15065_),
    .ZN(_15066_));
 AOI21_X1 _41456_ (.A(_15060_),
    .B1(_13990_),
    .B2(_13991_),
    .ZN(_15067_));
 BUF_X4 _41457_ (.A(_11257_),
    .Z(_15068_));
 AOI21_X1 _41458_ (.A(_15068_),
    .B1(_13986_),
    .B2(_13987_),
    .ZN(_15069_));
 OR2_X2 _41459_ (.A1(_15067_),
    .A2(_15069_),
    .ZN(_15070_));
 MUX2_X2 _41460_ (.A(_15066_),
    .B(_15070_),
    .S(_14926_),
    .Z(\icache.data_mem_data_li [229]));
 AOI21_X1 _41461_ (.A(_15018_),
    .B1(_14014_),
    .B2(_14015_),
    .ZN(_15071_));
 AOI21_X1 _41462_ (.A(_15027_),
    .B1(_14011_),
    .B2(_14012_),
    .ZN(_15072_));
 OR2_X4 _41463_ (.A1(_15071_),
    .A2(_15072_),
    .ZN(_15073_));
 AOI21_X1 _41464_ (.A(_15060_),
    .B1(_14005_),
    .B2(_14008_),
    .ZN(_15074_));
 AOI21_X1 _41465_ (.A(_15068_),
    .B1(_14002_),
    .B2(_14003_),
    .ZN(_15075_));
 OR2_X2 _41466_ (.A1(_15074_),
    .A2(_15075_),
    .ZN(_15076_));
 MUX2_X2 _41467_ (.A(_15073_),
    .B(_15076_),
    .S(_14926_),
    .Z(\icache.data_mem_data_li [230]));
 AOI21_X1 _41468_ (.A(_15018_),
    .B1(_14022_),
    .B2(_14023_),
    .ZN(_15077_));
 AOI21_X1 _41469_ (.A(_15027_),
    .B1(_14018_),
    .B2(_14019_),
    .ZN(_15078_));
 OR2_X4 _41470_ (.A1(_15077_),
    .A2(_15078_),
    .ZN(_15079_));
 AOI21_X1 _41471_ (.A(_15060_),
    .B1(_14029_),
    .B2(_14030_),
    .ZN(_15080_));
 AOI21_X1 _41472_ (.A(_15068_),
    .B1(_14026_),
    .B2(_14027_),
    .ZN(_15081_));
 OR2_X4 _41473_ (.A1(_15080_),
    .A2(_15081_),
    .ZN(_15082_));
 MUX2_X2 _41474_ (.A(_15079_),
    .B(_15082_),
    .S(_15025_),
    .Z(\icache.data_mem_data_li [231]));
 BUF_X8 _41475_ (.A(_08447_),
    .Z(_15083_));
 AOI21_X1 _41476_ (.A(_15083_),
    .B1(_14036_),
    .B2(_14037_),
    .ZN(_15084_));
 AOI21_X1 _41477_ (.A(_15027_),
    .B1(_14033_),
    .B2(_14034_),
    .ZN(_15085_));
 OR2_X4 _41478_ (.A1(_15084_),
    .A2(_15085_),
    .ZN(_15086_));
 AOI21_X1 _41479_ (.A(_15060_),
    .B1(_14044_),
    .B2(_14045_),
    .ZN(_15087_));
 AOI21_X1 _41480_ (.A(_15068_),
    .B1(_14041_),
    .B2(_14042_),
    .ZN(_15088_));
 OR2_X4 _41481_ (.A1(_15087_),
    .A2(_15088_),
    .ZN(_15089_));
 MUX2_X2 _41482_ (.A(_15086_),
    .B(_15089_),
    .S(_14926_),
    .Z(\icache.data_mem_data_li [232]));
 AOI21_X1 _41483_ (.A(_15083_),
    .B1(_14052_),
    .B2(_14053_),
    .ZN(_15090_));
 BUF_X8 _41484_ (.A(_08446_),
    .Z(_15091_));
 AOI21_X1 _41485_ (.A(_15091_),
    .B1(_14049_),
    .B2(_14050_),
    .ZN(_15092_));
 OR2_X4 _41486_ (.A1(_15090_),
    .A2(_15092_),
    .ZN(_15093_));
 AOI21_X1 _41487_ (.A(_15060_),
    .B1(_14061_),
    .B2(_14062_),
    .ZN(_15094_));
 AOI21_X1 _41488_ (.A(_15068_),
    .B1(_14056_),
    .B2(_14059_),
    .ZN(_15095_));
 OR2_X4 _41489_ (.A1(_15094_),
    .A2(_15095_),
    .ZN(_15096_));
 MUX2_X2 _41490_ (.A(_15093_),
    .B(_15096_),
    .S(_15025_),
    .Z(\icache.data_mem_data_li [233]));
 AOI21_X1 _41491_ (.A(_15083_),
    .B1(_14069_),
    .B2(_14070_),
    .ZN(_15097_));
 AOI21_X1 _41492_ (.A(_15091_),
    .B1(_14066_),
    .B2(_14067_),
    .ZN(_15098_));
 OR2_X4 _41493_ (.A1(_15097_),
    .A2(_15098_),
    .ZN(_15099_));
 AOI21_X1 _41494_ (.A(_15060_),
    .B1(_14076_),
    .B2(_14077_),
    .ZN(_15100_));
 AOI21_X1 _41495_ (.A(_15068_),
    .B1(_14073_),
    .B2(_14074_),
    .ZN(_15101_));
 OR2_X4 _41496_ (.A1(_15100_),
    .A2(_15101_),
    .ZN(_15102_));
 MUX2_X2 _41497_ (.A(_15099_),
    .B(_15102_),
    .S(_15025_),
    .Z(\icache.data_mem_data_li [234]));
 AOI21_X1 _41498_ (.A(_15083_),
    .B1(_14085_),
    .B2(_14086_),
    .ZN(_15103_));
 AOI21_X1 _41499_ (.A(_15091_),
    .B1(_14080_),
    .B2(_14083_),
    .ZN(_15104_));
 OR2_X4 _41500_ (.A1(_15103_),
    .A2(_15104_),
    .ZN(_15105_));
 AOI21_X1 _41501_ (.A(_15060_),
    .B1(_14092_),
    .B2(_14093_),
    .ZN(_15106_));
 AOI21_X1 _41502_ (.A(_15068_),
    .B1(_14089_),
    .B2(_14090_),
    .ZN(_15107_));
 OR2_X4 _41503_ (.A1(_15106_),
    .A2(_15107_),
    .ZN(_15108_));
 MUX2_X2 _41504_ (.A(_15105_),
    .B(_15108_),
    .S(_15025_),
    .Z(\icache.data_mem_data_li [235]));
 AOI21_X1 _41505_ (.A(_15083_),
    .B1(_14107_),
    .B2(_14108_),
    .ZN(_15109_));
 AOI21_X1 _41506_ (.A(_15091_),
    .B1(_14104_),
    .B2(_14105_),
    .ZN(_15110_));
 OR2_X4 _41507_ (.A1(_15109_),
    .A2(_15110_),
    .ZN(_15111_));
 AOI21_X1 _41508_ (.A(_15060_),
    .B1(_14099_),
    .B2(_14100_),
    .ZN(_15112_));
 AOI21_X1 _41509_ (.A(_15068_),
    .B1(_14096_),
    .B2(_14097_),
    .ZN(_15113_));
 OR2_X4 _41510_ (.A1(_15112_),
    .A2(_15113_),
    .ZN(_15114_));
 BUF_X16 _41511_ (.A(_13481_),
    .Z(_15115_));
 MUX2_X2 _41512_ (.A(_15111_),
    .B(_15114_),
    .S(_15115_),
    .Z(\icache.data_mem_data_li [236]));
 AOI21_X1 _41513_ (.A(_15083_),
    .B1(_14124_),
    .B2(_14125_),
    .ZN(_15116_));
 AOI21_X1 _41514_ (.A(_15091_),
    .B1(_14120_),
    .B2(_14121_),
    .ZN(_15117_));
 OR2_X4 _41515_ (.A1(_15116_),
    .A2(_15117_),
    .ZN(_15118_));
 AOI21_X1 _41516_ (.A(_15060_),
    .B1(_14116_),
    .B2(_14117_),
    .ZN(_15119_));
 AOI21_X1 _41517_ (.A(_15068_),
    .B1(_14113_),
    .B2(_14114_),
    .ZN(_15120_));
 OR2_X4 _41518_ (.A1(_15119_),
    .A2(_15120_),
    .ZN(_15121_));
 MUX2_X2 _41519_ (.A(_15118_),
    .B(_15121_),
    .S(_15115_),
    .Z(\icache.data_mem_data_li [237]));
 AOI21_X1 _41520_ (.A(_15083_),
    .B1(_14140_),
    .B2(_14141_),
    .ZN(_15122_));
 AOI21_X1 _41521_ (.A(_15091_),
    .B1(_14137_),
    .B2(_14138_),
    .ZN(_15123_));
 OR2_X4 _41522_ (.A1(_15122_),
    .A2(_15123_),
    .ZN(_15124_));
 BUF_X8 _41523_ (.A(_11239_),
    .Z(_15125_));
 AOI21_X1 _41524_ (.A(_15125_),
    .B1(_14133_),
    .B2(_14134_),
    .ZN(_15126_));
 AOI21_X1 _41525_ (.A(_15068_),
    .B1(_14128_),
    .B2(_14131_),
    .ZN(_15127_));
 OR2_X4 _41526_ (.A1(_15126_),
    .A2(_15127_),
    .ZN(_15128_));
 MUX2_X2 _41527_ (.A(_15124_),
    .B(_15128_),
    .S(_15025_),
    .Z(\icache.data_mem_data_li [238]));
 AOI21_X1 _41528_ (.A(_15083_),
    .B1(_14148_),
    .B2(_14149_),
    .ZN(_15129_));
 AOI21_X1 _41529_ (.A(_15091_),
    .B1(_14145_),
    .B2(_14146_),
    .ZN(_15130_));
 OR2_X4 _41530_ (.A1(_15129_),
    .A2(_15130_),
    .ZN(_15131_));
 AOI21_X1 _41531_ (.A(_15125_),
    .B1(_14155_),
    .B2(_14156_),
    .ZN(_15132_));
 BUF_X8 _41532_ (.A(_11257_),
    .Z(_15133_));
 AOI21_X1 _41533_ (.A(_15133_),
    .B1(_14152_),
    .B2(_14153_),
    .ZN(_15134_));
 OR2_X4 _41534_ (.A1(_15132_),
    .A2(_15134_),
    .ZN(_15135_));
 MUX2_X2 _41535_ (.A(_15131_),
    .B(_15135_),
    .S(_15115_),
    .Z(\icache.data_mem_data_li [239]));
 AOI21_X1 _41536_ (.A(_15083_),
    .B1(_14173_),
    .B2(_14174_),
    .ZN(_15136_));
 AOI21_X1 _41537_ (.A(_15091_),
    .B1(_14170_),
    .B2(_14171_),
    .ZN(_15137_));
 OR2_X4 _41538_ (.A1(_15136_),
    .A2(_15137_),
    .ZN(_15138_));
 AOI21_X2 _41539_ (.A(_15125_),
    .B1(_14164_),
    .B2(_14167_),
    .ZN(_15139_));
 AOI21_X1 _41540_ (.A(_15133_),
    .B1(_14161_),
    .B2(_14162_),
    .ZN(_15140_));
 OR2_X4 _41541_ (.A1(_15139_),
    .A2(_15140_),
    .ZN(_15141_));
 BUF_X4 _41542_ (.A(_14816_),
    .Z(_15142_));
 MUX2_X2 _41543_ (.A(_15138_),
    .B(_15141_),
    .S(_15142_),
    .Z(\icache.data_mem_data_li [240]));
 AOI21_X1 _41544_ (.A(_15083_),
    .B1(_14189_),
    .B2(_14190_),
    .ZN(_15143_));
 AOI21_X1 _41545_ (.A(_15091_),
    .B1(_14186_),
    .B2(_14187_),
    .ZN(_15144_));
 OR2_X4 _41546_ (.A1(_15143_),
    .A2(_15144_),
    .ZN(_15145_));
 AOI21_X1 _41547_ (.A(_15125_),
    .B1(_14182_),
    .B2(_14183_),
    .ZN(_15146_));
 AOI21_X1 _41548_ (.A(_15133_),
    .B1(_14177_),
    .B2(_14178_),
    .ZN(_15147_));
 OR2_X4 _41549_ (.A1(_15146_),
    .A2(_15147_),
    .ZN(_15148_));
 MUX2_X2 _41550_ (.A(_15145_),
    .B(_15148_),
    .S(_15115_),
    .Z(\icache.data_mem_data_li [241]));
 BUF_X8 _41551_ (.A(_08447_),
    .Z(_15149_));
 AOI21_X1 _41552_ (.A(_15149_),
    .B1(_14196_),
    .B2(_14197_),
    .ZN(_15150_));
 AOI21_X1 _41553_ (.A(_15091_),
    .B1(_14193_),
    .B2(_14194_),
    .ZN(_15151_));
 OR2_X4 _41554_ (.A1(_15150_),
    .A2(_15151_),
    .ZN(_15152_));
 AOI21_X1 _41555_ (.A(_15125_),
    .B1(_14204_),
    .B2(_14205_),
    .ZN(_15153_));
 AOI21_X2 _41556_ (.A(_15133_),
    .B1(_14201_),
    .B2(_14202_),
    .ZN(_15154_));
 OR2_X4 _41557_ (.A1(_15153_),
    .A2(_15154_),
    .ZN(_15155_));
 MUX2_X2 _41558_ (.A(_15152_),
    .B(_15155_),
    .S(_15142_),
    .Z(\icache.data_mem_data_li [242]));
 AOI21_X1 _41559_ (.A(_15149_),
    .B1(_14211_),
    .B2(_14212_),
    .ZN(_15156_));
 BUF_X8 _41560_ (.A(_08446_),
    .Z(_15157_));
 AOI21_X1 _41561_ (.A(_15157_),
    .B1(_14208_),
    .B2(_14209_),
    .ZN(_15158_));
 OR2_X4 _41562_ (.A1(_15156_),
    .A2(_15158_),
    .ZN(_15159_));
 AOI21_X1 _41563_ (.A(_15125_),
    .B1(_14220_),
    .B2(_14221_),
    .ZN(_15160_));
 AOI21_X2 _41564_ (.A(_15133_),
    .B1(_14215_),
    .B2(_14218_),
    .ZN(_15161_));
 OR2_X4 _41565_ (.A1(_15160_),
    .A2(_15161_),
    .ZN(_15162_));
 MUX2_X2 _41566_ (.A(_15159_),
    .B(_15162_),
    .S(_15142_),
    .Z(\icache.data_mem_data_li [243]));
 AOI21_X1 _41567_ (.A(_15149_),
    .B1(_14235_),
    .B2(_14236_),
    .ZN(_15163_));
 AOI21_X1 _41568_ (.A(_15157_),
    .B1(_14232_),
    .B2(_14233_),
    .ZN(_15164_));
 OR2_X4 _41569_ (.A1(_15163_),
    .A2(_15164_),
    .ZN(_15165_));
 AOI21_X2 _41570_ (.A(_15125_),
    .B1(_14228_),
    .B2(_14229_),
    .ZN(_15166_));
 AOI21_X1 _41571_ (.A(_15133_),
    .B1(_14224_),
    .B2(_14225_),
    .ZN(_15167_));
 OR2_X4 _41572_ (.A1(_15166_),
    .A2(_15167_),
    .ZN(_15168_));
 MUX2_X2 _41573_ (.A(_15165_),
    .B(_15168_),
    .S(_15142_),
    .Z(\icache.data_mem_data_li [244]));
 AOI21_X1 _41574_ (.A(_15149_),
    .B1(_14244_),
    .B2(_14245_),
    .ZN(_15169_));
 AOI21_X1 _41575_ (.A(_15157_),
    .B1(_14239_),
    .B2(_14242_),
    .ZN(_15170_));
 OR2_X4 _41576_ (.A1(_15169_),
    .A2(_15170_),
    .ZN(_15171_));
 AOI21_X1 _41577_ (.A(_15125_),
    .B1(_14251_),
    .B2(_14252_),
    .ZN(_15172_));
 AOI21_X1 _41578_ (.A(_15133_),
    .B1(_14248_),
    .B2(_14249_),
    .ZN(_15173_));
 OR2_X4 _41579_ (.A1(_15172_),
    .A2(_15173_),
    .ZN(_15174_));
 MUX2_X2 _41580_ (.A(_15171_),
    .B(_15174_),
    .S(_15142_),
    .Z(\icache.data_mem_data_li [245]));
 AOI21_X1 _41581_ (.A(_15149_),
    .B1(_14266_),
    .B2(_14267_),
    .ZN(_15175_));
 AOI21_X1 _41582_ (.A(_15157_),
    .B1(_14263_),
    .B2(_14264_),
    .ZN(_15176_));
 OR2_X4 _41583_ (.A1(_15175_),
    .A2(_15176_),
    .ZN(_15177_));
 AOI21_X1 _41584_ (.A(_15125_),
    .B1(_14258_),
    .B2(_14259_),
    .ZN(_15178_));
 AOI21_X1 _41585_ (.A(_15133_),
    .B1(_14255_),
    .B2(_14256_),
    .ZN(_15179_));
 OR2_X4 _41586_ (.A1(_15178_),
    .A2(_15179_),
    .ZN(_15180_));
 MUX2_X2 _41587_ (.A(_15177_),
    .B(_15180_),
    .S(_15115_),
    .Z(\icache.data_mem_data_li [246]));
 AOI21_X1 _41588_ (.A(_15149_),
    .B1(_14273_),
    .B2(_14274_),
    .ZN(_15181_));
 AOI21_X1 _41589_ (.A(_15157_),
    .B1(_14270_),
    .B2(_14271_),
    .ZN(_15182_));
 OR2_X4 _41590_ (.A1(_15181_),
    .A2(_15182_),
    .ZN(_15183_));
 AOI21_X1 _41591_ (.A(_15125_),
    .B1(_14282_),
    .B2(_14283_),
    .ZN(_15184_));
 AOI21_X1 _41592_ (.A(_15133_),
    .B1(_14278_),
    .B2(_14279_),
    .ZN(_15185_));
 OR2_X4 _41593_ (.A1(_15184_),
    .A2(_15185_),
    .ZN(_15186_));
 MUX2_X2 _41594_ (.A(_15183_),
    .B(_15186_),
    .S(_15142_),
    .Z(\icache.data_mem_data_li [247]));
 AOI21_X1 _41595_ (.A(_15149_),
    .B1(_14298_),
    .B2(_14299_),
    .ZN(_15187_));
 AOI21_X1 _41596_ (.A(_15157_),
    .B1(_14295_),
    .B2(_14296_),
    .ZN(_15188_));
 OR2_X4 _41597_ (.A1(_15187_),
    .A2(_15188_),
    .ZN(_15189_));
 AOI21_X1 _41598_ (.A(_11240_),
    .B1(_14291_),
    .B2(_14292_),
    .ZN(_15190_));
 AOI21_X1 _41599_ (.A(_15133_),
    .B1(_14286_),
    .B2(_14289_),
    .ZN(_15191_));
 OR2_X4 _41600_ (.A1(_15190_),
    .A2(_15191_),
    .ZN(_15192_));
 MUX2_X2 _41601_ (.A(_15189_),
    .B(_15192_),
    .S(_15115_),
    .Z(\icache.data_mem_data_li [248]));
 AOI21_X1 _41602_ (.A(_15149_),
    .B1(_14313_),
    .B2(_14314_),
    .ZN(_15193_));
 AOI21_X1 _41603_ (.A(_15157_),
    .B1(_14310_),
    .B2(_14311_),
    .ZN(_15194_));
 OR2_X4 _41604_ (.A1(_15193_),
    .A2(_15194_),
    .ZN(_15195_));
 AOI21_X1 _41605_ (.A(_11240_),
    .B1(_14306_),
    .B2(_14307_),
    .ZN(_15196_));
 AOI21_X2 _41606_ (.A(_11258_),
    .B1(_14302_),
    .B2(_14303_),
    .ZN(_15197_));
 OR2_X4 _41607_ (.A1(_15196_),
    .A2(_15197_),
    .ZN(_15198_));
 MUX2_X2 _41608_ (.A(_15195_),
    .B(_15198_),
    .S(_15142_),
    .Z(\icache.data_mem_data_li [249]));
 AOI21_X2 _41609_ (.A(_15149_),
    .B1(_14330_),
    .B2(_14331_),
    .ZN(_15199_));
 AOI21_X1 _41610_ (.A(_15157_),
    .B1(_14327_),
    .B2(_14328_),
    .ZN(_15200_));
 OR2_X4 _41611_ (.A1(_15199_),
    .A2(_15200_),
    .ZN(_15201_));
 AOI21_X1 _41612_ (.A(_11240_),
    .B1(_14321_),
    .B2(_14324_),
    .ZN(_15202_));
 AOI21_X1 _41613_ (.A(_11258_),
    .B1(_14318_),
    .B2(_14319_),
    .ZN(_15203_));
 OR2_X4 _41614_ (.A1(_15202_),
    .A2(_15203_),
    .ZN(_15204_));
 MUX2_X2 _41615_ (.A(_15201_),
    .B(_15204_),
    .S(_15142_),
    .Z(\icache.data_mem_data_li [250]));
 AOI21_X1 _41616_ (.A(_15149_),
    .B1(_14338_),
    .B2(_14339_),
    .ZN(_15205_));
 AOI21_X1 _41617_ (.A(_15157_),
    .B1(_14334_),
    .B2(_14335_),
    .ZN(_15206_));
 OR2_X4 _41618_ (.A1(_15205_),
    .A2(_15206_),
    .ZN(_15207_));
 AOI21_X1 _41619_ (.A(_11240_),
    .B1(_14345_),
    .B2(_14346_),
    .ZN(_15208_));
 AOI21_X1 _41620_ (.A(_11258_),
    .B1(_14342_),
    .B2(_14343_),
    .ZN(_15209_));
 OR2_X4 _41621_ (.A1(_15208_),
    .A2(_15209_),
    .ZN(_15210_));
 MUX2_X2 _41622_ (.A(_15207_),
    .B(_15210_),
    .S(_15142_),
    .Z(\icache.data_mem_data_li [251]));
 AOI21_X1 _41623_ (.A(_11546_),
    .B1(_14352_),
    .B2(_14353_),
    .ZN(_15211_));
 AOI21_X1 _41624_ (.A(_15157_),
    .B1(_14349_),
    .B2(_14350_),
    .ZN(_15212_));
 OR2_X4 _41625_ (.A1(_15211_),
    .A2(_15212_),
    .ZN(_15213_));
 AOI21_X1 _41626_ (.A(_11240_),
    .B1(_14359_),
    .B2(_14360_),
    .ZN(_15214_));
 AOI21_X1 _41627_ (.A(_11258_),
    .B1(_14356_),
    .B2(_14357_),
    .ZN(_15215_));
 OR2_X4 _41628_ (.A1(_15214_),
    .A2(_15215_),
    .ZN(_15216_));
 MUX2_X2 _41629_ (.A(_15213_),
    .B(_15216_),
    .S(_15142_),
    .Z(\icache.data_mem_data_li [252]));
 AOI21_X1 _41630_ (.A(_11546_),
    .B1(_14374_),
    .B2(_14375_),
    .ZN(_15217_));
 AOI21_X1 _41631_ (.A(_08493_),
    .B1(_14371_),
    .B2(_14372_),
    .ZN(_15218_));
 OR2_X4 _41632_ (.A1(_15217_),
    .A2(_15218_),
    .ZN(_15219_));
 AOI21_X1 _41633_ (.A(_11240_),
    .B1(_14367_),
    .B2(_14368_),
    .ZN(_15220_));
 AOI21_X1 _41634_ (.A(_11258_),
    .B1(_14364_),
    .B2(_14365_),
    .ZN(_15221_));
 OR2_X4 _41635_ (.A1(_15220_),
    .A2(_15221_),
    .ZN(_15222_));
 MUX2_X2 _41636_ (.A(_15219_),
    .B(_15222_),
    .S(_15115_),
    .Z(\icache.data_mem_data_li [253]));
 AOI21_X1 _41637_ (.A(_11546_),
    .B1(_14381_),
    .B2(_14382_),
    .ZN(_15223_));
 AOI21_X1 _41638_ (.A(_08493_),
    .B1(_14378_),
    .B2(_14379_),
    .ZN(_15224_));
 OR2_X4 _41639_ (.A1(_15223_),
    .A2(_15224_),
    .ZN(_15225_));
 AOI21_X1 _41640_ (.A(_11240_),
    .B1(_14388_),
    .B2(_14389_),
    .ZN(_15226_));
 AOI21_X1 _41641_ (.A(_11258_),
    .B1(_14385_),
    .B2(_14386_),
    .ZN(_15227_));
 OR2_X4 _41642_ (.A1(_15226_),
    .A2(_15227_),
    .ZN(_15228_));
 BUF_X16 _41643_ (.A(_14816_),
    .Z(_15229_));
 MUX2_X2 _41644_ (.A(_15225_),
    .B(_15228_),
    .S(_15229_),
    .Z(\icache.data_mem_data_li [254]));
 AOI21_X1 _41645_ (.A(_11546_),
    .B1(_14395_),
    .B2(_14396_),
    .ZN(_15230_));
 AOI21_X1 _41646_ (.A(_08493_),
    .B1(_14392_),
    .B2(_14393_),
    .ZN(_15231_));
 OR2_X4 _41647_ (.A1(_15230_),
    .A2(_15231_),
    .ZN(_15232_));
 AOI21_X2 _41648_ (.A(_11240_),
    .B1(_14402_),
    .B2(_14403_),
    .ZN(_15233_));
 AOI21_X1 _41649_ (.A(_11258_),
    .B1(_14399_),
    .B2(_14400_),
    .ZN(_15234_));
 OR2_X4 _41650_ (.A1(_15233_),
    .A2(_15234_),
    .ZN(_15235_));
 MUX2_X2 _41651_ (.A(_15232_),
    .B(_15235_),
    .S(_15115_),
    .Z(\icache.data_mem_data_li [255]));
 MUX2_X2 _41652_ (.A(_11275_),
    .B(_11291_),
    .S(_15229_),
    .Z(\icache.data_mem_data_li [256]));
 MUX2_X2 _41653_ (.A(_11310_),
    .B(_11327_),
    .S(_15115_),
    .Z(\icache.data_mem_data_li [257]));
 MUX2_X2 _41654_ (.A(_11346_),
    .B(_11363_),
    .S(_15115_),
    .Z(\icache.data_mem_data_li [258]));
 BUF_X16 _41655_ (.A(_13481_),
    .Z(_15236_));
 MUX2_X2 _41656_ (.A(_11380_),
    .B(_11395_),
    .S(_15236_),
    .Z(\icache.data_mem_data_li [259]));
 MUX2_X2 _41657_ (.A(_11412_),
    .B(_11429_),
    .S(_15236_),
    .Z(\icache.data_mem_data_li [260]));
 MUX2_X2 _41658_ (.A(_11447_),
    .B(_11463_),
    .S(_15236_),
    .Z(\icache.data_mem_data_li [261]));
 MUX2_X2 _41659_ (.A(_11481_),
    .B(_11496_),
    .S(_15236_),
    .Z(\icache.data_mem_data_li [262]));
 MUX2_X2 _41660_ (.A(_11514_),
    .B(_11529_),
    .S(_15229_),
    .Z(\icache.data_mem_data_li [263]));
 MUX2_X2 _41661_ (.A(_11545_),
    .B(_11562_),
    .S(_15236_),
    .Z(\icache.data_mem_data_li [264]));
 MUX2_X2 _41662_ (.A(_11581_),
    .B(_11597_),
    .S(_15229_),
    .Z(\icache.data_mem_data_li [265]));
 MUX2_X2 _41663_ (.A(_11613_),
    .B(_11630_),
    .S(_15229_),
    .Z(\icache.data_mem_data_li [266]));
 MUX2_X2 _41664_ (.A(_11649_),
    .B(_11664_),
    .S(_15229_),
    .Z(\icache.data_mem_data_li [267]));
 MUX2_X2 _41665_ (.A(_11686_),
    .B(_11701_),
    .S(_15236_),
    .Z(\icache.data_mem_data_li [268]));
 MUX2_X2 _41666_ (.A(_11719_),
    .B(_11735_),
    .S(_15236_),
    .Z(\icache.data_mem_data_li [269]));
 MUX2_X2 _41667_ (.A(_11752_),
    .B(_11768_),
    .S(_15236_),
    .Z(\icache.data_mem_data_li [270]));
 MUX2_X2 _41668_ (.A(_11787_),
    .B(_11802_),
    .S(_15236_),
    .Z(\icache.data_mem_data_li [271]));
 MUX2_X2 _41669_ (.A(_11819_),
    .B(_11834_),
    .S(_15229_),
    .Z(\icache.data_mem_data_li [272]));
 MUX2_X2 _41670_ (.A(_11854_),
    .B(_11869_),
    .S(_15236_),
    .Z(\icache.data_mem_data_li [273]));
 BUF_X4 _41671_ (.A(_13481_),
    .Z(_15237_));
 MUX2_X2 _41672_ (.A(_11885_),
    .B(_11902_),
    .S(_15237_),
    .Z(\icache.data_mem_data_li [274]));
 MUX2_X2 _41673_ (.A(_11917_),
    .B(_11935_),
    .S(_15237_),
    .Z(\icache.data_mem_data_li [275]));
 MUX2_X2 _41674_ (.A(_11954_),
    .B(_11969_),
    .S(_15229_),
    .Z(\icache.data_mem_data_li [276]));
 MUX2_X2 _41675_ (.A(_11986_),
    .B(_12002_),
    .S(_15237_),
    .Z(\icache.data_mem_data_li [277]));
 MUX2_X2 _41676_ (.A(_12020_),
    .B(_12035_),
    .S(_15229_),
    .Z(\icache.data_mem_data_li [278]));
 MUX2_X2 _41677_ (.A(_12052_),
    .B(_12068_),
    .S(_15237_),
    .Z(\icache.data_mem_data_li [279]));
 MUX2_X2 _41678_ (.A(_12087_),
    .B(_12102_),
    .S(_15237_),
    .Z(\icache.data_mem_data_li [280]));
 MUX2_X2 _41679_ (.A(_12118_),
    .B(_12136_),
    .S(_15237_),
    .Z(\icache.data_mem_data_li [281]));
 MUX2_X2 _41680_ (.A(_12154_),
    .B(_12169_),
    .S(_15237_),
    .Z(\icache.data_mem_data_li [282]));
 MUX2_X2 _41681_ (.A(_12186_),
    .B(_12202_),
    .S(_15237_),
    .Z(\icache.data_mem_data_li [283]));
 MUX2_X2 _41682_ (.A(_12219_),
    .B(_12235_),
    .S(_15237_),
    .Z(\icache.data_mem_data_li [284]));
 MUX2_X2 _41683_ (.A(_12253_),
    .B(_12269_),
    .S(_15237_),
    .Z(\icache.data_mem_data_li [285]));
 BUF_X8 _41684_ (.A(_13481_),
    .Z(_15238_));
 MUX2_X2 _41685_ (.A(_12284_),
    .B(_12303_),
    .S(_15238_),
    .Z(\icache.data_mem_data_li [286]));
 MUX2_X2 _41686_ (.A(_12321_),
    .B(_12336_),
    .S(_15229_),
    .Z(\icache.data_mem_data_li [287]));
 BUF_X32 _41687_ (.A(_14816_),
    .Z(_15239_));
 MUX2_X2 _41688_ (.A(_12357_),
    .B(_12372_),
    .S(_15239_),
    .Z(\icache.data_mem_data_li [288]));
 MUX2_X2 _41689_ (.A(_12389_),
    .B(_12404_),
    .S(_15238_),
    .Z(\icache.data_mem_data_li [289]));
 MUX2_X2 _41690_ (.A(_12420_),
    .B(_12438_),
    .S(_15238_),
    .Z(\icache.data_mem_data_li [290]));
 MUX2_X2 _41691_ (.A(_12454_),
    .B(_12472_),
    .S(_15238_),
    .Z(\icache.data_mem_data_li [291]));
 MUX2_X2 _41692_ (.A(_12490_),
    .B(_12505_),
    .S(_15238_),
    .Z(\icache.data_mem_data_li [292]));
 MUX2_X2 _41693_ (.A(_12523_),
    .B(_12538_),
    .S(_15238_),
    .Z(\icache.data_mem_data_li [293]));
 MUX2_X2 _41694_ (.A(_12554_),
    .B(_12570_),
    .S(_15238_),
    .Z(\icache.data_mem_data_li [294]));
 MUX2_X2 _41695_ (.A(_12588_),
    .B(_12604_),
    .S(_15239_),
    .Z(\icache.data_mem_data_li [295]));
 MUX2_X2 _41696_ (.A(_12624_),
    .B(_12639_),
    .S(_15238_),
    .Z(\icache.data_mem_data_li [296]));
 MUX2_X2 _41697_ (.A(_12659_),
    .B(_12674_),
    .S(_15239_),
    .Z(\icache.data_mem_data_li [297]));
 MUX2_X2 _41698_ (.A(_12694_),
    .B(_12709_),
    .S(_15239_),
    .Z(\icache.data_mem_data_li [298]));
 MUX2_X2 _41699_ (.A(_12726_),
    .B(_12741_),
    .S(_15239_),
    .Z(\icache.data_mem_data_li [299]));
 MUX2_X2 _41700_ (.A(_12758_),
    .B(_12773_),
    .S(_15238_),
    .Z(\icache.data_mem_data_li [300]));
 MUX2_X2 _41701_ (.A(_12792_),
    .B(_12807_),
    .S(_15238_),
    .Z(\icache.data_mem_data_li [301]));
 BUF_X32 _41702_ (.A(_08432_),
    .Z(_15240_));
 BUF_X4 _41703_ (.A(_15240_),
    .Z(_15241_));
 MUX2_X2 _41704_ (.A(_12824_),
    .B(_12839_),
    .S(_15241_),
    .Z(\icache.data_mem_data_li [302]));
 MUX2_X2 _41705_ (.A(_12857_),
    .B(_12872_),
    .S(_15241_),
    .Z(\icache.data_mem_data_li [303]));
 MUX2_X2 _41706_ (.A(_12889_),
    .B(_12905_),
    .S(_15239_),
    .Z(\icache.data_mem_data_li [304]));
 MUX2_X2 _41707_ (.A(_12923_),
    .B(_12939_),
    .S(_15241_),
    .Z(\icache.data_mem_data_li [305]));
 MUX2_X2 _41708_ (.A(_12955_),
    .B(_12972_),
    .S(_15241_),
    .Z(\icache.data_mem_data_li [306]));
 MUX2_X2 _41709_ (.A(_12990_),
    .B(_13006_),
    .S(_15241_),
    .Z(\icache.data_mem_data_li [307]));
 MUX2_X2 _41710_ (.A(_13024_),
    .B(_13039_),
    .S(_15239_),
    .Z(\icache.data_mem_data_li [308]));
 MUX2_X2 _41711_ (.A(_13056_),
    .B(_13072_),
    .S(_15241_),
    .Z(\icache.data_mem_data_li [309]));
 MUX2_X2 _41712_ (.A(_13089_),
    .B(_13105_),
    .S(_15239_),
    .Z(\icache.data_mem_data_li [310]));
 MUX2_X2 _41713_ (.A(_13120_),
    .B(_13137_),
    .S(_15241_),
    .Z(\icache.data_mem_data_li [311]));
 MUX2_X2 _41714_ (.A(_13155_),
    .B(_13170_),
    .S(_15241_),
    .Z(\icache.data_mem_data_li [312]));
 MUX2_X2 _41715_ (.A(_13190_),
    .B(_13205_),
    .S(_15241_),
    .Z(\icache.data_mem_data_li [313]));
 MUX2_X2 _41716_ (.A(_13221_),
    .B(_13237_),
    .S(_15241_),
    .Z(\icache.data_mem_data_li [314]));
 BUF_X32 _41717_ (.A(_15240_),
    .Z(_15242_));
 MUX2_X2 _41718_ (.A(_13253_),
    .B(_13271_),
    .S(_15242_),
    .Z(\icache.data_mem_data_li [315]));
 MUX2_X2 _41719_ (.A(_13286_),
    .B(_13304_),
    .S(_15242_),
    .Z(\icache.data_mem_data_li [316]));
 MUX2_X2 _41720_ (.A(_13320_),
    .B(_13335_),
    .S(_15242_),
    .Z(\icache.data_mem_data_li [317]));
 MUX2_X2 _41721_ (.A(_13355_),
    .B(_13370_),
    .S(_15242_),
    .Z(\icache.data_mem_data_li [318]));
 MUX2_X2 _41722_ (.A(_13386_),
    .B(_13401_),
    .S(_15239_),
    .Z(\icache.data_mem_data_li [319]));
 MUX2_X2 _41723_ (.A(_13408_),
    .B(_13416_),
    .S(_15242_),
    .Z(\icache.data_mem_data_li [320]));
 MUX2_X2 _41724_ (.A(_13425_),
    .B(_13432_),
    .S(_15242_),
    .Z(\icache.data_mem_data_li [321]));
 MUX2_X2 _41725_ (.A(_13440_),
    .B(_13447_),
    .S(_15242_),
    .Z(\icache.data_mem_data_li [322]));
 MUX2_X2 _41726_ (.A(_13456_),
    .B(_13463_),
    .S(_15242_),
    .Z(\icache.data_mem_data_li [323]));
 MUX2_X2 _41727_ (.A(_13471_),
    .B(_13480_),
    .S(_15239_),
    .Z(\icache.data_mem_data_li [324]));
 MUX2_X2 _41728_ (.A(_13490_),
    .B(_13499_),
    .S(_15242_),
    .Z(\icache.data_mem_data_li [325]));
 MUX2_X2 _41729_ (.A(_13508_),
    .B(_13515_),
    .S(_15242_),
    .Z(\icache.data_mem_data_li [326]));
 BUF_X8 _41730_ (.A(_15240_),
    .Z(_15243_));
 MUX2_X2 _41731_ (.A(_13523_),
    .B(_13530_),
    .S(_15243_),
    .Z(\icache.data_mem_data_li [327]));
 BUF_X16 _41732_ (.A(_14816_),
    .Z(_15244_));
 MUX2_X2 _41733_ (.A(_13540_),
    .B(_13547_),
    .S(_15244_),
    .Z(\icache.data_mem_data_li [328]));
 MUX2_X2 _41734_ (.A(_13555_),
    .B(_13562_),
    .S(_15243_),
    .Z(\icache.data_mem_data_li [329]));
 MUX2_X2 _41735_ (.A(_13569_),
    .B(_13577_),
    .S(_15243_),
    .Z(\icache.data_mem_data_li [330]));
 MUX2_X2 _41736_ (.A(_13584_),
    .B(_13593_),
    .S(_15243_),
    .Z(\icache.data_mem_data_li [331]));
 MUX2_X2 _41737_ (.A(_13601_),
    .B(_13608_),
    .S(_15243_),
    .Z(\icache.data_mem_data_li [332]));
 MUX2_X2 _41738_ (.A(_13617_),
    .B(_13624_),
    .S(_15243_),
    .Z(\icache.data_mem_data_li [333]));
 MUX2_X2 _41739_ (.A(_13631_),
    .B(_13639_),
    .S(_15244_),
    .Z(\icache.data_mem_data_li [334]));
 MUX2_X2 _41740_ (.A(_13646_),
    .B(_13655_),
    .S(_15244_),
    .Z(\icache.data_mem_data_li [335]));
 MUX2_X2 _41741_ (.A(_13664_),
    .B(_13671_),
    .S(_15244_),
    .Z(\icache.data_mem_data_li [336]));
 MUX2_X2 _41742_ (.A(_13679_),
    .B(_13686_),
    .S(_15243_),
    .Z(\icache.data_mem_data_li [337]));
 MUX2_X2 _41743_ (.A(_13696_),
    .B(_13703_),
    .S(_15243_),
    .Z(\icache.data_mem_data_li [338]));
 MUX2_X2 _41744_ (.A(_13712_),
    .B(_13719_),
    .S(_15243_),
    .Z(\icache.data_mem_data_li [339]));
 MUX2_X2 _41745_ (.A(_13727_),
    .B(_13734_),
    .S(_15244_),
    .Z(\icache.data_mem_data_li [340]));
 MUX2_X2 _41746_ (.A(_13741_),
    .B(_13750_),
    .S(_15243_),
    .Z(\icache.data_mem_data_li [341]));
 BUF_X4 _41747_ (.A(_15240_),
    .Z(_15245_));
 MUX2_X2 _41748_ (.A(_13758_),
    .B(_13765_),
    .S(_15245_),
    .Z(\icache.data_mem_data_li [342]));
 MUX2_X2 _41749_ (.A(_13774_),
    .B(_13781_),
    .S(_15245_),
    .Z(\icache.data_mem_data_li [343]));
 MUX2_X2 _41750_ (.A(_13788_),
    .B(_13796_),
    .S(_15245_),
    .Z(\icache.data_mem_data_li [344]));
 MUX2_X2 _41751_ (.A(_13804_),
    .B(_13812_),
    .S(_15244_),
    .Z(\icache.data_mem_data_li [345]));
 MUX2_X2 _41752_ (.A(_13821_),
    .B(_13828_),
    .S(_15244_),
    .Z(\icache.data_mem_data_li [346]));
 MUX2_X2 _41753_ (.A(_13836_),
    .B(_13843_),
    .S(_15245_),
    .Z(\icache.data_mem_data_li [347]));
 MUX2_X2 _41754_ (.A(_13853_),
    .B(_13860_),
    .S(_15245_),
    .Z(\icache.data_mem_data_li [348]));
 MUX2_X2 _41755_ (.A(_13868_),
    .B(_13875_),
    .S(_15245_),
    .Z(\icache.data_mem_data_li [349]));
 MUX2_X2 _41756_ (.A(_13882_),
    .B(_13890_),
    .S(_15245_),
    .Z(\icache.data_mem_data_li [350]));
 MUX2_X2 _41757_ (.A(_13897_),
    .B(_13906_),
    .S(_15244_),
    .Z(\icache.data_mem_data_li [351]));
 MUX2_X2 _41758_ (.A(_13914_),
    .B(_13921_),
    .S(_15245_),
    .Z(\icache.data_mem_data_li [352]));
 MUX2_X2 _41759_ (.A(_13931_),
    .B(_13938_),
    .S(_15245_),
    .Z(\icache.data_mem_data_li [353]));
 MUX2_X2 _41760_ (.A(_13945_),
    .B(_13953_),
    .S(_15245_),
    .Z(\icache.data_mem_data_li [354]));
 BUF_X8 _41761_ (.A(_15240_),
    .Z(_15246_));
 MUX2_X2 _41762_ (.A(_13960_),
    .B(_13969_),
    .S(_15246_),
    .Z(\icache.data_mem_data_li [355]));
 MUX2_X2 _41763_ (.A(_13978_),
    .B(_13985_),
    .S(_15244_),
    .Z(\icache.data_mem_data_li [356]));
 MUX2_X2 _41764_ (.A(_13993_),
    .B(_14000_),
    .S(_15246_),
    .Z(\icache.data_mem_data_li [357]));
 MUX2_X2 _41765_ (.A(_14010_),
    .B(_14017_),
    .S(_15246_),
    .Z(\icache.data_mem_data_li [358]));
 MUX2_X2 _41766_ (.A(_14025_),
    .B(_14032_),
    .S(_15246_),
    .Z(\icache.data_mem_data_li [359]));
 MUX2_X2 _41767_ (.A(_14039_),
    .B(_14047_),
    .S(_15244_),
    .Z(\icache.data_mem_data_li [360]));
 MUX2_X2 _41768_ (.A(_14055_),
    .B(_14064_),
    .S(_15246_),
    .Z(\icache.data_mem_data_li [361]));
 MUX2_X2 _41769_ (.A(_14072_),
    .B(_14079_),
    .S(_15246_),
    .Z(\icache.data_mem_data_li [362]));
 MUX2_X2 _41770_ (.A(_14088_),
    .B(_14095_),
    .S(_15246_),
    .Z(\icache.data_mem_data_li [363]));
 MUX2_X2 _41771_ (.A(_14102_),
    .B(_14110_),
    .S(_15246_),
    .Z(\icache.data_mem_data_li [364]));
 MUX2_X2 _41772_ (.A(_14119_),
    .B(_14127_),
    .S(_15246_),
    .Z(\icache.data_mem_data_li [365]));
 BUF_X32 _41773_ (.A(_14816_),
    .Z(_15247_));
 MUX2_X2 _41774_ (.A(_14136_),
    .B(_14143_),
    .S(_15247_),
    .Z(\icache.data_mem_data_li [366]));
 MUX2_X2 _41775_ (.A(_14151_),
    .B(_14158_),
    .S(_15247_),
    .Z(\icache.data_mem_data_li [367]));
 MUX2_X2 _41776_ (.A(_14169_),
    .B(_14176_),
    .S(_15247_),
    .Z(\icache.data_mem_data_li [368]));
 MUX2_X2 _41777_ (.A(_14185_),
    .B(_14192_),
    .S(_15246_),
    .Z(\icache.data_mem_data_li [369]));
 BUF_X8 _41778_ (.A(_15240_),
    .Z(_15248_));
 MUX2_X2 _41779_ (.A(_14199_),
    .B(_14207_),
    .S(_15248_),
    .Z(\icache.data_mem_data_li [370]));
 MUX2_X2 _41780_ (.A(_14214_),
    .B(_14223_),
    .S(_15248_),
    .Z(\icache.data_mem_data_li [371]));
 MUX2_X2 _41781_ (.A(_14231_),
    .B(_14238_),
    .S(_15247_),
    .Z(\icache.data_mem_data_li [372]));
 MUX2_X2 _41782_ (.A(_14247_),
    .B(_14254_),
    .S(_15248_),
    .Z(\icache.data_mem_data_li [373]));
 MUX2_X2 _41783_ (.A(_14261_),
    .B(_14269_),
    .S(_15248_),
    .Z(\icache.data_mem_data_li [374]));
 MUX2_X2 _41784_ (.A(_14276_),
    .B(_14285_),
    .S(_15248_),
    .Z(\icache.data_mem_data_li [375]));
 MUX2_X2 _41785_ (.A(_14294_),
    .B(_14301_),
    .S(_15248_),
    .Z(\icache.data_mem_data_li [376]));
 MUX2_X2 _41786_ (.A(_14309_),
    .B(_14316_),
    .S(_15247_),
    .Z(\icache.data_mem_data_li [377]));
 MUX2_X2 _41787_ (.A(_14326_),
    .B(_14333_),
    .S(_15247_),
    .Z(\icache.data_mem_data_li [378]));
 MUX2_X2 _41788_ (.A(_14341_),
    .B(_14348_),
    .S(_15248_),
    .Z(\icache.data_mem_data_li [379]));
 MUX2_X2 _41789_ (.A(_14355_),
    .B(_14362_),
    .S(_15248_),
    .Z(\icache.data_mem_data_li [380]));
 MUX2_X2 _41790_ (.A(_14370_),
    .B(_14377_),
    .S(_15248_),
    .Z(\icache.data_mem_data_li [381]));
 MUX2_X2 _41791_ (.A(_14384_),
    .B(_14391_),
    .S(_15248_),
    .Z(\icache.data_mem_data_li [382]));
 MUX2_X2 _41792_ (.A(_14398_),
    .B(_14405_),
    .S(_15247_),
    .Z(\icache.data_mem_data_li [383]));
 BUF_X16 _41793_ (.A(_15240_),
    .Z(_15249_));
 MUX2_X2 _41794_ (.A(_14408_),
    .B(_14412_),
    .S(_15249_),
    .Z(\icache.data_mem_data_li [384]));
 MUX2_X2 _41795_ (.A(_14415_),
    .B(_14419_),
    .S(_15247_),
    .Z(\icache.data_mem_data_li [385]));
 MUX2_X2 _41796_ (.A(_14422_),
    .B(_14425_),
    .S(_15249_),
    .Z(\icache.data_mem_data_li [386]));
 MUX2_X2 _41797_ (.A(_14428_),
    .B(_14431_),
    .S(_15249_),
    .Z(\icache.data_mem_data_li [387]));
 MUX2_X2 _41798_ (.A(_14435_),
    .B(_14438_),
    .S(_15249_),
    .Z(\icache.data_mem_data_li [388]));
 MUX2_X2 _41799_ (.A(_14442_),
    .B(_14445_),
    .S(_15247_),
    .Z(\icache.data_mem_data_li [389]));
 MUX2_X2 _41800_ (.A(_14448_),
    .B(_14451_),
    .S(_15247_),
    .Z(\icache.data_mem_data_li [390]));
 MUX2_X2 _41801_ (.A(_14455_),
    .B(_14458_),
    .S(_15249_),
    .Z(\icache.data_mem_data_li [391]));
 BUF_X8 _41802_ (.A(_14816_),
    .Z(_15250_));
 MUX2_X2 _41803_ (.A(_14461_),
    .B(_14464_),
    .S(_15250_),
    .Z(\icache.data_mem_data_li [392]));
 MUX2_X2 _41804_ (.A(_14467_),
    .B(_14470_),
    .S(_15249_),
    .Z(\icache.data_mem_data_li [393]));
 MUX2_X2 _41805_ (.A(_14473_),
    .B(_14477_),
    .S(_15250_),
    .Z(\icache.data_mem_data_li [394]));
 MUX2_X2 _41806_ (.A(_14480_),
    .B(_14484_),
    .S(_15249_),
    .Z(\icache.data_mem_data_li [395]));
 MUX2_X2 _41807_ (.A(_14487_),
    .B(_14490_),
    .S(_15250_),
    .Z(\icache.data_mem_data_li [396]));
 MUX2_X2 _41808_ (.A(_14493_),
    .B(_14496_),
    .S(_15250_),
    .Z(\icache.data_mem_data_li [397]));
 MUX2_X2 _41809_ (.A(_14500_),
    .B(_14503_),
    .S(_15249_),
    .Z(\icache.data_mem_data_li [398]));
 MUX2_X2 _41810_ (.A(_14508_),
    .B(_14511_),
    .S(_15250_),
    .Z(\icache.data_mem_data_li [399]));
 MUX2_X2 _41811_ (.A(_14514_),
    .B(_14517_),
    .S(_15249_),
    .Z(\icache.data_mem_data_li [400]));
 MUX2_X2 _41812_ (.A(_14520_),
    .B(_14523_),
    .S(_15250_),
    .Z(\icache.data_mem_data_li [401]));
 MUX2_X2 _41813_ (.A(_14526_),
    .B(_14529_),
    .S(_15249_),
    .Z(\icache.data_mem_data_li [402]));
 BUF_X8 _41814_ (.A(_15240_),
    .Z(_15251_));
 MUX2_X2 _41815_ (.A(_14532_),
    .B(_14535_),
    .S(_15251_),
    .Z(\icache.data_mem_data_li [403]));
 MUX2_X2 _41816_ (.A(_14538_),
    .B(_14542_),
    .S(_15251_),
    .Z(\icache.data_mem_data_li [404]));
 MUX2_X2 _41817_ (.A(_14545_),
    .B(_14549_),
    .S(_15251_),
    .Z(\icache.data_mem_data_li [405]));
 MUX2_X2 _41818_ (.A(_14552_),
    .B(_14555_),
    .S(_15250_),
    .Z(\icache.data_mem_data_li [406]));
 MUX2_X2 _41819_ (.A(_14558_),
    .B(_14561_),
    .S(_15251_),
    .Z(\icache.data_mem_data_li [407]));
 MUX2_X2 _41820_ (.A(_14565_),
    .B(_14568_),
    .S(_15250_),
    .Z(\icache.data_mem_data_li [408]));
 MUX2_X2 _41821_ (.A(_14572_),
    .B(_14575_),
    .S(_15251_),
    .Z(\icache.data_mem_data_li [409]));
 MUX2_X2 _41822_ (.A(_14578_),
    .B(_14581_),
    .S(_15251_),
    .Z(\icache.data_mem_data_li [410]));
 MUX2_X2 _41823_ (.A(_14584_),
    .B(_14587_),
    .S(_15251_),
    .Z(\icache.data_mem_data_li [411]));
 MUX2_X2 _41824_ (.A(_14590_),
    .B(_14593_),
    .S(_15251_),
    .Z(\icache.data_mem_data_li [412]));
 MUX2_X2 _41825_ (.A(_14597_),
    .B(_14600_),
    .S(_15250_),
    .Z(\icache.data_mem_data_li [413]));
 MUX2_X2 _41826_ (.A(_14603_),
    .B(_14607_),
    .S(_15251_),
    .Z(\icache.data_mem_data_li [414]));
 MUX2_X2 _41827_ (.A(_14610_),
    .B(_14614_),
    .S(_15250_),
    .Z(\icache.data_mem_data_li [415]));
 MUX2_X2 _41828_ (.A(_14618_),
    .B(_14621_),
    .S(_15251_),
    .Z(\icache.data_mem_data_li [416]));
 BUF_X8 _41829_ (.A(_14816_),
    .Z(_15252_));
 MUX2_X2 _41830_ (.A(_14624_),
    .B(_14627_),
    .S(_15252_),
    .Z(\icache.data_mem_data_li [417]));
 BUF_X8 _41831_ (.A(_15240_),
    .Z(_15253_));
 MUX2_X2 _41832_ (.A(_14631_),
    .B(_14634_),
    .S(_15253_),
    .Z(\icache.data_mem_data_li [418]));
 MUX2_X2 _41833_ (.A(_14638_),
    .B(_14641_),
    .S(_15253_),
    .Z(\icache.data_mem_data_li [419]));
 MUX2_X2 _41834_ (.A(_14644_),
    .B(_14647_),
    .S(_15253_),
    .Z(\icache.data_mem_data_li [420]));
 MUX2_X2 _41835_ (.A(_14650_),
    .B(_14653_),
    .S(_15252_),
    .Z(\icache.data_mem_data_li [421]));
 MUX2_X2 _41836_ (.A(_14656_),
    .B(_14659_),
    .S(_15252_),
    .Z(\icache.data_mem_data_li [422]));
 MUX2_X2 _41837_ (.A(_14662_),
    .B(_14665_),
    .S(_15253_),
    .Z(\icache.data_mem_data_li [423]));
 MUX2_X2 _41838_ (.A(_14668_),
    .B(_14672_),
    .S(_15252_),
    .Z(\icache.data_mem_data_li [424]));
 MUX2_X2 _41839_ (.A(_14675_),
    .B(_14679_),
    .S(_15253_),
    .Z(\icache.data_mem_data_li [425]));
 MUX2_X2 _41840_ (.A(_14682_),
    .B(_14685_),
    .S(_15252_),
    .Z(\icache.data_mem_data_li [426]));
 MUX2_X2 _41841_ (.A(_14688_),
    .B(_14691_),
    .S(_15253_),
    .Z(\icache.data_mem_data_li [427]));
 MUX2_X2 _41842_ (.A(_14695_),
    .B(_14698_),
    .S(_15252_),
    .Z(\icache.data_mem_data_li [428]));
 MUX2_X2 _41843_ (.A(_14702_),
    .B(_14705_),
    .S(_15252_),
    .Z(\icache.data_mem_data_li [429]));
 MUX2_X2 _41844_ (.A(_14708_),
    .B(_14711_),
    .S(_15253_),
    .Z(\icache.data_mem_data_li [430]));
 MUX2_X2 _41845_ (.A(_14714_),
    .B(_14717_),
    .S(_15252_),
    .Z(\icache.data_mem_data_li [431]));
 MUX2_X2 _41846_ (.A(_14720_),
    .B(_14723_),
    .S(_15253_),
    .Z(\icache.data_mem_data_li [432]));
 MUX2_X2 _41847_ (.A(_14727_),
    .B(_14730_),
    .S(_15252_),
    .Z(\icache.data_mem_data_li [433]));
 MUX2_X2 _41848_ (.A(_14733_),
    .B(_14737_),
    .S(_15253_),
    .Z(\icache.data_mem_data_li [434]));
 MUX2_X2 _41849_ (.A(_14740_),
    .B(_14744_),
    .S(_15253_),
    .Z(\icache.data_mem_data_li [435]));
 BUF_X8 _41850_ (.A(_15240_),
    .Z(_15254_));
 MUX2_X2 _41851_ (.A(_14747_),
    .B(_14750_),
    .S(_15254_),
    .Z(\icache.data_mem_data_li [436]));
 MUX2_X2 _41852_ (.A(_14753_),
    .B(_14756_),
    .S(_15254_),
    .Z(\icache.data_mem_data_li [437]));
 MUX2_X2 _41853_ (.A(_14760_),
    .B(_14763_),
    .S(_15252_),
    .Z(\icache.data_mem_data_li [438]));
 MUX2_X2 _41854_ (.A(_14768_),
    .B(_14771_),
    .S(_15254_),
    .Z(\icache.data_mem_data_li [439]));
 BUF_X8 _41855_ (.A(_08431_),
    .Z(_15255_));
 MUX2_X2 _41856_ (.A(_14774_),
    .B(_14777_),
    .S(_15255_),
    .Z(\icache.data_mem_data_li [440]));
 MUX2_X2 _41857_ (.A(_14780_),
    .B(_14783_),
    .S(_15254_),
    .Z(\icache.data_mem_data_li [441]));
 MUX2_X2 _41858_ (.A(_14786_),
    .B(_14789_),
    .S(_15254_),
    .Z(\icache.data_mem_data_li [442]));
 MUX2_X2 _41859_ (.A(_14792_),
    .B(_14795_),
    .S(_15254_),
    .Z(\icache.data_mem_data_li [443]));
 MUX2_X2 _41860_ (.A(_14798_),
    .B(_14802_),
    .S(_15254_),
    .Z(\icache.data_mem_data_li [444]));
 MUX2_X2 _41861_ (.A(_14805_),
    .B(_14809_),
    .S(_15255_),
    .Z(\icache.data_mem_data_li [445]));
 MUX2_X2 _41862_ (.A(_14812_),
    .B(_14815_),
    .S(_15254_),
    .Z(\icache.data_mem_data_li [446]));
 MUX2_X2 _41863_ (.A(_14820_),
    .B(_14823_),
    .S(_15255_),
    .Z(\icache.data_mem_data_li [447]));
 MUX2_X2 _41864_ (.A(_14827_),
    .B(_14830_),
    .S(_15254_),
    .Z(\icache.data_mem_data_li [448]));
 MUX2_X2 _41865_ (.A(_14834_),
    .B(_14837_),
    .S(_15255_),
    .Z(\icache.data_mem_data_li [449]));
 MUX2_X2 _41866_ (.A(_14840_),
    .B(_14843_),
    .S(_15254_),
    .Z(\icache.data_mem_data_li [450]));
 BUF_X8 _41867_ (.A(_08432_),
    .Z(_15256_));
 MUX2_X2 _41868_ (.A(_14846_),
    .B(_14849_),
    .S(_15256_),
    .Z(\icache.data_mem_data_li [451]));
 MUX2_X2 _41869_ (.A(_14852_),
    .B(_14855_),
    .S(_15256_),
    .Z(\icache.data_mem_data_li [452]));
 MUX2_X2 _41870_ (.A(_14858_),
    .B(_14861_),
    .S(_15255_),
    .Z(\icache.data_mem_data_li [453]));
 MUX2_X2 _41871_ (.A(_14864_),
    .B(_14868_),
    .S(_15255_),
    .Z(\icache.data_mem_data_li [454]));
 MUX2_X2 _41872_ (.A(_14871_),
    .B(_14875_),
    .S(_15256_),
    .Z(\icache.data_mem_data_li [455]));
 MUX2_X2 _41873_ (.A(_14878_),
    .B(_14881_),
    .S(_15255_),
    .Z(\icache.data_mem_data_li [456]));
 MUX2_X2 _41874_ (.A(_14884_),
    .B(_14887_),
    .S(_15256_),
    .Z(\icache.data_mem_data_li [457]));
 MUX2_X2 _41875_ (.A(_14891_),
    .B(_14894_),
    .S(_15256_),
    .Z(\icache.data_mem_data_li [458]));
 MUX2_X2 _41876_ (.A(_14898_),
    .B(_14901_),
    .S(_15256_),
    .Z(\icache.data_mem_data_li [459]));
 MUX2_X2 _41877_ (.A(_14904_),
    .B(_14907_),
    .S(_15255_),
    .Z(\icache.data_mem_data_li [460]));
 MUX2_X2 _41878_ (.A(_14910_),
    .B(_14913_),
    .S(_15255_),
    .Z(\icache.data_mem_data_li [461]));
 MUX2_X2 _41879_ (.A(_14916_),
    .B(_14919_),
    .S(_15256_),
    .Z(\icache.data_mem_data_li [462]));
 MUX2_X2 _41880_ (.A(_14922_),
    .B(_14925_),
    .S(_15255_),
    .Z(\icache.data_mem_data_li [463]));
 MUX2_X2 _41881_ (.A(_14929_),
    .B(_14933_),
    .S(_15256_),
    .Z(\icache.data_mem_data_li [464]));
 BUF_X8 _41882_ (.A(_08431_),
    .Z(_15257_));
 MUX2_X2 _41883_ (.A(_14937_),
    .B(_14941_),
    .S(_15257_),
    .Z(\icache.data_mem_data_li [465]));
 MUX2_X2 _41884_ (.A(_14944_),
    .B(_14947_),
    .S(_15256_),
    .Z(\icache.data_mem_data_li [466]));
 MUX2_X2 _41885_ (.A(_14950_),
    .B(_14953_),
    .S(_15256_),
    .Z(\icache.data_mem_data_li [467]));
 BUF_X4 _41886_ (.A(_08432_),
    .Z(_15258_));
 MUX2_X2 _41887_ (.A(_14957_),
    .B(_14960_),
    .S(_15258_),
    .Z(\icache.data_mem_data_li [468]));
 MUX2_X2 _41888_ (.A(_14964_),
    .B(_14967_),
    .S(_15258_),
    .Z(\icache.data_mem_data_li [469]));
 MUX2_X2 _41889_ (.A(_14970_),
    .B(_14973_),
    .S(_15257_),
    .Z(\icache.data_mem_data_li [470]));
 MUX2_X2 _41890_ (.A(_14976_),
    .B(_14979_),
    .S(_15258_),
    .Z(\icache.data_mem_data_li [471]));
 MUX2_X2 _41891_ (.A(_14982_),
    .B(_14985_),
    .S(_15257_),
    .Z(\icache.data_mem_data_li [472]));
 MUX2_X2 _41892_ (.A(_14988_),
    .B(_14991_),
    .S(_15258_),
    .Z(\icache.data_mem_data_li [473]));
 MUX2_X2 _41893_ (.A(_14994_),
    .B(_14998_),
    .S(_15258_),
    .Z(\icache.data_mem_data_li [474]));
 MUX2_X2 _41894_ (.A(_15001_),
    .B(_15005_),
    .S(_15258_),
    .Z(\icache.data_mem_data_li [475]));
 MUX2_X2 _41895_ (.A(_15008_),
    .B(_15011_),
    .S(_15258_),
    .Z(\icache.data_mem_data_li [476]));
 MUX2_X2 _41896_ (.A(_15014_),
    .B(_15017_),
    .S(_15257_),
    .Z(\icache.data_mem_data_li [477]));
 MUX2_X2 _41897_ (.A(_15021_),
    .B(_15024_),
    .S(_15258_),
    .Z(\icache.data_mem_data_li [478]));
 MUX2_X2 _41898_ (.A(_15029_),
    .B(_15032_),
    .S(_15257_),
    .Z(\icache.data_mem_data_li [479]));
 MUX2_X2 _41899_ (.A(_15035_),
    .B(_15038_),
    .S(_15258_),
    .Z(\icache.data_mem_data_li [480]));
 MUX2_X2 _41900_ (.A(_15041_),
    .B(_15044_),
    .S(_15257_),
    .Z(\icache.data_mem_data_li [481]));
 MUX2_X2 _41901_ (.A(_15047_),
    .B(_15050_),
    .S(_15258_),
    .Z(\icache.data_mem_data_li [482]));
 BUF_X8 _41902_ (.A(_08432_),
    .Z(_15259_));
 MUX2_X2 _41903_ (.A(_15053_),
    .B(_15056_),
    .S(_15259_),
    .Z(\icache.data_mem_data_li [483]));
 MUX2_X2 _41904_ (.A(_15059_),
    .B(_15063_),
    .S(_15259_),
    .Z(\icache.data_mem_data_li [484]));
 MUX2_X2 _41905_ (.A(_15066_),
    .B(_15070_),
    .S(_15257_),
    .Z(\icache.data_mem_data_li [485]));
 MUX2_X2 _41906_ (.A(_15073_),
    .B(_15076_),
    .S(_15257_),
    .Z(\icache.data_mem_data_li [486]));
 MUX2_X2 _41907_ (.A(_15079_),
    .B(_15082_),
    .S(_15259_),
    .Z(\icache.data_mem_data_li [487]));
 MUX2_X2 _41908_ (.A(_15086_),
    .B(_15089_),
    .S(_15257_),
    .Z(\icache.data_mem_data_li [488]));
 MUX2_X2 _41909_ (.A(_15093_),
    .B(_15096_),
    .S(_15259_),
    .Z(\icache.data_mem_data_li [489]));
 MUX2_X2 _41910_ (.A(_15099_),
    .B(_15102_),
    .S(_15259_),
    .Z(\icache.data_mem_data_li [490]));
 MUX2_X2 _41911_ (.A(_15105_),
    .B(_15108_),
    .S(_15259_),
    .Z(\icache.data_mem_data_li [491]));
 MUX2_X2 _41912_ (.A(_15111_),
    .B(_15114_),
    .S(_15257_),
    .Z(\icache.data_mem_data_li [492]));
 MUX2_X2 _41913_ (.A(_15118_),
    .B(_15121_),
    .S(_08495_),
    .Z(\icache.data_mem_data_li [493]));
 MUX2_X2 _41914_ (.A(_15124_),
    .B(_15128_),
    .S(_15259_),
    .Z(\icache.data_mem_data_li [494]));
 MUX2_X2 _41915_ (.A(_15131_),
    .B(_15135_),
    .S(_08495_),
    .Z(\icache.data_mem_data_li [495]));
 MUX2_X2 _41916_ (.A(_15138_),
    .B(_15141_),
    .S(_15259_),
    .Z(\icache.data_mem_data_li [496]));
 MUX2_X2 _41917_ (.A(_15145_),
    .B(_15148_),
    .S(_08495_),
    .Z(\icache.data_mem_data_li [497]));
 MUX2_X2 _41918_ (.A(_15152_),
    .B(_15155_),
    .S(_15259_),
    .Z(\icache.data_mem_data_li [498]));
 MUX2_X2 _41919_ (.A(_15159_),
    .B(_15162_),
    .S(_15259_),
    .Z(\icache.data_mem_data_li [499]));
 MUX2_X2 _41920_ (.A(_15165_),
    .B(_15168_),
    .S(_08433_),
    .Z(\icache.data_mem_data_li [500]));
 MUX2_X2 _41921_ (.A(_15171_),
    .B(_15174_),
    .S(_08433_),
    .Z(\icache.data_mem_data_li [501]));
 MUX2_X2 _41922_ (.A(_15177_),
    .B(_15180_),
    .S(_08495_),
    .Z(\icache.data_mem_data_li [502]));
 MUX2_X2 _41923_ (.A(_15183_),
    .B(_15186_),
    .S(_08433_),
    .Z(\icache.data_mem_data_li [503]));
 MUX2_X2 _41924_ (.A(_15189_),
    .B(_15192_),
    .S(_08495_),
    .Z(\icache.data_mem_data_li [504]));
 MUX2_X2 _41925_ (.A(_15195_),
    .B(_15198_),
    .S(_08433_),
    .Z(\icache.data_mem_data_li [505]));
 MUX2_X2 _41926_ (.A(_15201_),
    .B(_15204_),
    .S(_08433_),
    .Z(\icache.data_mem_data_li [506]));
 MUX2_X2 _41927_ (.A(_15207_),
    .B(_15210_),
    .S(_08433_),
    .Z(\icache.data_mem_data_li [507]));
 MUX2_X2 _41928_ (.A(_15213_),
    .B(_15216_),
    .S(_08433_),
    .Z(\icache.data_mem_data_li [508]));
 MUX2_X2 _41929_ (.A(_15219_),
    .B(_15222_),
    .S(_08495_),
    .Z(\icache.data_mem_data_li [509]));
 MUX2_X2 _41930_ (.A(_15225_),
    .B(_15228_),
    .S(_08433_),
    .Z(\icache.data_mem_data_li [510]));
 MUX2_X2 _41931_ (.A(_15232_),
    .B(_15235_),
    .S(_08495_),
    .Z(\icache.data_mem_data_li [511]));
 AND2_X1 _41932_ (.A1(_07618_),
    .A2(_07978_),
    .ZN(_15260_));
 INV_X1 _41933_ (.A(_10734_),
    .ZN(_15261_));
 OAI21_X1 _41934_ (.A(_15260_),
    .B1(_15261_),
    .B2(\icache.lce.lce_cmd_inst.syn_ack_cnt_r ),
    .ZN(_15262_));
 INV_X1 _41935_ (.A(_15260_),
    .ZN(_15263_));
 AOI21_X1 _41936_ (.A(_07605_),
    .B1(_15263_),
    .B2(_00599_),
    .ZN(_15264_));
 AND2_X1 _41937_ (.A1(_15262_),
    .A2(_15264_),
    .ZN(_15265_));
 MUX2_X1 _41938_ (.A(_15265_),
    .B(lce_data_cmd_ready_i),
    .S(_07608_),
    .Z(_15266_));
 INV_X1 _41939_ (.A(_08497_),
    .ZN(_15267_));
 NAND2_X1 _41940_ (.A1(_08424_),
    .A2(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [3]),
    .ZN(_15268_));
 NAND2_X1 _41941_ (.A1(net1396),
    .A2(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [521]),
    .ZN(_15269_));
 NAND2_X4 _41942_ (.A1(_15268_),
    .A2(_15269_),
    .ZN(_15270_));
 NAND2_X1 _41943_ (.A1(_08424_),
    .A2(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [4]),
    .ZN(_15271_));
 NAND2_X1 _41944_ (.A1(net1393),
    .A2(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [522]),
    .ZN(_15272_));
 AOI21_X1 _41945_ (.A(_15270_),
    .B1(_15271_),
    .B2(_15272_),
    .ZN(_15273_));
 AND2_X2 _41946_ (.A1(_15273_),
    .A2(_00075_),
    .ZN(_15274_));
 INV_X1 _41947_ (.A(_15274_),
    .ZN(_15275_));
 NOR2_X1 _41948_ (.A1(_08499_),
    .A2(_15275_),
    .ZN(_15276_));
 INV_X1 _41949_ (.A(_15276_),
    .ZN(_15277_));
 AND2_X2 _41950_ (.A1(_08037_),
    .A2(_15277_),
    .ZN(_15278_));
 AOI21_X2 _41951_ (.A(_00075_),
    .B1(_08497_),
    .B2(_10726_),
    .ZN(_15279_));
 NOR2_X1 _41952_ (.A1(_15278_),
    .A2(_15279_),
    .ZN(_15280_));
 INV_X1 _41953_ (.A(_00075_),
    .ZN(_15281_));
 AOI221_X4 _41954_ (.A(_07890_),
    .B1(_00599_),
    .B2(_15267_),
    .C1(_15280_),
    .C2(_15281_),
    .ZN(_15282_));
 OAI21_X1 _41955_ (.A(_08723_),
    .B1(_15266_),
    .B2(_15282_),
    .ZN(_15283_));
 NAND3_X1 _41956_ (.A1(_10739_),
    .A2(\icache.lce.lce_cmd_inst.state_r [1]),
    .A3(_07605_),
    .ZN(_15284_));
 NAND2_X1 _41957_ (.A1(_15283_),
    .A2(_15284_),
    .ZN(_05403_));
 NOR3_X1 _41958_ (.A1(_07604_),
    .A2(_07605_),
    .A3(lce_data_cmd_ready_i),
    .ZN(_15285_));
 AND2_X1 _41959_ (.A1(_15280_),
    .A2(_15281_),
    .ZN(_15286_));
 OAI21_X1 _41960_ (.A(_07896_),
    .B1(_08497_),
    .B2(_00598_),
    .ZN(_15287_));
 OAI221_X2 _41961_ (.A(_08662_),
    .B1(_07896_),
    .B2(_15285_),
    .C1(_15286_),
    .C2(_15287_),
    .ZN(_15288_));
 NAND2_X1 _41962_ (.A1(_15288_),
    .A2(_15284_),
    .ZN(_05404_));
 AOI21_X1 _41963_ (.A(_15262_),
    .B1(\icache.lce.lce_cmd_inst.syn_ack_cnt_r ),
    .B2(_15261_),
    .ZN(_15289_));
 AND2_X1 _41964_ (.A1(_00598_),
    .A2(_00599_),
    .ZN(_15290_));
 INV_X1 _41965_ (.A(_00600_),
    .ZN(_15291_));
 OAI211_X1 _41966_ (.A(_08674_),
    .B(_15290_),
    .C1(_15260_),
    .C2(_15291_),
    .ZN(_15292_));
 NAND2_X1 _41967_ (.A1(_08662_),
    .A2(\icache.lce.lce_cmd_inst.syn_ack_cnt_r ),
    .ZN(_15293_));
 OAI22_X1 _41968_ (.A1(_15289_),
    .A2(_15292_),
    .B1(_15290_),
    .B2(_15293_),
    .ZN(_05405_));
 AND3_X2 _41969_ (.A1(\icache.lce.lce_cmd_inst.state_r [1]),
    .A2(_00599_),
    .A3(lce_data_cmd_ready_i),
    .ZN(_15294_));
 INV_X32 _41970_ (.A(net1419),
    .ZN(_15295_));
 BUF_X32 _41971_ (.A(_15295_),
    .Z(_15296_));
 BUF_X32 _41972_ (.A(_15296_),
    .Z(_15297_));
 NAND2_X2 _41973_ (.A1(\icache.lce.lce_cmd_inst.state_r [1]),
    .A2(_00599_),
    .ZN(_15298_));
 AOI211_X1 _41974_ (.A(_11219_),
    .B(_15294_),
    .C1(_15297_),
    .C2(_15298_),
    .ZN(_05401_));
 NOR2_X1 _41975_ (.A1(_08516_),
    .A2(net1418),
    .ZN(_15299_));
 NAND2_X4 _41976_ (.A1(_07607_),
    .A2(_15299_),
    .ZN(_15300_));
 BUF_X8 _41977_ (.A(_15300_),
    .Z(_15301_));
 BUF_X16 _41978_ (.A(_15301_),
    .Z(_15302_));
 BUF_X8 _41979_ (.A(_15302_),
    .Z(_15303_));
 NAND2_X1 _41980_ (.A1(_15303_),
    .A2(\icache.lce.lce_cmd_inst.data_r [0]),
    .ZN(_15304_));
 INV_X8 _41981_ (.A(net1307),
    .ZN(_15305_));
 BUF_X16 _41982_ (.A(_15305_),
    .Z(_15306_));
 AND2_X1 _41983_ (.A1(_15306_),
    .A2(\icache.data_mems_6__data_mem.data_o [0]),
    .ZN(_15307_));
 BUF_X16 _41984_ (.A(net1310),
    .Z(_15308_));
 AND2_X1 _41985_ (.A1(_15308_),
    .A2(\icache.data_mems_7__data_mem.data_o [0]),
    .ZN(_15309_));
 INV_X8 _41986_ (.A(net1303),
    .ZN(_15310_));
 BUF_X16 _41987_ (.A(_15310_),
    .Z(_15311_));
 OR3_X1 _41988_ (.A1(_15307_),
    .A2(_15309_),
    .A3(_15311_),
    .ZN(_15312_));
 BUF_X16 _41989_ (.A(\icache.read_mux_butterfly.mux_stage_2__mux_swap_0__swap_inst.N0 ),
    .Z(_15313_));
 BUF_X16 _41990_ (.A(_15313_),
    .Z(_15314_));
 BUF_X8 _41991_ (.A(_15314_),
    .Z(_15315_));
 BUF_X16 _41992_ (.A(net1311),
    .Z(_15316_));
 BUF_X16 _41993_ (.A(_15316_),
    .Z(_15317_));
 BUF_X16 _41994_ (.A(_15317_),
    .Z(_15318_));
 NAND2_X1 _41995_ (.A1(_15318_),
    .A2(\icache.data_mems_5__data_mem.data_o [0]),
    .ZN(_15319_));
 BUF_X16 _41996_ (.A(_15310_),
    .Z(_15320_));
 BUF_X16 _41997_ (.A(_15320_),
    .Z(_15321_));
 BUF_X16 _41998_ (.A(net1312),
    .Z(_15322_));
 BUF_X16 _41999_ (.A(_15322_),
    .Z(_15323_));
 BUF_X16 _42000_ (.A(_15323_),
    .Z(_15324_));
 INV_X1 _42001_ (.A(\icache.data_mems_4__data_mem.data_o [0]),
    .ZN(_15325_));
 OAI211_X4 _42002_ (.A(_15319_),
    .B(_15321_),
    .C1(_15324_),
    .C2(_15325_),
    .ZN(_15326_));
 AND3_X1 _42003_ (.A1(_15312_),
    .A2(_15315_),
    .A3(_15326_),
    .ZN(_15327_));
 BUF_X16 _42004_ (.A(_15313_),
    .Z(_15328_));
 BUF_X16 _42005_ (.A(_15328_),
    .Z(_15329_));
 BUF_X16 _42006_ (.A(_15310_),
    .Z(_15330_));
 BUF_X16 _42007_ (.A(_15330_),
    .Z(_15331_));
 BUF_X16 _42008_ (.A(_15331_),
    .Z(_15332_));
 INV_X4 _42009_ (.A(\icache.data_mems_0__data_mem.data_o [0]),
    .ZN(_15333_));
 BUF_X16 _42010_ (.A(_15316_),
    .Z(_15334_));
 BUF_X8 _42011_ (.A(_15334_),
    .Z(_15335_));
 NOR2_X1 _42012_ (.A1(_15333_),
    .A2(_15335_),
    .ZN(_15336_));
 BUF_X16 _42013_ (.A(net1311),
    .Z(_15337_));
 BUF_X16 _42014_ (.A(_15337_),
    .Z(_15338_));
 AND2_X1 _42015_ (.A1(\icache.data_mems_1__data_mem.data_o [0]),
    .A2(_15338_),
    .ZN(_15339_));
 OAI21_X1 _42016_ (.A(_15332_),
    .B1(_15336_),
    .B2(_15339_),
    .ZN(_15340_));
 BUF_X16 _42017_ (.A(net1305),
    .Z(_15341_));
 BUF_X16 _42018_ (.A(_15341_),
    .Z(_15342_));
 BUF_X16 _42019_ (.A(_15342_),
    .Z(_15343_));
 INV_X1 _42020_ (.A(\icache.data_mems_2__data_mem.data_o [0]),
    .ZN(_15344_));
 NOR2_X1 _42021_ (.A1(_15344_),
    .A2(_15335_),
    .ZN(_15345_));
 BUF_X16 _42022_ (.A(_15337_),
    .Z(_15346_));
 AND2_X1 _42023_ (.A1(_15346_),
    .A2(\icache.data_mems_3__data_mem.data_o [0]),
    .ZN(_15347_));
 OAI21_X2 _42024_ (.A(_15343_),
    .B1(_15345_),
    .B2(_15347_),
    .ZN(_15348_));
 AOI21_X1 _42025_ (.A(_15329_),
    .B1(_15340_),
    .B2(_15348_),
    .ZN(_15349_));
 NOR2_X2 _42026_ (.A1(_15327_),
    .A2(_15349_),
    .ZN(_15350_));
 BUF_X16 _42027_ (.A(_15301_),
    .Z(_15351_));
 BUF_X8 _42028_ (.A(_15351_),
    .Z(_15352_));
 OAI21_X1 _42029_ (.A(_15304_),
    .B1(_15350_),
    .B2(_15352_),
    .ZN(_04889_));
 NAND2_X1 _42030_ (.A1(_15303_),
    .A2(\icache.lce.lce_cmd_inst.data_r [511]),
    .ZN(_15353_));
 BUF_X16 _42031_ (.A(_15328_),
    .Z(_15354_));
 AND2_X1 _42032_ (.A1(_15306_),
    .A2(\icache.data_mems_7__data_mem.data_o [63]),
    .ZN(_15355_));
 AND2_X1 _42033_ (.A1(_15308_),
    .A2(\icache.data_mems_6__data_mem.data_o [63]),
    .ZN(_15356_));
 OAI21_X2 _42034_ (.A(_15332_),
    .B1(_15355_),
    .B2(_15356_),
    .ZN(_15357_));
 INV_X1 _42035_ (.A(\icache.data_mems_5__data_mem.data_o [63]),
    .ZN(_15358_));
 BUF_X16 _42036_ (.A(_15316_),
    .Z(_15359_));
 NOR2_X1 _42037_ (.A1(_15358_),
    .A2(_15359_),
    .ZN(_15360_));
 BUF_X16 _42038_ (.A(net1308),
    .Z(_15361_));
 BUF_X16 _42039_ (.A(_15361_),
    .Z(_15362_));
 AND2_X1 _42040_ (.A1(_15362_),
    .A2(\icache.data_mems_4__data_mem.data_o [63]),
    .ZN(_15363_));
 OAI21_X2 _42041_ (.A(_15343_),
    .B1(_15360_),
    .B2(_15363_),
    .ZN(_15364_));
 AOI21_X2 _42042_ (.A(_15354_),
    .B1(_15357_),
    .B2(_15364_),
    .ZN(_15365_));
 INV_X16 _42043_ (.A(\icache.read_mux_butterfly.mux_stage_2__mux_swap_0__swap_inst.N0 ),
    .ZN(_15366_));
 BUF_X16 _42044_ (.A(_15366_),
    .Z(_15367_));
 BUF_X16 _42045_ (.A(_15367_),
    .Z(_15368_));
 BUF_X16 _42046_ (.A(_15341_),
    .Z(_15369_));
 BUF_X16 _42047_ (.A(_15369_),
    .Z(_15370_));
 BUF_X16 _42048_ (.A(_15305_),
    .Z(_15371_));
 BUF_X16 _42049_ (.A(_15371_),
    .Z(_15372_));
 AND2_X1 _42050_ (.A1(_15372_),
    .A2(\icache.data_mems_1__data_mem.data_o [63]),
    .ZN(_15373_));
 BUF_X16 _42051_ (.A(net1311),
    .Z(_15374_));
 BUF_X16 _42052_ (.A(_15374_),
    .Z(_15375_));
 AND2_X1 _42053_ (.A1(_15375_),
    .A2(\icache.data_mems_0__data_mem.data_o [63]),
    .ZN(_15376_));
 OAI21_X2 _42054_ (.A(_15370_),
    .B1(_15373_),
    .B2(_15376_),
    .ZN(_15377_));
 BUF_X16 _42055_ (.A(_15330_),
    .Z(_15378_));
 BUF_X16 _42056_ (.A(_15378_),
    .Z(_15379_));
 INV_X4 _42057_ (.A(\icache.data_mems_3__data_mem.data_o [63]),
    .ZN(_15380_));
 NOR2_X1 _42058_ (.A1(_15380_),
    .A2(_15335_),
    .ZN(_15381_));
 AND2_X1 _42059_ (.A1(_15346_),
    .A2(\icache.data_mems_2__data_mem.data_o [63]),
    .ZN(_15382_));
 OAI21_X2 _42060_ (.A(_15379_),
    .B1(_15381_),
    .B2(_15382_),
    .ZN(_15383_));
 AOI21_X2 _42061_ (.A(_15368_),
    .B1(_15377_),
    .B2(_15383_),
    .ZN(_15384_));
 NOR2_X4 _42062_ (.A1(_15365_),
    .A2(_15384_),
    .ZN(_15385_));
 OAI21_X1 _42063_ (.A(_15353_),
    .B1(_15385_),
    .B2(_15352_),
    .ZN(_05346_));
 NAND2_X1 _42064_ (.A1(_15303_),
    .A2(\icache.lce.lce_cmd_inst.data_r [510]),
    .ZN(_15386_));
 BUF_X8 _42065_ (.A(_15316_),
    .Z(_15387_));
 OR2_X1 _42066_ (.A1(_15387_),
    .A2(\icache.data_mems_7__data_mem.data_o [62]),
    .ZN(_15388_));
 INV_X2 _42067_ (.A(\icache.data_mems_6__data_mem.data_o [62]),
    .ZN(_15389_));
 BUF_X16 _42068_ (.A(_15361_),
    .Z(_15390_));
 BUF_X8 _42069_ (.A(_15390_),
    .Z(_15391_));
 NAND2_X1 _42070_ (.A1(_15389_),
    .A2(_15391_),
    .ZN(_15392_));
 NAND2_X1 _42071_ (.A1(_15388_),
    .A2(_15392_),
    .ZN(_15393_));
 BUF_X16 _42072_ (.A(_15330_),
    .Z(_15394_));
 BUF_X16 _42073_ (.A(_15394_),
    .Z(_15395_));
 NAND2_X1 _42074_ (.A1(_15393_),
    .A2(_15395_),
    .ZN(_15396_));
 BUF_X16 _42075_ (.A(_15305_),
    .Z(_15397_));
 BUF_X16 _42076_ (.A(_15397_),
    .Z(_15398_));
 INV_X4 _42077_ (.A(\icache.data_mems_5__data_mem.data_o [62]),
    .ZN(_15399_));
 NAND2_X1 _42078_ (.A1(_15398_),
    .A2(_15399_),
    .ZN(_15400_));
 INV_X2 _42079_ (.A(\icache.data_mems_4__data_mem.data_o [62]),
    .ZN(_15401_));
 BUF_X16 _42080_ (.A(_15362_),
    .Z(_15402_));
 NAND2_X1 _42081_ (.A1(_15401_),
    .A2(_15402_),
    .ZN(_15403_));
 NAND2_X1 _42082_ (.A1(_15400_),
    .A2(_15403_),
    .ZN(_15404_));
 BUF_X16 _42083_ (.A(_15341_),
    .Z(_15405_));
 BUF_X16 _42084_ (.A(_15405_),
    .Z(_15406_));
 NAND2_X1 _42085_ (.A1(_15404_),
    .A2(_15406_),
    .ZN(_15407_));
 BUF_X16 _42086_ (.A(_15366_),
    .Z(_15408_));
 BUF_X16 _42087_ (.A(_15408_),
    .Z(_15409_));
 NAND3_X1 _42088_ (.A1(_15396_),
    .A2(_15407_),
    .A3(_15409_),
    .ZN(_15410_));
 BUF_X8 _42089_ (.A(_15361_),
    .Z(_15411_));
 OR2_X1 _42090_ (.A1(_15411_),
    .A2(\icache.data_mems_1__data_mem.data_o [62]),
    .ZN(_15412_));
 INV_X8 _42091_ (.A(\icache.data_mems_0__data_mem.data_o [62]),
    .ZN(_15413_));
 NAND2_X1 _42092_ (.A1(_15413_),
    .A2(_15323_),
    .ZN(_15414_));
 NAND2_X1 _42093_ (.A1(_15412_),
    .A2(_15414_),
    .ZN(_15415_));
 NAND2_X1 _42094_ (.A1(_15415_),
    .A2(_15406_),
    .ZN(_15416_));
 BUF_X16 _42095_ (.A(_15371_),
    .Z(_15417_));
 INV_X8 _42096_ (.A(\icache.data_mems_3__data_mem.data_o [62]),
    .ZN(_15418_));
 NAND2_X1 _42097_ (.A1(_15417_),
    .A2(_15418_),
    .ZN(_15419_));
 INV_X4 _42098_ (.A(\icache.data_mems_2__data_mem.data_o [62]),
    .ZN(_15420_));
 BUF_X16 _42099_ (.A(_15374_),
    .Z(_15421_));
 NAND2_X1 _42100_ (.A1(_15420_),
    .A2(_15421_),
    .ZN(_15422_));
 NAND2_X1 _42101_ (.A1(_15419_),
    .A2(_15422_),
    .ZN(_15423_));
 BUF_X16 _42102_ (.A(_15310_),
    .Z(_15424_));
 BUF_X16 _42103_ (.A(_15424_),
    .Z(_15425_));
 NAND2_X1 _42104_ (.A1(_15423_),
    .A2(_15425_),
    .ZN(_15426_));
 NAND3_X1 _42105_ (.A1(_15416_),
    .A2(_15426_),
    .A3(_15315_),
    .ZN(_15427_));
 AND2_X2 _42106_ (.A1(_15410_),
    .A2(_15427_),
    .ZN(_15428_));
 OAI21_X1 _42107_ (.A(_15386_),
    .B1(_15428_),
    .B2(_15352_),
    .ZN(_05345_));
 NAND2_X1 _42108_ (.A1(_15303_),
    .A2(\icache.lce.lce_cmd_inst.data_r [509]),
    .ZN(_15429_));
 BUF_X16 _42109_ (.A(_15313_),
    .Z(_15430_));
 BUF_X16 _42110_ (.A(_15430_),
    .Z(_15431_));
 BUF_X16 _42111_ (.A(_15330_),
    .Z(_15432_));
 BUF_X16 _42112_ (.A(_15432_),
    .Z(_15433_));
 INV_X1 _42113_ (.A(\icache.data_mems_7__data_mem.data_o [61]),
    .ZN(_15434_));
 BUF_X16 _42114_ (.A(_15316_),
    .Z(_15435_));
 BUF_X16 _42115_ (.A(_15435_),
    .Z(_15436_));
 NOR2_X1 _42116_ (.A1(_15434_),
    .A2(_15436_),
    .ZN(_15437_));
 BUF_X16 _42117_ (.A(_15337_),
    .Z(_15438_));
 AND2_X1 _42118_ (.A1(_15438_),
    .A2(\icache.data_mems_6__data_mem.data_o [61]),
    .ZN(_15439_));
 OAI21_X2 _42119_ (.A(_15433_),
    .B1(_15437_),
    .B2(_15439_),
    .ZN(_15440_));
 OR2_X1 _42120_ (.A1(_15338_),
    .A2(\icache.data_mems_5__data_mem.data_o [61]),
    .ZN(_15441_));
 INV_X1 _42121_ (.A(\icache.data_mems_4__data_mem.data_o [61]),
    .ZN(_15442_));
 BUF_X16 _42122_ (.A(_15359_),
    .Z(_15443_));
 NAND2_X2 _42123_ (.A1(_15442_),
    .A2(_15443_),
    .ZN(_15444_));
 BUF_X16 _42124_ (.A(_15341_),
    .Z(_15445_));
 BUF_X16 _42125_ (.A(_15445_),
    .Z(_15446_));
 NAND3_X2 _42126_ (.A1(_15441_),
    .A2(_15444_),
    .A3(_15446_),
    .ZN(_15447_));
 AOI21_X2 _42127_ (.A(_15431_),
    .B1(_15440_),
    .B2(_15447_),
    .ZN(_15448_));
 BUF_X16 _42128_ (.A(_15367_),
    .Z(_15449_));
 BUF_X16 _42129_ (.A(_15331_),
    .Z(_15450_));
 INV_X4 _42130_ (.A(\icache.data_mems_3__data_mem.data_o [61]),
    .ZN(_15451_));
 BUF_X16 _42131_ (.A(_15435_),
    .Z(_15452_));
 NOR2_X1 _42132_ (.A1(_15451_),
    .A2(_15452_),
    .ZN(_15453_));
 BUF_X16 _42133_ (.A(_15374_),
    .Z(_15454_));
 AND2_X1 _42134_ (.A1(_15454_),
    .A2(\icache.data_mems_2__data_mem.data_o [61]),
    .ZN(_15455_));
 OAI21_X2 _42135_ (.A(_15450_),
    .B1(_15453_),
    .B2(_15455_),
    .ZN(_15456_));
 BUF_X16 _42136_ (.A(_15322_),
    .Z(_15457_));
 OR2_X1 _42137_ (.A1(_15457_),
    .A2(\icache.data_mems_1__data_mem.data_o [61]),
    .ZN(_15458_));
 INV_X4 _42138_ (.A(\icache.data_mems_0__data_mem.data_o [61]),
    .ZN(_15459_));
 BUF_X16 _42139_ (.A(_15316_),
    .Z(_15460_));
 BUF_X16 _42140_ (.A(_15460_),
    .Z(_15461_));
 NAND2_X2 _42141_ (.A1(_15459_),
    .A2(_15461_),
    .ZN(_15462_));
 BUF_X16 _42142_ (.A(_15341_),
    .Z(_15463_));
 BUF_X16 _42143_ (.A(_15463_),
    .Z(_15464_));
 NAND3_X2 _42144_ (.A1(_15458_),
    .A2(_15462_),
    .A3(_15464_),
    .ZN(_15465_));
 AOI21_X2 _42145_ (.A(_15449_),
    .B1(_15456_),
    .B2(_15465_),
    .ZN(_15466_));
 NOR2_X4 _42146_ (.A1(_15448_),
    .A2(_15466_),
    .ZN(_15467_));
 OAI21_X1 _42147_ (.A(_15429_),
    .B1(_15467_),
    .B2(_15352_),
    .ZN(_05343_));
 NAND2_X1 _42148_ (.A1(_15303_),
    .A2(\icache.lce.lce_cmd_inst.data_r [508]),
    .ZN(_15468_));
 INV_X1 _42149_ (.A(\icache.data_mems_1__data_mem.data_o [60]),
    .ZN(_15469_));
 NOR2_X1 _42150_ (.A1(_15469_),
    .A2(_15435_),
    .ZN(_15470_));
 BUF_X16 _42151_ (.A(net1313),
    .Z(_15471_));
 AND2_X1 _42152_ (.A1(_15471_),
    .A2(\icache.data_mems_0__data_mem.data_o [60]),
    .ZN(_15472_));
 OR3_X1 _42153_ (.A1(_15470_),
    .A2(_15472_),
    .A3(_15424_),
    .ZN(_15473_));
 BUF_X16 _42154_ (.A(_15314_),
    .Z(_15474_));
 BUF_X16 _42155_ (.A(_15308_),
    .Z(_15475_));
 NAND2_X1 _42156_ (.A1(_15475_),
    .A2(\icache.data_mems_2__data_mem.data_o [60]),
    .ZN(_15476_));
 BUF_X8 _42157_ (.A(_15320_),
    .Z(_15477_));
 BUF_X16 _42158_ (.A(_15337_),
    .Z(_15478_));
 BUF_X16 _42159_ (.A(_15478_),
    .Z(_15479_));
 INV_X1 _42160_ (.A(\icache.data_mems_3__data_mem.data_o [60]),
    .ZN(_15480_));
 OAI211_X2 _42161_ (.A(_15476_),
    .B(_15477_),
    .C1(_15479_),
    .C2(_15480_),
    .ZN(_15481_));
 AND3_X1 _42162_ (.A1(_15473_),
    .A2(_15474_),
    .A3(_15481_),
    .ZN(_15482_));
 BUF_X16 _42163_ (.A(net1306),
    .Z(_15483_));
 BUF_X16 _42164_ (.A(_15483_),
    .Z(_15484_));
 INV_X2 _42165_ (.A(\icache.data_mems_5__data_mem.data_o [60]),
    .ZN(_15485_));
 BUF_X8 _42166_ (.A(_15316_),
    .Z(_15486_));
 NOR2_X1 _42167_ (.A1(_15485_),
    .A2(_15486_),
    .ZN(_15487_));
 BUF_X8 _42168_ (.A(_15361_),
    .Z(_15488_));
 AND2_X1 _42169_ (.A1(_15488_),
    .A2(\icache.data_mems_4__data_mem.data_o [60]),
    .ZN(_15489_));
 OAI21_X1 _42170_ (.A(_15484_),
    .B1(_15487_),
    .B2(_15489_),
    .ZN(_15490_));
 BUF_X16 _42171_ (.A(_15371_),
    .Z(_15491_));
 INV_X8 _42172_ (.A(\icache.data_mems_7__data_mem.data_o [60]),
    .ZN(_15492_));
 NAND2_X1 _42173_ (.A1(_15491_),
    .A2(_15492_),
    .ZN(_15493_));
 INV_X4 _42174_ (.A(\icache.data_mems_6__data_mem.data_o [60]),
    .ZN(_15494_));
 BUF_X16 _42175_ (.A(_15337_),
    .Z(_15495_));
 NAND2_X1 _42176_ (.A1(_15494_),
    .A2(_15495_),
    .ZN(_15496_));
 BUF_X16 _42177_ (.A(_15330_),
    .Z(_15497_));
 NAND3_X1 _42178_ (.A1(_15493_),
    .A2(_15496_),
    .A3(_15497_),
    .ZN(_15498_));
 AOI21_X1 _42179_ (.A(_15329_),
    .B1(_15490_),
    .B2(_15498_),
    .ZN(_15499_));
 NOR2_X2 _42180_ (.A1(_15482_),
    .A2(_15499_),
    .ZN(_15500_));
 OAI21_X1 _42181_ (.A(_15468_),
    .B1(_15500_),
    .B2(_15352_),
    .ZN(_05342_));
 NAND2_X1 _42182_ (.A1(_15303_),
    .A2(\icache.lce.lce_cmd_inst.data_r [493]),
    .ZN(_15501_));
 BUF_X16 _42183_ (.A(_15366_),
    .Z(_15502_));
 BUF_X16 _42184_ (.A(_15502_),
    .Z(_15503_));
 INV_X8 _42185_ (.A(\icache.data_mems_1__data_mem.data_o [45]),
    .ZN(_15504_));
 BUF_X16 _42186_ (.A(_15316_),
    .Z(_15505_));
 NOR2_X1 _42187_ (.A1(_15504_),
    .A2(_15505_),
    .ZN(_15506_));
 AND2_X1 _42188_ (.A1(_15390_),
    .A2(\icache.data_mems_0__data_mem.data_o [45]),
    .ZN(_15507_));
 OR3_X1 _42189_ (.A1(_15506_),
    .A2(_15507_),
    .A3(_15424_),
    .ZN(_15508_));
 OR2_X1 _42190_ (.A1(_15411_),
    .A2(\icache.data_mems_3__data_mem.data_o [45]),
    .ZN(_15509_));
 INV_X4 _42191_ (.A(\icache.data_mems_2__data_mem.data_o [45]),
    .ZN(_15510_));
 BUF_X16 _42192_ (.A(_15362_),
    .Z(_15511_));
 NAND2_X1 _42193_ (.A1(_15510_),
    .A2(_15511_),
    .ZN(_15512_));
 NAND2_X1 _42194_ (.A1(_15509_),
    .A2(_15512_),
    .ZN(_15513_));
 BUF_X16 _42195_ (.A(_15311_),
    .Z(_15514_));
 NAND2_X1 _42196_ (.A1(_15513_),
    .A2(_15514_),
    .ZN(_15515_));
 AOI21_X1 _42197_ (.A(_15503_),
    .B1(_15508_),
    .B2(_15515_),
    .ZN(_15516_));
 INV_X1 _42198_ (.A(\icache.data_mems_5__data_mem.data_o [45]),
    .ZN(_15517_));
 BUF_X16 _42199_ (.A(_15337_),
    .Z(_15518_));
 NOR2_X1 _42200_ (.A1(_15517_),
    .A2(_15518_),
    .ZN(_15519_));
 AND2_X1 _42201_ (.A1(_15488_),
    .A2(\icache.data_mems_4__data_mem.data_o [45]),
    .ZN(_15520_));
 OAI21_X1 _42202_ (.A(_15484_),
    .B1(_15519_),
    .B2(_15520_),
    .ZN(_15521_));
 BUF_X16 _42203_ (.A(_15366_),
    .Z(_15522_));
 BUF_X16 _42204_ (.A(_15371_),
    .Z(_15523_));
 INV_X1 _42205_ (.A(\icache.data_mems_7__data_mem.data_o [45]),
    .ZN(_15524_));
 NAND2_X1 _42206_ (.A1(_15523_),
    .A2(_15524_),
    .ZN(_15525_));
 INV_X4 _42207_ (.A(\icache.data_mems_6__data_mem.data_o [45]),
    .ZN(_15526_));
 NAND2_X1 _42208_ (.A1(_15526_),
    .A2(_15495_),
    .ZN(_15527_));
 NAND3_X2 _42209_ (.A1(_15525_),
    .A2(_15527_),
    .A3(_15378_),
    .ZN(_15528_));
 AND3_X1 _42210_ (.A1(_15521_),
    .A2(_15522_),
    .A3(_15528_),
    .ZN(_15529_));
 OR2_X4 _42211_ (.A1(_15516_),
    .A2(_15529_),
    .ZN(_15530_));
 OAI21_X1 _42212_ (.A(_15501_),
    .B1(_15530_),
    .B2(_15352_),
    .ZN(_05325_));
 NAND2_X1 _42213_ (.A1(_15303_),
    .A2(\icache.lce.lce_cmd_inst.data_r [494]),
    .ZN(_15531_));
 INV_X8 _42214_ (.A(\icache.data_mems_1__data_mem.data_o [46]),
    .ZN(_15532_));
 BUF_X16 _42215_ (.A(_15316_),
    .Z(_15533_));
 NOR2_X1 _42216_ (.A1(_15532_),
    .A2(_15533_),
    .ZN(_15534_));
 AND2_X1 _42217_ (.A1(_15362_),
    .A2(\icache.data_mems_0__data_mem.data_o [46]),
    .ZN(_15535_));
 OR3_X1 _42218_ (.A1(_15534_),
    .A2(_15535_),
    .A3(_15311_),
    .ZN(_15536_));
 BUF_X16 _42219_ (.A(_15371_),
    .Z(_15537_));
 INV_X4 _42220_ (.A(\icache.data_mems_3__data_mem.data_o [46]),
    .ZN(_15538_));
 NAND2_X1 _42221_ (.A1(_15537_),
    .A2(_15538_),
    .ZN(_15539_));
 INV_X2 _42222_ (.A(\icache.data_mems_2__data_mem.data_o [46]),
    .ZN(_15540_));
 BUF_X16 _42223_ (.A(_15337_),
    .Z(_15541_));
 NAND2_X1 _42224_ (.A1(_15540_),
    .A2(_15541_),
    .ZN(_15542_));
 NAND2_X1 _42225_ (.A1(_15539_),
    .A2(_15542_),
    .ZN(_15543_));
 BUF_X16 _42226_ (.A(_15330_),
    .Z(_15544_));
 BUF_X16 _42227_ (.A(_15544_),
    .Z(_15545_));
 NAND2_X1 _42228_ (.A1(_15543_),
    .A2(_15545_),
    .ZN(_15546_));
 AND3_X1 _42229_ (.A1(_15536_),
    .A2(_15474_),
    .A3(_15546_),
    .ZN(_15547_));
 BUF_X16 _42230_ (.A(_15305_),
    .Z(_15548_));
 AND2_X1 _42231_ (.A1(_15548_),
    .A2(\icache.data_mems_7__data_mem.data_o [46]),
    .ZN(_15549_));
 BUF_X16 _42232_ (.A(_15361_),
    .Z(_15550_));
 AND2_X1 _42233_ (.A1(_15550_),
    .A2(\icache.data_mems_6__data_mem.data_o [46]),
    .ZN(_15551_));
 OAI21_X2 _42234_ (.A(_15332_),
    .B1(_15549_),
    .B2(_15551_),
    .ZN(_15552_));
 BUF_X16 _42235_ (.A(_15342_),
    .Z(_15553_));
 BUF_X8 _42236_ (.A(_15371_),
    .Z(_15554_));
 AND2_X1 _42237_ (.A1(_15554_),
    .A2(\icache.data_mems_5__data_mem.data_o [46]),
    .ZN(_15555_));
 BUF_X8 _42238_ (.A(_15361_),
    .Z(_15556_));
 AND2_X1 _42239_ (.A1(_15556_),
    .A2(\icache.data_mems_4__data_mem.data_o [46]),
    .ZN(_15557_));
 OAI21_X2 _42240_ (.A(_15553_),
    .B1(_15555_),
    .B2(_15557_),
    .ZN(_15558_));
 AOI21_X2 _42241_ (.A(_15329_),
    .B1(_15552_),
    .B2(_15558_),
    .ZN(_15559_));
 NOR2_X4 _42242_ (.A1(_15547_),
    .A2(_15559_),
    .ZN(_15560_));
 OAI21_X1 _42243_ (.A(_15531_),
    .B1(_15560_),
    .B2(_15352_),
    .ZN(_05326_));
 NAND2_X1 _42244_ (.A1(_15303_),
    .A2(\icache.lce.lce_cmd_inst.data_r [495]),
    .ZN(_15561_));
 OR2_X1 _42245_ (.A1(_15486_),
    .A2(\icache.data_mems_3__data_mem.data_o [47]),
    .ZN(_15562_));
 INV_X4 _42246_ (.A(\icache.data_mems_2__data_mem.data_o [47]),
    .ZN(_15563_));
 BUF_X16 _42247_ (.A(_15471_),
    .Z(_15564_));
 NAND2_X1 _42248_ (.A1(_15563_),
    .A2(_15564_),
    .ZN(_15565_));
 NAND2_X1 _42249_ (.A1(_15562_),
    .A2(_15565_),
    .ZN(_15566_));
 BUF_X16 _42250_ (.A(_15497_),
    .Z(_15567_));
 NAND2_X1 _42251_ (.A1(_15566_),
    .A2(_15567_),
    .ZN(_15568_));
 BUF_X16 _42252_ (.A(_15397_),
    .Z(_15569_));
 INV_X1 _42253_ (.A(\icache.data_mems_1__data_mem.data_o [47]),
    .ZN(_15570_));
 NAND2_X1 _42254_ (.A1(_15569_),
    .A2(_15570_),
    .ZN(_15571_));
 INV_X8 _42255_ (.A(\icache.data_mems_0__data_mem.data_o [47]),
    .ZN(_15572_));
 BUF_X16 _42256_ (.A(_15362_),
    .Z(_15573_));
 NAND2_X1 _42257_ (.A1(_15572_),
    .A2(_15573_),
    .ZN(_15574_));
 NAND2_X2 _42258_ (.A1(_15571_),
    .A2(_15574_),
    .ZN(_15575_));
 BUF_X16 _42259_ (.A(_15463_),
    .Z(_15576_));
 NAND2_X1 _42260_ (.A1(_15575_),
    .A2(_15576_),
    .ZN(_15577_));
 NAND2_X1 _42261_ (.A1(_15568_),
    .A2(_15577_),
    .ZN(_15578_));
 BUF_X16 _42262_ (.A(_15314_),
    .Z(_15579_));
 BUF_X16 _42263_ (.A(_15579_),
    .Z(_15580_));
 NAND2_X1 _42264_ (.A1(_15578_),
    .A2(_15580_),
    .ZN(_15581_));
 OR2_X1 _42265_ (.A1(_15486_),
    .A2(\icache.data_mems_5__data_mem.data_o [47]),
    .ZN(_15582_));
 INV_X2 _42266_ (.A(\icache.data_mems_4__data_mem.data_o [47]),
    .ZN(_15583_));
 NAND2_X1 _42267_ (.A1(_15583_),
    .A2(_15564_),
    .ZN(_15584_));
 NAND2_X1 _42268_ (.A1(_15582_),
    .A2(_15584_),
    .ZN(_15585_));
 BUF_X16 _42269_ (.A(_15341_),
    .Z(_15586_));
 BUF_X8 _42270_ (.A(_15586_),
    .Z(_15587_));
 NAND2_X1 _42271_ (.A1(_15585_),
    .A2(_15587_),
    .ZN(_15588_));
 INV_X1 _42272_ (.A(\icache.data_mems_7__data_mem.data_o [47]),
    .ZN(_15589_));
 NAND2_X1 _42273_ (.A1(_15569_),
    .A2(_15589_),
    .ZN(_15590_));
 INV_X1 _42274_ (.A(\icache.data_mems_6__data_mem.data_o [47]),
    .ZN(_15591_));
 NAND2_X1 _42275_ (.A1(_15591_),
    .A2(_15573_),
    .ZN(_15592_));
 NAND2_X2 _42276_ (.A1(_15590_),
    .A2(_15592_),
    .ZN(_15593_));
 BUF_X16 _42277_ (.A(_15378_),
    .Z(_15594_));
 NAND2_X1 _42278_ (.A1(_15593_),
    .A2(_15594_),
    .ZN(_15595_));
 NAND2_X1 _42279_ (.A1(_15588_),
    .A2(_15595_),
    .ZN(_15596_));
 BUF_X16 _42280_ (.A(_15502_),
    .Z(_15597_));
 BUF_X16 _42281_ (.A(_15597_),
    .Z(_15598_));
 NAND2_X1 _42282_ (.A1(_15596_),
    .A2(_15598_),
    .ZN(_15599_));
 NAND2_X2 _42283_ (.A1(_15581_),
    .A2(_15599_),
    .ZN(_15600_));
 OAI21_X1 _42284_ (.A(_15561_),
    .B1(_15600_),
    .B2(_15352_),
    .ZN(_05327_));
 BUF_X16 _42285_ (.A(_15301_),
    .Z(_15601_));
 BUF_X16 _42286_ (.A(_15601_),
    .Z(_15602_));
 NAND2_X1 _42287_ (.A1(_15602_),
    .A2(\icache.lce.lce_cmd_inst.data_r [496]),
    .ZN(_15603_));
 OR2_X1 _42288_ (.A1(_15435_),
    .A2(\icache.data_mems_1__data_mem.data_o [48]),
    .ZN(_15604_));
 INV_X8 _42289_ (.A(\icache.data_mems_0__data_mem.data_o [48]),
    .ZN(_15605_));
 BUF_X8 _42290_ (.A(_15374_),
    .Z(_15606_));
 NAND2_X2 _42291_ (.A1(_15605_),
    .A2(_15606_),
    .ZN(_15607_));
 NAND2_X1 _42292_ (.A1(_15604_),
    .A2(_15607_),
    .ZN(_15608_));
 BUF_X16 _42293_ (.A(_15341_),
    .Z(_15609_));
 BUF_X16 _42294_ (.A(_15609_),
    .Z(_15610_));
 NAND2_X1 _42295_ (.A1(_15608_),
    .A2(_15610_),
    .ZN(_15611_));
 BUF_X16 _42296_ (.A(_15397_),
    .Z(_15612_));
 INV_X8 _42297_ (.A(\icache.data_mems_3__data_mem.data_o [48]),
    .ZN(_15613_));
 NAND2_X1 _42298_ (.A1(_15612_),
    .A2(_15613_),
    .ZN(_15614_));
 INV_X4 _42299_ (.A(\icache.data_mems_2__data_mem.data_o [48]),
    .ZN(_15615_));
 BUF_X16 _42300_ (.A(_15374_),
    .Z(_15616_));
 NAND2_X1 _42301_ (.A1(_15615_),
    .A2(_15616_),
    .ZN(_15617_));
 NAND2_X1 _42302_ (.A1(_15614_),
    .A2(_15617_),
    .ZN(_15618_));
 BUF_X16 _42303_ (.A(_15544_),
    .Z(_15619_));
 NAND2_X1 _42304_ (.A1(_15618_),
    .A2(_15619_),
    .ZN(_15620_));
 BUF_X16 _42305_ (.A(_15314_),
    .Z(_15621_));
 AND3_X1 _42306_ (.A1(_15611_),
    .A2(_15620_),
    .A3(_15621_),
    .ZN(_15622_));
 INV_X8 _42307_ (.A(\icache.data_mems_7__data_mem.data_o [48]),
    .ZN(_15623_));
 NOR2_X2 _42308_ (.A1(_15623_),
    .A2(_15436_),
    .ZN(_15624_));
 AND2_X1 _42309_ (.A1(_15375_),
    .A2(\icache.data_mems_6__data_mem.data_o [48]),
    .ZN(_15625_));
 OAI21_X4 _42310_ (.A(_15332_),
    .B1(_15624_),
    .B2(_15625_),
    .ZN(_15626_));
 BUF_X16 _42311_ (.A(_15523_),
    .Z(_15627_));
 INV_X1 _42312_ (.A(\icache.data_mems_5__data_mem.data_o [48]),
    .ZN(_15628_));
 NAND2_X2 _42313_ (.A1(_15627_),
    .A2(_15628_),
    .ZN(_15629_));
 INV_X2 _42314_ (.A(\icache.data_mems_4__data_mem.data_o [48]),
    .ZN(_15630_));
 NAND2_X2 _42315_ (.A1(_15630_),
    .A2(_15461_),
    .ZN(_15631_));
 NAND3_X4 _42316_ (.A1(_15629_),
    .A2(_15631_),
    .A3(_15576_),
    .ZN(_15632_));
 AOI21_X2 _42317_ (.A(_15329_),
    .B1(_15626_),
    .B2(_15632_),
    .ZN(_15633_));
 NOR2_X4 _42318_ (.A1(_15622_),
    .A2(_15633_),
    .ZN(_15634_));
 OAI21_X1 _42319_ (.A(_15603_),
    .B1(_15634_),
    .B2(_15352_),
    .ZN(_05328_));
 NAND2_X1 _42320_ (.A1(_15602_),
    .A2(\icache.lce.lce_cmd_inst.data_r [497]),
    .ZN(_15635_));
 BUF_X16 _42321_ (.A(_15371_),
    .Z(_15636_));
 AND2_X1 _42322_ (.A1(_15636_),
    .A2(\icache.data_mems_3__data_mem.data_o [49]),
    .ZN(_15637_));
 AND2_X1 _42323_ (.A1(_15564_),
    .A2(\icache.data_mems_2__data_mem.data_o [49]),
    .ZN(_15638_));
 OAI21_X2 _42324_ (.A(_15433_),
    .B1(_15637_),
    .B2(_15638_),
    .ZN(_15639_));
 INV_X4 _42325_ (.A(\icache.data_mems_1__data_mem.data_o [49]),
    .ZN(_15640_));
 NOR2_X1 _42326_ (.A1(_15640_),
    .A2(_15436_),
    .ZN(_15641_));
 AND2_X1 _42327_ (.A1(_15375_),
    .A2(\icache.data_mems_0__data_mem.data_o [49]),
    .ZN(_15642_));
 OAI21_X2 _42328_ (.A(_15370_),
    .B1(_15641_),
    .B2(_15642_),
    .ZN(_15643_));
 BUF_X16 _42329_ (.A(_15313_),
    .Z(_15644_));
 BUF_X16 _42330_ (.A(_15644_),
    .Z(_15645_));
 NAND3_X2 _42331_ (.A1(_15639_),
    .A2(_15643_),
    .A3(_15645_),
    .ZN(_15646_));
 AND2_X1 _42332_ (.A1(_15372_),
    .A2(\icache.data_mems_7__data_mem.data_o [49]),
    .ZN(_15647_));
 AND2_X1 _42333_ (.A1(_15454_),
    .A2(\icache.data_mems_6__data_mem.data_o [49]),
    .ZN(_15648_));
 OAI21_X2 _42334_ (.A(_15450_),
    .B1(_15647_),
    .B2(_15648_),
    .ZN(_15649_));
 BUF_X16 _42335_ (.A(_15463_),
    .Z(_15650_));
 INV_X1 _42336_ (.A(\icache.data_mems_5__data_mem.data_o [49]),
    .ZN(_15651_));
 NOR2_X2 _42337_ (.A1(_15651_),
    .A2(_15318_),
    .ZN(_15652_));
 AND2_X1 _42338_ (.A1(_15438_),
    .A2(\icache.data_mems_4__data_mem.data_o [49]),
    .ZN(_15653_));
 OAI21_X2 _42339_ (.A(_15650_),
    .B1(_15652_),
    .B2(_15653_),
    .ZN(_15654_));
 BUF_X16 _42340_ (.A(_15366_),
    .Z(_15655_));
 BUF_X32 _42341_ (.A(_15655_),
    .Z(_15656_));
 NAND3_X2 _42342_ (.A1(_15649_),
    .A2(_15654_),
    .A3(_15656_),
    .ZN(_15657_));
 NAND2_X4 _42343_ (.A1(_15646_),
    .A2(_15657_),
    .ZN(_15658_));
 OAI21_X1 _42344_ (.A(_15635_),
    .B1(_15658_),
    .B2(_15352_),
    .ZN(_05329_));
 NAND2_X1 _42345_ (.A1(_15602_),
    .A2(\icache.lce.lce_cmd_inst.data_r [498]),
    .ZN(_15659_));
 BUF_X16 _42346_ (.A(_15483_),
    .Z(_15660_));
 AND2_X1 _42347_ (.A1(_15554_),
    .A2(\icache.data_mems_5__data_mem.data_o [50]),
    .ZN(_15661_));
 AND2_X1 _42348_ (.A1(_15556_),
    .A2(\icache.data_mems_4__data_mem.data_o [50]),
    .ZN(_15662_));
 OAI21_X1 _42349_ (.A(_15660_),
    .B1(_15661_),
    .B2(_15662_),
    .ZN(_15663_));
 BUF_X16 _42350_ (.A(_15320_),
    .Z(_15664_));
 INV_X4 _42351_ (.A(\icache.data_mems_7__data_mem.data_o [50]),
    .ZN(_15665_));
 NOR2_X1 _42352_ (.A1(_15665_),
    .A2(_15486_),
    .ZN(_15666_));
 AND2_X1 _42353_ (.A1(_15488_),
    .A2(\icache.data_mems_6__data_mem.data_o [50]),
    .ZN(_15667_));
 OAI21_X1 _42354_ (.A(_15664_),
    .B1(_15666_),
    .B2(_15667_),
    .ZN(_15668_));
 AND3_X1 _42355_ (.A1(_15663_),
    .A2(_15655_),
    .A3(_15668_),
    .ZN(_15669_));
 BUF_X8 _42356_ (.A(_15502_),
    .Z(_15670_));
 BUF_X16 _42357_ (.A(_15397_),
    .Z(_15671_));
 NAND2_X1 _42358_ (.A1(_15671_),
    .A2(\icache.data_mems_1__data_mem.data_o [50]),
    .ZN(_15672_));
 BUF_X16 _42359_ (.A(_15483_),
    .Z(_15673_));
 BUF_X16 _42360_ (.A(_15417_),
    .Z(_15674_));
 INV_X8 _42361_ (.A(\icache.data_mems_0__data_mem.data_o [50]),
    .ZN(_15675_));
 OAI211_X4 _42362_ (.A(_15672_),
    .B(_15673_),
    .C1(_15674_),
    .C2(_15675_),
    .ZN(_15676_));
 NAND2_X1 _42363_ (.A1(_15569_),
    .A2(\icache.data_mems_3__data_mem.data_o [50]),
    .ZN(_15677_));
 BUF_X16 _42364_ (.A(_15320_),
    .Z(_15678_));
 BUF_X8 _42365_ (.A(_15523_),
    .Z(_15679_));
 INV_X4 _42366_ (.A(\icache.data_mems_2__data_mem.data_o [50]),
    .ZN(_15680_));
 OAI211_X2 _42367_ (.A(_15677_),
    .B(_15678_),
    .C1(_15679_),
    .C2(_15680_),
    .ZN(_15681_));
 AOI21_X2 _42368_ (.A(_15670_),
    .B1(_15676_),
    .B2(_15681_),
    .ZN(_15682_));
 OR2_X4 _42369_ (.A1(_15669_),
    .A2(_15682_),
    .ZN(_15683_));
 BUF_X16 _42370_ (.A(_15351_),
    .Z(_15684_));
 OAI21_X1 _42371_ (.A(_15659_),
    .B1(_15683_),
    .B2(_15684_),
    .ZN(_05330_));
 NAND2_X1 _42372_ (.A1(_15602_),
    .A2(\icache.lce.lce_cmd_inst.data_r [499]),
    .ZN(_15685_));
 BUF_X16 _42373_ (.A(_15313_),
    .Z(_15686_));
 INV_X1 _42374_ (.A(\icache.data_mems_5__data_mem.data_o [51]),
    .ZN(_15687_));
 NOR2_X1 _42375_ (.A1(_15687_),
    .A2(_15435_),
    .ZN(_15688_));
 AND2_X1 _42376_ (.A1(_15471_),
    .A2(\icache.data_mems_4__data_mem.data_o [51]),
    .ZN(_15689_));
 OR3_X1 _42377_ (.A1(_15688_),
    .A2(_15689_),
    .A3(_15424_),
    .ZN(_15690_));
 NAND2_X1 _42378_ (.A1(_15636_),
    .A2(\icache.data_mems_7__data_mem.data_o [51]),
    .ZN(_15691_));
 BUF_X16 _42379_ (.A(_15523_),
    .Z(_15692_));
 INV_X2 _42380_ (.A(\icache.data_mems_6__data_mem.data_o [51]),
    .ZN(_15693_));
 OAI211_X4 _42381_ (.A(_15691_),
    .B(_15477_),
    .C1(_15692_),
    .C2(_15693_),
    .ZN(_15694_));
 AOI21_X1 _42382_ (.A(_15686_),
    .B1(_15690_),
    .B2(_15694_),
    .ZN(_15695_));
 AND2_X1 _42383_ (.A1(_15548_),
    .A2(\icache.data_mems_3__data_mem.data_o [51]),
    .ZN(_15696_));
 AND2_X1 _42384_ (.A1(_15488_),
    .A2(\icache.data_mems_2__data_mem.data_o [51]),
    .ZN(_15697_));
 OAI21_X2 _42385_ (.A(_15664_),
    .B1(_15696_),
    .B2(_15697_),
    .ZN(_15698_));
 BUF_X16 _42386_ (.A(_15313_),
    .Z(_15699_));
 BUF_X16 _42387_ (.A(_15361_),
    .Z(_15700_));
 OR2_X2 _42388_ (.A1(_15700_),
    .A2(\icache.data_mems_1__data_mem.data_o [51]),
    .ZN(_15701_));
 INV_X8 _42389_ (.A(\icache.data_mems_0__data_mem.data_o [51]),
    .ZN(_15702_));
 NAND2_X2 _42390_ (.A1(_15702_),
    .A2(_15495_),
    .ZN(_15703_));
 NAND3_X4 _42391_ (.A1(_15701_),
    .A2(_15703_),
    .A3(_15586_),
    .ZN(_15704_));
 AND3_X1 _42392_ (.A1(_15698_),
    .A2(_15699_),
    .A3(_15704_),
    .ZN(_15705_));
 OR2_X2 _42393_ (.A1(_15695_),
    .A2(_15705_),
    .ZN(_15706_));
 OAI21_X1 _42394_ (.A(_15685_),
    .B1(_15706_),
    .B2(_15684_),
    .ZN(_05331_));
 NAND2_X1 _42395_ (.A1(_15602_),
    .A2(\icache.lce.lce_cmd_inst.data_r [500]),
    .ZN(_15707_));
 BUF_X16 _42396_ (.A(_15432_),
    .Z(_15708_));
 AND2_X1 _42397_ (.A1(_15306_),
    .A2(\icache.data_mems_7__data_mem.data_o [52]),
    .ZN(_15709_));
 AND2_X1 _42398_ (.A1(_15471_),
    .A2(\icache.data_mems_6__data_mem.data_o [52]),
    .ZN(_15710_));
 OAI21_X2 _42399_ (.A(_15708_),
    .B1(_15709_),
    .B2(_15710_),
    .ZN(_15711_));
 BUF_X16 _42400_ (.A(_15369_),
    .Z(_15712_));
 INV_X1 _42401_ (.A(\icache.data_mems_5__data_mem.data_o [52]),
    .ZN(_15713_));
 BUF_X16 _42402_ (.A(_15316_),
    .Z(_15714_));
 NOR2_X1 _42403_ (.A1(_15713_),
    .A2(_15714_),
    .ZN(_15715_));
 AND2_X1 _42404_ (.A1(_15362_),
    .A2(\icache.data_mems_4__data_mem.data_o [52]),
    .ZN(_15716_));
 OAI21_X2 _42405_ (.A(_15712_),
    .B1(_15715_),
    .B2(_15716_),
    .ZN(_15717_));
 AOI21_X2 _42406_ (.A(_15431_),
    .B1(_15711_),
    .B2(_15717_),
    .ZN(_15718_));
 BUF_X8 _42407_ (.A(_15548_),
    .Z(_15719_));
 NAND2_X1 _42408_ (.A1(_15719_),
    .A2(\icache.data_mems_3__data_mem.data_o [52]),
    .ZN(_15720_));
 BUF_X16 _42409_ (.A(_15417_),
    .Z(_15721_));
 INV_X8 _42410_ (.A(\icache.data_mems_2__data_mem.data_o [52]),
    .ZN(_15722_));
 OAI211_X1 _42411_ (.A(_15720_),
    .B(_15321_),
    .C1(_15721_),
    .C2(_15722_),
    .ZN(_15723_));
 BUF_X16 _42412_ (.A(_15313_),
    .Z(_15724_));
 BUF_X16 _42413_ (.A(_15550_),
    .Z(_15725_));
 NAND2_X1 _42414_ (.A1(_15725_),
    .A2(\icache.data_mems_0__data_mem.data_o [52]),
    .ZN(_15726_));
 BUF_X8 _42415_ (.A(_15483_),
    .Z(_15727_));
 BUF_X8 _42416_ (.A(_15478_),
    .Z(_15728_));
 INV_X1 _42417_ (.A(\icache.data_mems_1__data_mem.data_o [52]),
    .ZN(_15729_));
 OAI211_X2 _42418_ (.A(_15726_),
    .B(_15727_),
    .C1(_15728_),
    .C2(_15729_),
    .ZN(_15730_));
 AND3_X1 _42419_ (.A1(_15723_),
    .A2(_15724_),
    .A3(_15730_),
    .ZN(_15731_));
 NOR2_X4 _42420_ (.A1(_15718_),
    .A2(_15731_),
    .ZN(_15732_));
 OAI21_X1 _42421_ (.A(_15707_),
    .B1(_15732_),
    .B2(_15684_),
    .ZN(_05334_));
 NAND2_X1 _42422_ (.A1(_15602_),
    .A2(\icache.lce.lce_cmd_inst.data_r [501]),
    .ZN(_15733_));
 BUF_X16 _42423_ (.A(_15313_),
    .Z(_15734_));
 BUF_X16 _42424_ (.A(_15734_),
    .Z(_15735_));
 BUF_X16 _42425_ (.A(_15371_),
    .Z(_15736_));
 AND2_X1 _42426_ (.A1(_15736_),
    .A2(\icache.data_mems_1__data_mem.data_o [53]),
    .ZN(_15737_));
 BUF_X16 _42427_ (.A(_15374_),
    .Z(_15738_));
 AND2_X1 _42428_ (.A1(_15738_),
    .A2(\icache.data_mems_0__data_mem.data_o [53]),
    .ZN(_15739_));
 BUF_X16 _42429_ (.A(_15544_),
    .Z(_15740_));
 NOR3_X2 _42430_ (.A1(_15737_),
    .A2(_15739_),
    .A3(_15740_),
    .ZN(_15741_));
 OR2_X1 _42431_ (.A1(_15457_),
    .A2(\icache.data_mems_3__data_mem.data_o [53]),
    .ZN(_15742_));
 INV_X8 _42432_ (.A(\icache.data_mems_2__data_mem.data_o [53]),
    .ZN(_15743_));
 NAND2_X1 _42433_ (.A1(_15743_),
    .A2(_15461_),
    .ZN(_15744_));
 AOI21_X2 _42434_ (.A(_15610_),
    .B1(_15742_),
    .B2(_15744_),
    .ZN(_15745_));
 OAI21_X2 _42435_ (.A(_15735_),
    .B1(_15741_),
    .B2(_15745_),
    .ZN(_15746_));
 BUF_X16 _42436_ (.A(_15523_),
    .Z(_15747_));
 INV_X1 _42437_ (.A(\icache.data_mems_7__data_mem.data_o [53]),
    .ZN(_15748_));
 NAND2_X2 _42438_ (.A1(_15747_),
    .A2(_15748_),
    .ZN(_15749_));
 INV_X2 _42439_ (.A(\icache.data_mems_6__data_mem.data_o [53]),
    .ZN(_15750_));
 BUF_X16 _42440_ (.A(_15337_),
    .Z(_15751_));
 BUF_X16 _42441_ (.A(_15751_),
    .Z(_15752_));
 NAND2_X2 _42442_ (.A1(_15750_),
    .A2(_15752_),
    .ZN(_15753_));
 BUF_X16 _42443_ (.A(_15432_),
    .Z(_15754_));
 NAND3_X2 _42444_ (.A1(_15749_),
    .A2(_15753_),
    .A3(_15754_),
    .ZN(_15755_));
 BUF_X16 _42445_ (.A(_15554_),
    .Z(_15756_));
 INV_X1 _42446_ (.A(\icache.data_mems_5__data_mem.data_o [53]),
    .ZN(_15757_));
 NAND2_X1 _42447_ (.A1(_15756_),
    .A2(_15757_),
    .ZN(_15758_));
 INV_X2 _42448_ (.A(\icache.data_mems_4__data_mem.data_o [53]),
    .ZN(_15759_));
 NAND2_X1 _42449_ (.A1(_15759_),
    .A2(_15443_),
    .ZN(_15760_));
 BUF_X16 _42450_ (.A(_15660_),
    .Z(_15761_));
 NAND3_X2 _42451_ (.A1(_15758_),
    .A2(_15760_),
    .A3(_15761_),
    .ZN(_15762_));
 NAND3_X2 _42452_ (.A1(_15755_),
    .A2(_15762_),
    .A3(_15656_),
    .ZN(_15763_));
 NAND2_X4 _42453_ (.A1(_15746_),
    .A2(_15763_),
    .ZN(_15764_));
 OAI21_X1 _42454_ (.A(_15733_),
    .B1(_15764_),
    .B2(_15684_),
    .ZN(_05335_));
 NAND2_X1 _42455_ (.A1(_15602_),
    .A2(\icache.lce.lce_cmd_inst.data_r [502]),
    .ZN(_15765_));
 OR2_X1 _42456_ (.A1(_15387_),
    .A2(\icache.data_mems_5__data_mem.data_o [54]),
    .ZN(_15766_));
 INV_X2 _42457_ (.A(\icache.data_mems_4__data_mem.data_o [54]),
    .ZN(_15767_));
 NAND2_X1 _42458_ (.A1(_15767_),
    .A2(_15391_),
    .ZN(_15768_));
 NAND2_X1 _42459_ (.A1(_15766_),
    .A2(_15768_),
    .ZN(_15769_));
 BUF_X16 _42460_ (.A(_15609_),
    .Z(_15770_));
 NAND2_X1 _42461_ (.A1(_15769_),
    .A2(_15770_),
    .ZN(_15771_));
 BUF_X16 _42462_ (.A(_15397_),
    .Z(_15772_));
 INV_X4 _42463_ (.A(\icache.data_mems_7__data_mem.data_o [54]),
    .ZN(_15773_));
 NAND2_X1 _42464_ (.A1(_15772_),
    .A2(_15773_),
    .ZN(_15774_));
 INV_X4 _42465_ (.A(\icache.data_mems_6__data_mem.data_o [54]),
    .ZN(_15775_));
 BUF_X16 _42466_ (.A(_15374_),
    .Z(_15776_));
 NAND2_X1 _42467_ (.A1(_15775_),
    .A2(_15776_),
    .ZN(_15777_));
 NAND2_X2 _42468_ (.A1(_15774_),
    .A2(_15777_),
    .ZN(_15778_));
 BUF_X16 _42469_ (.A(_15544_),
    .Z(_15779_));
 NAND2_X1 _42470_ (.A1(_15778_),
    .A2(_15779_),
    .ZN(_15780_));
 AOI21_X1 _42471_ (.A(_15686_),
    .B1(_15771_),
    .B2(_15780_),
    .ZN(_15781_));
 INV_X4 _42472_ (.A(\icache.data_mems_3__data_mem.data_o [54]),
    .ZN(_15782_));
 NOR2_X1 _42473_ (.A1(_15782_),
    .A2(_15533_),
    .ZN(_15783_));
 BUF_X8 _42474_ (.A(_15361_),
    .Z(_15784_));
 AND2_X1 _42475_ (.A1(_15784_),
    .A2(\icache.data_mems_2__data_mem.data_o [54]),
    .ZN(_15785_));
 OAI21_X1 _42476_ (.A(_15664_),
    .B1(_15783_),
    .B2(_15785_),
    .ZN(_15786_));
 INV_X1 _42477_ (.A(\icache.data_mems_1__data_mem.data_o [54]),
    .ZN(_15787_));
 NOR2_X1 _42478_ (.A1(_15787_),
    .A2(_15533_),
    .ZN(_15788_));
 AND2_X1 _42479_ (.A1(_15784_),
    .A2(\icache.data_mems_0__data_mem.data_o [54]),
    .ZN(_15789_));
 OAI21_X2 _42480_ (.A(_15445_),
    .B1(_15788_),
    .B2(_15789_),
    .ZN(_15790_));
 AND3_X1 _42481_ (.A1(_15786_),
    .A2(_15790_),
    .A3(_15328_),
    .ZN(_15791_));
 OR2_X2 _42482_ (.A1(_15781_),
    .A2(_15791_),
    .ZN(_15792_));
 OAI21_X1 _42483_ (.A(_15765_),
    .B1(_15792_),
    .B2(_15684_),
    .ZN(_05336_));
 NAND2_X1 _42484_ (.A1(_15602_),
    .A2(\icache.lce.lce_cmd_inst.data_r [503]),
    .ZN(_15793_));
 OR2_X1 _42485_ (.A1(_15387_),
    .A2(\icache.data_mems_1__data_mem.data_o [55]),
    .ZN(_15794_));
 INV_X8 _42486_ (.A(\icache.data_mems_0__data_mem.data_o [55]),
    .ZN(_15795_));
 NAND2_X1 _42487_ (.A1(_15795_),
    .A2(_15391_),
    .ZN(_15796_));
 NAND2_X1 _42488_ (.A1(_15794_),
    .A2(_15796_),
    .ZN(_15797_));
 NAND2_X1 _42489_ (.A1(_15797_),
    .A2(_15770_),
    .ZN(_15798_));
 INV_X4 _42490_ (.A(\icache.data_mems_3__data_mem.data_o [55]),
    .ZN(_15799_));
 NAND2_X1 _42491_ (.A1(_15772_),
    .A2(_15799_),
    .ZN(_15800_));
 INV_X8 _42492_ (.A(\icache.data_mems_2__data_mem.data_o [55]),
    .ZN(_15801_));
 NAND2_X1 _42493_ (.A1(_15801_),
    .A2(_15776_),
    .ZN(_15802_));
 NAND2_X1 _42494_ (.A1(_15800_),
    .A2(_15802_),
    .ZN(_15803_));
 BUF_X16 _42495_ (.A(_15311_),
    .Z(_15804_));
 NAND2_X1 _42496_ (.A1(_15803_),
    .A2(_15804_),
    .ZN(_15805_));
 AOI21_X1 _42497_ (.A(_15503_),
    .B1(_15798_),
    .B2(_15805_),
    .ZN(_15806_));
 INV_X4 _42498_ (.A(\icache.data_mems_7__data_mem.data_o [55]),
    .ZN(_15807_));
 NAND2_X1 _42499_ (.A1(_15537_),
    .A2(_15807_),
    .ZN(_15808_));
 INV_X4 _42500_ (.A(\icache.data_mems_6__data_mem.data_o [55]),
    .ZN(_15809_));
 BUF_X16 _42501_ (.A(_15374_),
    .Z(_15810_));
 NAND2_X1 _42502_ (.A1(_15809_),
    .A2(_15810_),
    .ZN(_15811_));
 BUF_X16 _42503_ (.A(_15330_),
    .Z(_15812_));
 NAND3_X1 _42504_ (.A1(_15808_),
    .A2(_15811_),
    .A3(_15812_),
    .ZN(_15813_));
 INV_X2 _42505_ (.A(\icache.data_mems_5__data_mem.data_o [55]),
    .ZN(_15814_));
 NAND2_X1 _42506_ (.A1(_15491_),
    .A2(_15814_),
    .ZN(_15815_));
 INV_X2 _42507_ (.A(\icache.data_mems_4__data_mem.data_o [55]),
    .ZN(_15816_));
 NAND2_X1 _42508_ (.A1(_15816_),
    .A2(_15478_),
    .ZN(_15817_));
 NAND3_X1 _42509_ (.A1(_15815_),
    .A2(_15817_),
    .A3(_15586_),
    .ZN(_15818_));
 BUF_X16 _42510_ (.A(_15366_),
    .Z(_15819_));
 AND3_X1 _42511_ (.A1(_15813_),
    .A2(_15818_),
    .A3(_15819_),
    .ZN(_15820_));
 OR2_X2 _42512_ (.A1(_15806_),
    .A2(_15820_),
    .ZN(_15821_));
 OAI21_X1 _42513_ (.A(_15793_),
    .B1(_15821_),
    .B2(_15684_),
    .ZN(_05337_));
 NAND2_X1 _42514_ (.A1(_15602_),
    .A2(\icache.lce.lce_cmd_inst.data_r [504]),
    .ZN(_15822_));
 OR2_X1 _42515_ (.A1(_15387_),
    .A2(\icache.data_mems_1__data_mem.data_o [56]),
    .ZN(_15823_));
 INV_X8 _42516_ (.A(\icache.data_mems_0__data_mem.data_o [56]),
    .ZN(_15824_));
 NAND2_X1 _42517_ (.A1(_15824_),
    .A2(_15391_),
    .ZN(_15825_));
 NAND2_X1 _42518_ (.A1(_15823_),
    .A2(_15825_),
    .ZN(_15826_));
 NAND2_X1 _42519_ (.A1(_15826_),
    .A2(_15770_),
    .ZN(_15827_));
 OR2_X1 _42520_ (.A1(_15317_),
    .A2(\icache.data_mems_3__data_mem.data_o [56]),
    .ZN(_15828_));
 INV_X8 _42521_ (.A(\icache.data_mems_2__data_mem.data_o [56]),
    .ZN(_15829_));
 NAND2_X1 _42522_ (.A1(_15829_),
    .A2(_15402_),
    .ZN(_15830_));
 NAND2_X1 _42523_ (.A1(_15828_),
    .A2(_15830_),
    .ZN(_15831_));
 NAND2_X1 _42524_ (.A1(_15831_),
    .A2(_15804_),
    .ZN(_15832_));
 BUF_X16 _42525_ (.A(_15313_),
    .Z(_15833_));
 BUF_X16 _42526_ (.A(_15833_),
    .Z(_15834_));
 NAND3_X1 _42527_ (.A1(_15827_),
    .A2(_15832_),
    .A3(_15834_),
    .ZN(_15835_));
 BUF_X16 _42528_ (.A(_15397_),
    .Z(_15836_));
 INV_X1 _42529_ (.A(\icache.data_mems_5__data_mem.data_o [56]),
    .ZN(_15837_));
 NAND2_X1 _42530_ (.A1(_15836_),
    .A2(_15837_),
    .ZN(_15838_));
 INV_X1 _42531_ (.A(\icache.data_mems_4__data_mem.data_o [56]),
    .ZN(_15839_));
 NAND2_X1 _42532_ (.A1(_15839_),
    .A2(_15323_),
    .ZN(_15840_));
 NAND2_X1 _42533_ (.A1(_15838_),
    .A2(_15840_),
    .ZN(_15841_));
 NAND2_X1 _42534_ (.A1(_15841_),
    .A2(_15406_),
    .ZN(_15842_));
 INV_X1 _42535_ (.A(\icache.data_mems_7__data_mem.data_o [56]),
    .ZN(_15843_));
 NAND2_X1 _42536_ (.A1(_15417_),
    .A2(_15843_),
    .ZN(_15844_));
 INV_X1 _42537_ (.A(\icache.data_mems_6__data_mem.data_o [56]),
    .ZN(_15845_));
 NAND2_X1 _42538_ (.A1(_15845_),
    .A2(_15421_),
    .ZN(_15846_));
 NAND2_X1 _42539_ (.A1(_15844_),
    .A2(_15846_),
    .ZN(_15847_));
 NAND2_X1 _42540_ (.A1(_15847_),
    .A2(_15425_),
    .ZN(_15848_));
 BUF_X16 _42541_ (.A(_15408_),
    .Z(_15849_));
 NAND3_X1 _42542_ (.A1(_15842_),
    .A2(_15848_),
    .A3(_15849_),
    .ZN(_15850_));
 AND2_X4 _42543_ (.A1(_15835_),
    .A2(_15850_),
    .ZN(_15851_));
 OAI21_X1 _42544_ (.A(_15822_),
    .B1(_15851_),
    .B2(_15684_),
    .ZN(_05338_));
 NAND2_X1 _42545_ (.A1(_15602_),
    .A2(\icache.lce.lce_cmd_inst.data_r [505]),
    .ZN(_15852_));
 BUF_X16 _42546_ (.A(_15660_),
    .Z(_15853_));
 AND2_X1 _42547_ (.A1(_15372_),
    .A2(\icache.data_mems_5__data_mem.data_o [57]),
    .ZN(_15854_));
 AND2_X1 _42548_ (.A1(_15438_),
    .A2(\icache.data_mems_4__data_mem.data_o [57]),
    .ZN(_15855_));
 OAI21_X2 _42549_ (.A(_15853_),
    .B1(_15854_),
    .B2(_15855_),
    .ZN(_15856_));
 OR2_X1 _42550_ (.A1(_15338_),
    .A2(\icache.data_mems_7__data_mem.data_o [57]),
    .ZN(_15857_));
 INV_X2 _42551_ (.A(\icache.data_mems_6__data_mem.data_o [57]),
    .ZN(_15858_));
 NAND2_X1 _42552_ (.A1(_15858_),
    .A2(_15443_),
    .ZN(_15859_));
 BUF_X16 _42553_ (.A(_15331_),
    .Z(_15860_));
 NAND3_X2 _42554_ (.A1(_15857_),
    .A2(_15859_),
    .A3(_15860_),
    .ZN(_15861_));
 AOI21_X2 _42555_ (.A(_15431_),
    .B1(_15856_),
    .B2(_15861_),
    .ZN(_15862_));
 INV_X4 _42556_ (.A(\icache.data_mems_3__data_mem.data_o [57]),
    .ZN(_15863_));
 NOR2_X1 _42557_ (.A1(_15863_),
    .A2(_15318_),
    .ZN(_15864_));
 AND2_X1 _42558_ (.A1(_15616_),
    .A2(\icache.data_mems_2__data_mem.data_o [57]),
    .ZN(_15865_));
 OAI21_X2 _42559_ (.A(_15332_),
    .B1(_15864_),
    .B2(_15865_),
    .ZN(_15866_));
 INV_X1 _42560_ (.A(\icache.data_mems_1__data_mem.data_o [57]),
    .ZN(_15867_));
 NOR2_X1 _42561_ (.A1(_15867_),
    .A2(_15335_),
    .ZN(_15868_));
 AND2_X1 _42562_ (.A1(_15346_),
    .A2(\icache.data_mems_0__data_mem.data_o [57]),
    .ZN(_15869_));
 OAI21_X2 _42563_ (.A(_15553_),
    .B1(_15868_),
    .B2(_15869_),
    .ZN(_15870_));
 AOI21_X2 _42564_ (.A(_15449_),
    .B1(_15866_),
    .B2(_15870_),
    .ZN(_15871_));
 NOR2_X4 _42565_ (.A1(_15862_),
    .A2(_15871_),
    .ZN(_15872_));
 OAI21_X1 _42566_ (.A(_15852_),
    .B1(_15872_),
    .B2(_15684_),
    .ZN(_05339_));
 BUF_X4 _42567_ (.A(_15601_),
    .Z(_15873_));
 NAND2_X1 _42568_ (.A1(_15873_),
    .A2(\icache.lce.lce_cmd_inst.data_r [506]),
    .ZN(_15874_));
 AND2_X1 _42569_ (.A1(_15554_),
    .A2(\icache.data_mems_3__data_mem.data_o [58]),
    .ZN(_15875_));
 BUF_X16 _42570_ (.A(_15361_),
    .Z(_15876_));
 AND2_X1 _42571_ (.A1(_15876_),
    .A2(\icache.data_mems_2__data_mem.data_o [58]),
    .ZN(_15877_));
 OR3_X1 _42572_ (.A1(_15875_),
    .A2(_15877_),
    .A3(_15609_),
    .ZN(_15878_));
 INV_X1 _42573_ (.A(\icache.data_mems_1__data_mem.data_o [58]),
    .ZN(_15879_));
 NOR2_X2 _42574_ (.A1(_15879_),
    .A2(_15751_),
    .ZN(_15880_));
 AND2_X1 _42575_ (.A1(_15700_),
    .A2(\icache.data_mems_0__data_mem.data_o [58]),
    .ZN(_15881_));
 OR3_X1 _42576_ (.A1(_15880_),
    .A2(_15881_),
    .A3(_15544_),
    .ZN(_15882_));
 NAND2_X1 _42577_ (.A1(_15878_),
    .A2(_15882_),
    .ZN(_15883_));
 NAND2_X1 _42578_ (.A1(_15883_),
    .A2(_15580_),
    .ZN(_15884_));
 INV_X1 _42579_ (.A(\icache.data_mems_5__data_mem.data_o [58]),
    .ZN(_15885_));
 NAND2_X1 _42580_ (.A1(_15612_),
    .A2(_15885_),
    .ZN(_15886_));
 INV_X1 _42581_ (.A(\icache.data_mems_4__data_mem.data_o [58]),
    .ZN(_15887_));
 NAND2_X1 _42582_ (.A1(_15887_),
    .A2(_15616_),
    .ZN(_15888_));
 NAND2_X1 _42583_ (.A1(_15886_),
    .A2(_15888_),
    .ZN(_15889_));
 NAND2_X1 _42584_ (.A1(_15889_),
    .A2(_15587_),
    .ZN(_15890_));
 INV_X4 _42585_ (.A(\icache.data_mems_7__data_mem.data_o [58]),
    .ZN(_15891_));
 NAND2_X1 _42586_ (.A1(_15736_),
    .A2(_15891_),
    .ZN(_15892_));
 INV_X1 _42587_ (.A(\icache.data_mems_6__data_mem.data_o [58]),
    .ZN(_15893_));
 NAND2_X1 _42588_ (.A1(_15893_),
    .A2(_15606_),
    .ZN(_15894_));
 NAND2_X1 _42589_ (.A1(_15892_),
    .A2(_15894_),
    .ZN(_15895_));
 NAND2_X1 _42590_ (.A1(_15895_),
    .A2(_15594_),
    .ZN(_15896_));
 NAND2_X1 _42591_ (.A1(_15890_),
    .A2(_15896_),
    .ZN(_15897_));
 NAND2_X2 _42592_ (.A1(_15897_),
    .A2(_15598_),
    .ZN(_15898_));
 NAND2_X4 _42593_ (.A1(_15884_),
    .A2(_15898_),
    .ZN(_15899_));
 OAI21_X1 _42594_ (.A(_15874_),
    .B1(_15899_),
    .B2(_15684_),
    .ZN(_05340_));
 NAND2_X1 _42595_ (.A1(_15873_),
    .A2(\icache.lce.lce_cmd_inst.data_r [413]),
    .ZN(_15900_));
 BUF_X16 _42596_ (.A(_15660_),
    .Z(_15901_));
 AND2_X1 _42597_ (.A1(_15636_),
    .A2(\icache.data_mems_4__data_mem.data_o [29]),
    .ZN(_15902_));
 AND2_X1 _42598_ (.A1(_15457_),
    .A2(\icache.data_mems_5__data_mem.data_o [29]),
    .ZN(_15903_));
 OAI21_X1 _42599_ (.A(_15901_),
    .B1(_15902_),
    .B2(_15903_),
    .ZN(_15904_));
 BUF_X16 _42600_ (.A(_15597_),
    .Z(_15905_));
 BUF_X16 _42601_ (.A(_15362_),
    .Z(_15906_));
 OR2_X1 _42602_ (.A1(_15906_),
    .A2(\icache.data_mems_6__data_mem.data_o [29]),
    .ZN(_15907_));
 INV_X2 _42603_ (.A(\icache.data_mems_7__data_mem.data_o [29]),
    .ZN(_15908_));
 BUF_X16 _42604_ (.A(_15751_),
    .Z(_15909_));
 NAND2_X1 _42605_ (.A1(_15908_),
    .A2(_15909_),
    .ZN(_15910_));
 BUF_X16 _42606_ (.A(_15497_),
    .Z(_15911_));
 NAND3_X2 _42607_ (.A1(_15907_),
    .A2(_15910_),
    .A3(_15911_),
    .ZN(_15912_));
 NAND3_X1 _42608_ (.A1(_15904_),
    .A2(_15905_),
    .A3(_15912_),
    .ZN(_15913_));
 INV_X8 _42609_ (.A(\icache.data_mems_2__data_mem.data_o [29]),
    .ZN(_15914_));
 NOR2_X2 _42610_ (.A1(_15914_),
    .A2(_15443_),
    .ZN(_15915_));
 BUF_X16 _42611_ (.A(_15374_),
    .Z(_15916_));
 AND2_X2 _42612_ (.A1(_15916_),
    .A2(\icache.data_mems_3__data_mem.data_o [29]),
    .ZN(_15917_));
 OAI21_X4 _42613_ (.A(_15450_),
    .B1(_15915_),
    .B2(_15917_),
    .ZN(_15918_));
 INV_X8 _42614_ (.A(\icache.data_mems_0__data_mem.data_o [29]),
    .ZN(_15919_));
 NAND2_X2 _42615_ (.A1(_15679_),
    .A2(_15919_),
    .ZN(_15920_));
 INV_X1 _42616_ (.A(\icache.data_mems_1__data_mem.data_o [29]),
    .ZN(_15921_));
 BUF_X16 _42617_ (.A(_15460_),
    .Z(_15922_));
 NAND2_X2 _42618_ (.A1(_15921_),
    .A2(_15922_),
    .ZN(_15923_));
 NAND3_X2 _42619_ (.A1(_15920_),
    .A2(_15923_),
    .A3(_15464_),
    .ZN(_15924_));
 NAND3_X2 _42620_ (.A1(_15918_),
    .A2(_15645_),
    .A3(_15924_),
    .ZN(_15925_));
 NAND2_X4 _42621_ (.A1(_15913_),
    .A2(_15925_),
    .ZN(_15926_));
 OAI21_X1 _42622_ (.A(_15900_),
    .B1(_15926_),
    .B2(_15684_),
    .ZN(_05237_));
 NAND2_X1 _42623_ (.A1(_15873_),
    .A2(\icache.lce.lce_cmd_inst.data_r [414]),
    .ZN(_15927_));
 OR2_X1 _42624_ (.A1(_15334_),
    .A2(\icache.data_mems_4__data_mem.data_o [30]),
    .ZN(_15928_));
 INV_X1 _42625_ (.A(\icache.data_mems_5__data_mem.data_o [30]),
    .ZN(_15929_));
 NAND2_X1 _42626_ (.A1(_15929_),
    .A2(_15776_),
    .ZN(_15930_));
 NAND2_X1 _42627_ (.A1(_15928_),
    .A2(_15930_),
    .ZN(_15931_));
 BUF_X16 _42628_ (.A(_15405_),
    .Z(_15932_));
 NAND2_X1 _42629_ (.A1(_15931_),
    .A2(_15932_),
    .ZN(_15933_));
 OR2_X1 _42630_ (.A1(_15556_),
    .A2(\icache.data_mems_6__data_mem.data_o [30]),
    .ZN(_15934_));
 INV_X8 _42631_ (.A(\icache.data_mems_7__data_mem.data_o [30]),
    .ZN(_15935_));
 NAND2_X1 _42632_ (.A1(_15935_),
    .A2(_15541_),
    .ZN(_15936_));
 NAND2_X1 _42633_ (.A1(_15934_),
    .A2(_15936_),
    .ZN(_15937_));
 BUF_X16 _42634_ (.A(_15311_),
    .Z(_15938_));
 NAND2_X1 _42635_ (.A1(_15937_),
    .A2(_15938_),
    .ZN(_15939_));
 BUF_X16 _42636_ (.A(_15502_),
    .Z(_15940_));
 AND3_X1 _42637_ (.A1(_15933_),
    .A2(_15939_),
    .A3(_15940_),
    .ZN(_15941_));
 AND2_X1 _42638_ (.A1(_15548_),
    .A2(\icache.data_mems_2__data_mem.data_o [30]),
    .ZN(_15942_));
 AND2_X1 _42639_ (.A1(_15556_),
    .A2(\icache.data_mems_3__data_mem.data_o [30]),
    .ZN(_15943_));
 OAI21_X2 _42640_ (.A(_15678_),
    .B1(_15942_),
    .B2(_15943_),
    .ZN(_15944_));
 OR2_X1 _42641_ (.A1(_15556_),
    .A2(\icache.data_mems_0__data_mem.data_o [30]),
    .ZN(_15945_));
 INV_X4 _42642_ (.A(\icache.data_mems_1__data_mem.data_o [30]),
    .ZN(_15946_));
 NAND2_X1 _42643_ (.A1(_15946_),
    .A2(_15810_),
    .ZN(_15947_));
 NAND3_X1 _42644_ (.A1(_15945_),
    .A2(_15947_),
    .A3(_15484_),
    .ZN(_15948_));
 AOI21_X2 _42645_ (.A(_15449_),
    .B1(_15944_),
    .B2(_15948_),
    .ZN(_15949_));
 NOR2_X4 _42646_ (.A1(_15941_),
    .A2(_15949_),
    .ZN(_15950_));
 BUF_X8 _42647_ (.A(_15351_),
    .Z(_15951_));
 OAI21_X1 _42648_ (.A(_15927_),
    .B1(_15950_),
    .B2(_15951_),
    .ZN(_05238_));
 NAND2_X1 _42649_ (.A1(_15873_),
    .A2(\icache.lce.lce_cmd_inst.data_r [415]),
    .ZN(_15952_));
 OR2_X1 _42650_ (.A1(_15334_),
    .A2(\icache.data_mems_4__data_mem.data_o [31]),
    .ZN(_15953_));
 INV_X1 _42651_ (.A(\icache.data_mems_5__data_mem.data_o [31]),
    .ZN(_15954_));
 BUF_X16 _42652_ (.A(_15362_),
    .Z(_15955_));
 NAND2_X1 _42653_ (.A1(_15954_),
    .A2(_15955_),
    .ZN(_15956_));
 NAND3_X1 _42654_ (.A1(_15953_),
    .A2(_15956_),
    .A3(_15660_),
    .ZN(_15957_));
 INV_X8 _42655_ (.A(\icache.data_mems_6__data_mem.data_o [31]),
    .ZN(_15958_));
 NAND2_X1 _42656_ (.A1(_15836_),
    .A2(_15958_),
    .ZN(_15959_));
 INV_X8 _42657_ (.A(\icache.data_mems_7__data_mem.data_o [31]),
    .ZN(_15960_));
 NAND2_X1 _42658_ (.A1(_15960_),
    .A2(_15810_),
    .ZN(_15961_));
 NAND3_X1 _42659_ (.A1(_15959_),
    .A2(_15961_),
    .A3(_15664_),
    .ZN(_15962_));
 AND3_X1 _42660_ (.A1(_15957_),
    .A2(_15962_),
    .A3(_15522_),
    .ZN(_15963_));
 NAND2_X1 _42661_ (.A1(_15671_),
    .A2(\icache.data_mems_0__data_mem.data_o [31]),
    .ZN(_15964_));
 INV_X4 _42662_ (.A(\icache.data_mems_1__data_mem.data_o [31]),
    .ZN(_15965_));
 OAI211_X2 _42663_ (.A(_15964_),
    .B(_15673_),
    .C1(_15674_),
    .C2(_15965_),
    .ZN(_15966_));
 BUF_X16 _42664_ (.A(_15784_),
    .Z(_15967_));
 NAND2_X1 _42665_ (.A1(_15967_),
    .A2(\icache.data_mems_3__data_mem.data_o [31]),
    .ZN(_15968_));
 INV_X1 _42666_ (.A(\icache.data_mems_2__data_mem.data_o [31]),
    .ZN(_15969_));
 OAI211_X1 _42667_ (.A(_15968_),
    .B(_15678_),
    .C1(_15728_),
    .C2(_15969_),
    .ZN(_15970_));
 AOI21_X1 _42668_ (.A(_15670_),
    .B1(_15966_),
    .B2(_15970_),
    .ZN(_15971_));
 OR2_X4 _42669_ (.A1(_15963_),
    .A2(_15971_),
    .ZN(_15972_));
 OAI21_X1 _42670_ (.A(_15952_),
    .B1(_15972_),
    .B2(_15951_),
    .ZN(_05239_));
 NAND2_X1 _42671_ (.A1(_15873_),
    .A2(\icache.lce.lce_cmd_inst.data_r [416]),
    .ZN(_15973_));
 AND2_X1 _42672_ (.A1(_15636_),
    .A2(\icache.data_mems_6__data_mem.data_o [32]),
    .ZN(_15974_));
 AND2_X1 _42673_ (.A1(_15457_),
    .A2(\icache.data_mems_7__data_mem.data_o [32]),
    .ZN(_15975_));
 OAI21_X2 _42674_ (.A(_15433_),
    .B1(_15974_),
    .B2(_15975_),
    .ZN(_15976_));
 OR2_X1 _42675_ (.A1(_15906_),
    .A2(\icache.data_mems_4__data_mem.data_o [32]),
    .ZN(_15977_));
 INV_X1 _42676_ (.A(\icache.data_mems_5__data_mem.data_o [32]),
    .ZN(_15978_));
 NAND2_X2 _42677_ (.A1(_15978_),
    .A2(_15909_),
    .ZN(_15979_));
 NAND3_X2 _42678_ (.A1(_15977_),
    .A2(_15979_),
    .A3(_15446_),
    .ZN(_15980_));
 NAND3_X2 _42679_ (.A1(_15976_),
    .A2(_15905_),
    .A3(_15980_),
    .ZN(_15981_));
 INV_X8 _42680_ (.A(\icache.data_mems_2__data_mem.data_o [32]),
    .ZN(_15982_));
 NAND2_X4 _42681_ (.A1(_15674_),
    .A2(_15982_),
    .ZN(_15983_));
 INV_X2 _42682_ (.A(\icache.data_mems_3__data_mem.data_o [32]),
    .ZN(_15984_));
 BUF_X16 _42683_ (.A(_15337_),
    .Z(_15985_));
 BUF_X16 _42684_ (.A(_15985_),
    .Z(_15986_));
 NAND2_X1 _42685_ (.A1(_15984_),
    .A2(_15986_),
    .ZN(_15987_));
 BUF_X16 _42686_ (.A(_15497_),
    .Z(_15988_));
 NAND3_X2 _42687_ (.A1(_15983_),
    .A2(_15987_),
    .A3(_15988_),
    .ZN(_15989_));
 INV_X8 _42688_ (.A(\icache.data_mems_0__data_mem.data_o [32]),
    .ZN(_15990_));
 NAND2_X2 _42689_ (.A1(_15679_),
    .A2(_15990_),
    .ZN(_15991_));
 INV_X1 _42690_ (.A(\icache.data_mems_1__data_mem.data_o [32]),
    .ZN(_15992_));
 NAND2_X2 _42691_ (.A1(_15992_),
    .A2(_15922_),
    .ZN(_15993_));
 BUF_X16 _42692_ (.A(_15463_),
    .Z(_15994_));
 NAND3_X4 _42693_ (.A1(_15991_),
    .A2(_15993_),
    .A3(_15994_),
    .ZN(_15995_));
 BUF_X16 _42694_ (.A(_15644_),
    .Z(_15996_));
 NAND3_X2 _42695_ (.A1(_15989_),
    .A2(_15995_),
    .A3(_15996_),
    .ZN(_15997_));
 NAND2_X4 _42696_ (.A1(_15981_),
    .A2(_15997_),
    .ZN(_15998_));
 OAI21_X1 _42697_ (.A(_15973_),
    .B1(_15998_),
    .B2(_15951_),
    .ZN(_05240_));
 NAND2_X1 _42698_ (.A1(_15873_),
    .A2(\icache.lce.lce_cmd_inst.data_r [417]),
    .ZN(_15999_));
 INV_X8 _42699_ (.A(\icache.data_mems_0__data_mem.data_o [33]),
    .ZN(_16000_));
 BUF_X16 _42700_ (.A(_15505_),
    .Z(_16001_));
 NOR2_X4 _42701_ (.A1(_16000_),
    .A2(_16001_),
    .ZN(_16002_));
 AND2_X1 _42702_ (.A1(_15457_),
    .A2(\icache.data_mems_1__data_mem.data_o [33]),
    .ZN(_16003_));
 NOR3_X2 _42703_ (.A1(_16002_),
    .A2(_16003_),
    .A3(_15740_),
    .ZN(_16004_));
 BUF_X16 _42704_ (.A(_15609_),
    .Z(_16005_));
 OR2_X1 _42705_ (.A1(_15906_),
    .A2(\icache.data_mems_2__data_mem.data_o [33]),
    .ZN(_16006_));
 INV_X8 _42706_ (.A(\icache.data_mems_3__data_mem.data_o [33]),
    .ZN(_16007_));
 BUF_X16 _42707_ (.A(_15751_),
    .Z(_16008_));
 NAND2_X4 _42708_ (.A1(_16007_),
    .A2(_16008_),
    .ZN(_16009_));
 AOI21_X2 _42709_ (.A(_16005_),
    .B1(_16006_),
    .B2(_16009_),
    .ZN(_16010_));
 OAI21_X2 _42710_ (.A(_15735_),
    .B1(_16004_),
    .B2(_16010_),
    .ZN(_16011_));
 BUF_X16 _42711_ (.A(_15366_),
    .Z(_16012_));
 BUF_X16 _42712_ (.A(_16012_),
    .Z(_16013_));
 BUF_X16 _42713_ (.A(_15378_),
    .Z(_16014_));
 BUF_X16 _42714_ (.A(_15322_),
    .Z(_16015_));
 OR2_X1 _42715_ (.A1(_16015_),
    .A2(\icache.data_mems_4__data_mem.data_o [33]),
    .ZN(_16016_));
 INV_X1 _42716_ (.A(\icache.data_mems_5__data_mem.data_o [33]),
    .ZN(_16017_));
 BUF_X16 _42717_ (.A(_15478_),
    .Z(_16018_));
 NAND2_X2 _42718_ (.A1(_16017_),
    .A2(_16018_),
    .ZN(_16019_));
 AOI21_X2 _42719_ (.A(_16014_),
    .B1(_16016_),
    .B2(_16019_),
    .ZN(_16020_));
 BUF_X16 _42720_ (.A(_15609_),
    .Z(_16021_));
 INV_X8 _42721_ (.A(\icache.data_mems_6__data_mem.data_o [33]),
    .ZN(_16022_));
 NAND2_X2 _42722_ (.A1(_15679_),
    .A2(_16022_),
    .ZN(_16023_));
 INV_X1 _42723_ (.A(\icache.data_mems_7__data_mem.data_o [33]),
    .ZN(_16024_));
 NAND2_X2 _42724_ (.A1(_16024_),
    .A2(_15922_),
    .ZN(_16025_));
 AOI21_X4 _42725_ (.A(_16021_),
    .B1(_16023_),
    .B2(_16025_),
    .ZN(_16026_));
 OAI21_X2 _42726_ (.A(_16013_),
    .B1(_16020_),
    .B2(_16026_),
    .ZN(_16027_));
 NAND2_X4 _42727_ (.A1(_16011_),
    .A2(_16027_),
    .ZN(_16028_));
 OAI21_X1 _42728_ (.A(_15999_),
    .B1(_16028_),
    .B2(_15951_),
    .ZN(_05241_));
 NAND2_X1 _42729_ (.A1(_15873_),
    .A2(\icache.lce.lce_cmd_inst.data_r [418]),
    .ZN(_16029_));
 AND2_X1 _42730_ (.A1(_15306_),
    .A2(\icache.data_mems_4__data_mem.data_o [34]),
    .ZN(_16030_));
 AND2_X1 _42731_ (.A1(_15308_),
    .A2(\icache.data_mems_5__data_mem.data_o [34]),
    .ZN(_16031_));
 OR3_X1 _42732_ (.A1(_16030_),
    .A2(_16031_),
    .A3(_15311_),
    .ZN(_16032_));
 BUF_X8 _42733_ (.A(_15502_),
    .Z(_16033_));
 NAND2_X1 _42734_ (.A1(_15719_),
    .A2(\icache.data_mems_6__data_mem.data_o [34]),
    .ZN(_16034_));
 BUF_X16 _42735_ (.A(_15417_),
    .Z(_16035_));
 INV_X8 _42736_ (.A(\icache.data_mems_7__data_mem.data_o [34]),
    .ZN(_16036_));
 OAI211_X2 _42737_ (.A(_16034_),
    .B(_15321_),
    .C1(_16035_),
    .C2(_16036_),
    .ZN(_16037_));
 AND3_X2 _42738_ (.A1(_16032_),
    .A2(_16033_),
    .A3(_16037_),
    .ZN(_16038_));
 AND2_X1 _42739_ (.A1(_15372_),
    .A2(\icache.data_mems_0__data_mem.data_o [34]),
    .ZN(_16039_));
 AND2_X1 _42740_ (.A1(_15375_),
    .A2(\icache.data_mems_1__data_mem.data_o [34]),
    .ZN(_16040_));
 OAI21_X2 _42741_ (.A(_15370_),
    .B1(_16039_),
    .B2(_16040_),
    .ZN(_16041_));
 INV_X8 _42742_ (.A(\icache.data_mems_2__data_mem.data_o [34]),
    .ZN(_16042_));
 NOR2_X1 _42743_ (.A1(_16042_),
    .A2(_15335_),
    .ZN(_16043_));
 AND2_X1 _42744_ (.A1(_15346_),
    .A2(\icache.data_mems_3__data_mem.data_o [34]),
    .ZN(_16044_));
 OAI21_X2 _42745_ (.A(_15379_),
    .B1(_16043_),
    .B2(_16044_),
    .ZN(_16045_));
 AOI21_X2 _42746_ (.A(_15449_),
    .B1(_16041_),
    .B2(_16045_),
    .ZN(_16046_));
 NOR2_X4 _42747_ (.A1(_16038_),
    .A2(_16046_),
    .ZN(_16047_));
 OAI21_X1 _42748_ (.A(_16029_),
    .B1(_16047_),
    .B2(_15951_),
    .ZN(_05242_));
 NAND2_X1 _42749_ (.A1(_15873_),
    .A2(\icache.lce.lce_cmd_inst.data_r [419]),
    .ZN(_16048_));
 BUF_X16 _42750_ (.A(_15502_),
    .Z(_16049_));
 INV_X8 _42751_ (.A(\icache.data_mems_2__data_mem.data_o [35]),
    .ZN(_16050_));
 NOR2_X4 _42752_ (.A1(_16050_),
    .A2(_15435_),
    .ZN(_16051_));
 AND2_X1 _42753_ (.A1(_15471_),
    .A2(\icache.data_mems_3__data_mem.data_o [35]),
    .ZN(_16052_));
 BUF_X16 _42754_ (.A(_15341_),
    .Z(_16053_));
 OR3_X1 _42755_ (.A1(_16051_),
    .A2(_16052_),
    .A3(_16053_),
    .ZN(_16054_));
 NAND2_X1 _42756_ (.A1(_15636_),
    .A2(\icache.data_mems_0__data_mem.data_o [35]),
    .ZN(_16055_));
 BUF_X8 _42757_ (.A(_15483_),
    .Z(_16056_));
 INV_X1 _42758_ (.A(\icache.data_mems_1__data_mem.data_o [35]),
    .ZN(_16057_));
 OAI211_X2 _42759_ (.A(_16055_),
    .B(_16056_),
    .C1(_15692_),
    .C2(_16057_),
    .ZN(_16058_));
 AOI21_X1 _42760_ (.A(_16049_),
    .B1(_16054_),
    .B2(_16058_),
    .ZN(_16059_));
 AND2_X1 _42761_ (.A1(_15306_),
    .A2(\icache.data_mems_6__data_mem.data_o [35]),
    .ZN(_16060_));
 BUF_X16 _42762_ (.A(_15361_),
    .Z(_16061_));
 AND2_X1 _42763_ (.A1(_16061_),
    .A2(\icache.data_mems_7__data_mem.data_o [35]),
    .ZN(_16062_));
 OAI21_X1 _42764_ (.A(_15664_),
    .B1(_16060_),
    .B2(_16062_),
    .ZN(_16063_));
 INV_X2 _42765_ (.A(\icache.data_mems_4__data_mem.data_o [35]),
    .ZN(_16064_));
 NAND2_X2 _42766_ (.A1(_15491_),
    .A2(_16064_),
    .ZN(_16065_));
 INV_X1 _42767_ (.A(\icache.data_mems_5__data_mem.data_o [35]),
    .ZN(_16066_));
 BUF_X16 _42768_ (.A(_15337_),
    .Z(_16067_));
 NAND2_X2 _42769_ (.A1(_16066_),
    .A2(_16067_),
    .ZN(_16068_));
 NAND3_X1 _42770_ (.A1(_16065_),
    .A2(_16068_),
    .A3(_15586_),
    .ZN(_16069_));
 AND3_X1 _42771_ (.A1(_16063_),
    .A2(_15522_),
    .A3(_16069_),
    .ZN(_16070_));
 OR2_X4 _42772_ (.A1(_16059_),
    .A2(_16070_),
    .ZN(_16071_));
 OAI21_X1 _42773_ (.A(_16048_),
    .B1(_16071_),
    .B2(_15951_),
    .ZN(_05243_));
 NAND2_X1 _42774_ (.A1(_15873_),
    .A2(\icache.lce.lce_cmd_inst.data_r [420]),
    .ZN(_16072_));
 OR2_X2 _42775_ (.A1(_15475_),
    .A2(\icache.data_mems_0__data_mem.data_o [36]),
    .ZN(_16073_));
 INV_X2 _42776_ (.A(\icache.data_mems_1__data_mem.data_o [36]),
    .ZN(_16074_));
 NAND2_X2 _42777_ (.A1(_16074_),
    .A2(_15479_),
    .ZN(_16075_));
 NAND3_X2 _42778_ (.A1(_16073_),
    .A2(_16075_),
    .A3(_15712_),
    .ZN(_16076_));
 INV_X1 _42779_ (.A(\icache.data_mems_2__data_mem.data_o [36]),
    .ZN(_16077_));
 NAND2_X2 _42780_ (.A1(_16035_),
    .A2(_16077_),
    .ZN(_16078_));
 INV_X1 _42781_ (.A(\icache.data_mems_3__data_mem.data_o [36]),
    .ZN(_16079_));
 NAND2_X2 _42782_ (.A1(_16079_),
    .A2(_15728_),
    .ZN(_16080_));
 NAND3_X2 _42783_ (.A1(_16078_),
    .A2(_16080_),
    .A3(_15911_),
    .ZN(_16081_));
 NAND3_X2 _42784_ (.A1(_16076_),
    .A2(_16081_),
    .A3(_15645_),
    .ZN(_16082_));
 BUF_X16 _42785_ (.A(_15390_),
    .Z(_16083_));
 OR2_X2 _42786_ (.A1(_16083_),
    .A2(\icache.data_mems_6__data_mem.data_o [36]),
    .ZN(_16084_));
 INV_X8 _42787_ (.A(\icache.data_mems_7__data_mem.data_o [36]),
    .ZN(_16085_));
 NAND2_X2 _42788_ (.A1(_16085_),
    .A2(_15986_),
    .ZN(_16086_));
 NAND3_X2 _42789_ (.A1(_16084_),
    .A2(_16086_),
    .A3(_15988_),
    .ZN(_16087_));
 INV_X2 _42790_ (.A(\icache.data_mems_4__data_mem.data_o [36]),
    .ZN(_16088_));
 NAND2_X2 _42791_ (.A1(_15627_),
    .A2(_16088_),
    .ZN(_16089_));
 INV_X1 _42792_ (.A(\icache.data_mems_5__data_mem.data_o [36]),
    .ZN(_16090_));
 NAND2_X2 _42793_ (.A1(_16090_),
    .A2(_15461_),
    .ZN(_16091_));
 NAND3_X2 _42794_ (.A1(_16089_),
    .A2(_16091_),
    .A3(_15994_),
    .ZN(_16092_));
 NAND3_X2 _42795_ (.A1(_16087_),
    .A2(_16092_),
    .A3(_15656_),
    .ZN(_16093_));
 NAND2_X4 _42796_ (.A1(_16082_),
    .A2(_16093_),
    .ZN(_16094_));
 OAI21_X1 _42797_ (.A(_16072_),
    .B1(_16094_),
    .B2(_15951_),
    .ZN(_05245_));
 NAND2_X1 _42798_ (.A1(_15873_),
    .A2(\icache.lce.lce_cmd_inst.data_r [421]),
    .ZN(_16095_));
 AND2_X1 _42799_ (.A1(_15636_),
    .A2(\icache.data_mems_4__data_mem.data_o [37]),
    .ZN(_16096_));
 AND2_X1 _42800_ (.A1(_15564_),
    .A2(\icache.data_mems_5__data_mem.data_o [37]),
    .ZN(_16097_));
 OAI21_X2 _42801_ (.A(_15853_),
    .B1(_16096_),
    .B2(_16097_),
    .ZN(_16098_));
 BUF_X16 _42802_ (.A(_15812_),
    .Z(_16099_));
 INV_X8 _42803_ (.A(\icache.data_mems_6__data_mem.data_o [37]),
    .ZN(_16100_));
 NOR2_X1 _42804_ (.A1(_16100_),
    .A2(_15436_),
    .ZN(_16101_));
 AND2_X1 _42805_ (.A1(_15375_),
    .A2(\icache.data_mems_7__data_mem.data_o [37]),
    .ZN(_16102_));
 OAI21_X2 _42806_ (.A(_16099_),
    .B1(_16101_),
    .B2(_16102_),
    .ZN(_16103_));
 AOI21_X2 _42807_ (.A(_15431_),
    .B1(_16098_),
    .B2(_16103_),
    .ZN(_16104_));
 INV_X8 _42808_ (.A(\icache.data_mems_2__data_mem.data_o [37]),
    .ZN(_16105_));
 NOR2_X1 _42809_ (.A1(_16105_),
    .A2(_15452_),
    .ZN(_16106_));
 AND2_X1 _42810_ (.A1(_15454_),
    .A2(\icache.data_mems_3__data_mem.data_o [37]),
    .ZN(_16107_));
 OAI21_X2 _42811_ (.A(_15332_),
    .B1(_16106_),
    .B2(_16107_),
    .ZN(_16108_));
 INV_X2 _42812_ (.A(\icache.data_mems_0__data_mem.data_o [37]),
    .ZN(_16109_));
 NAND2_X1 _42813_ (.A1(_15627_),
    .A2(_16109_),
    .ZN(_16110_));
 INV_X1 _42814_ (.A(\icache.data_mems_1__data_mem.data_o [37]),
    .ZN(_16111_));
 BUF_X16 _42815_ (.A(_15460_),
    .Z(_16112_));
 NAND2_X1 _42816_ (.A1(_16111_),
    .A2(_16112_),
    .ZN(_16113_));
 NAND3_X2 _42817_ (.A1(_16110_),
    .A2(_16113_),
    .A3(_15576_),
    .ZN(_16114_));
 AOI21_X2 _42818_ (.A(_15449_),
    .B1(_16108_),
    .B2(_16114_),
    .ZN(_16115_));
 NOR2_X4 _42819_ (.A1(_16104_),
    .A2(_16115_),
    .ZN(_16116_));
 OAI21_X1 _42820_ (.A(_16095_),
    .B1(_16116_),
    .B2(_15951_),
    .ZN(_05246_));
 BUF_X8 _42821_ (.A(_15601_),
    .Z(_16117_));
 NAND2_X1 _42822_ (.A1(_16117_),
    .A2(\icache.lce.lce_cmd_inst.data_r [422]),
    .ZN(_16118_));
 AND2_X1 _42823_ (.A1(_15306_),
    .A2(\icache.data_mems_4__data_mem.data_o [38]),
    .ZN(_16119_));
 AND2_X1 _42824_ (.A1(_15308_),
    .A2(\icache.data_mems_5__data_mem.data_o [38]),
    .ZN(_16120_));
 OR3_X1 _42825_ (.A1(_16119_),
    .A2(_16120_),
    .A3(_15424_),
    .ZN(_16121_));
 NAND2_X1 _42826_ (.A1(_15719_),
    .A2(\icache.data_mems_6__data_mem.data_o [38]),
    .ZN(_16122_));
 INV_X8 _42827_ (.A(\icache.data_mems_7__data_mem.data_o [38]),
    .ZN(_16123_));
 OAI211_X1 _42828_ (.A(_16122_),
    .B(_15321_),
    .C1(_16035_),
    .C2(_16123_),
    .ZN(_16124_));
 AND3_X1 _42829_ (.A1(_16121_),
    .A2(_16033_),
    .A3(_16124_),
    .ZN(_16125_));
 AND2_X1 _42830_ (.A1(_15306_),
    .A2(\icache.data_mems_2__data_mem.data_o [38]),
    .ZN(_16126_));
 AND2_X1 _42831_ (.A1(_15471_),
    .A2(\icache.data_mems_3__data_mem.data_o [38]),
    .ZN(_16127_));
 OAI21_X2 _42832_ (.A(_15332_),
    .B1(_16126_),
    .B2(_16127_),
    .ZN(_16128_));
 INV_X8 _42833_ (.A(\icache.data_mems_0__data_mem.data_o [38]),
    .ZN(_16129_));
 NOR2_X2 _42834_ (.A1(_16129_),
    .A2(_15714_),
    .ZN(_16130_));
 AND2_X1 _42835_ (.A1(_15322_),
    .A2(\icache.data_mems_1__data_mem.data_o [38]),
    .ZN(_16131_));
 OAI21_X4 _42836_ (.A(_15553_),
    .B1(_16130_),
    .B2(_16131_),
    .ZN(_16132_));
 AOI21_X2 _42837_ (.A(_15449_),
    .B1(_16128_),
    .B2(_16132_),
    .ZN(_16133_));
 NOR2_X4 _42838_ (.A1(_16125_),
    .A2(_16133_),
    .ZN(_16134_));
 OAI21_X1 _42839_ (.A(_16118_),
    .B1(_16134_),
    .B2(_15951_),
    .ZN(_05247_));
 NAND2_X1 _42840_ (.A1(_16117_),
    .A2(\icache.lce.lce_cmd_inst.data_r [423]),
    .ZN(_16135_));
 AND2_X1 _42841_ (.A1(_15636_),
    .A2(\icache.data_mems_6__data_mem.data_o [39]),
    .ZN(_16136_));
 AND2_X1 _42842_ (.A1(_15564_),
    .A2(\icache.data_mems_7__data_mem.data_o [39]),
    .ZN(_16137_));
 OAI21_X1 _42843_ (.A(_15433_),
    .B1(_16136_),
    .B2(_16137_),
    .ZN(_16138_));
 INV_X1 _42844_ (.A(\icache.data_mems_4__data_mem.data_o [39]),
    .ZN(_16139_));
 NOR2_X1 _42845_ (.A1(_16139_),
    .A2(_15436_),
    .ZN(_16140_));
 AND2_X1 _42846_ (.A1(_15375_),
    .A2(\icache.data_mems_5__data_mem.data_o [39]),
    .ZN(_16141_));
 OAI21_X2 _42847_ (.A(_15370_),
    .B1(_16140_),
    .B2(_16141_),
    .ZN(_16142_));
 BUF_X16 _42848_ (.A(_16012_),
    .Z(_16143_));
 NAND3_X1 _42849_ (.A1(_16138_),
    .A2(_16142_),
    .A3(_16143_),
    .ZN(_16144_));
 AND2_X1 _42850_ (.A1(_15372_),
    .A2(\icache.data_mems_2__data_mem.data_o [39]),
    .ZN(_16145_));
 AND2_X1 _42851_ (.A1(_15454_),
    .A2(\icache.data_mems_3__data_mem.data_o [39]),
    .ZN(_16146_));
 OAI21_X2 _42852_ (.A(_15450_),
    .B1(_16145_),
    .B2(_16146_),
    .ZN(_16147_));
 OR2_X1 _42853_ (.A1(_15457_),
    .A2(\icache.data_mems_0__data_mem.data_o [39]),
    .ZN(_16148_));
 INV_X8 _42854_ (.A(\icache.data_mems_1__data_mem.data_o [39]),
    .ZN(_16149_));
 NAND2_X1 _42855_ (.A1(_16149_),
    .A2(_16112_),
    .ZN(_16150_));
 NAND3_X2 _42856_ (.A1(_16148_),
    .A2(_16150_),
    .A3(_15464_),
    .ZN(_16151_));
 NAND3_X1 _42857_ (.A1(_16147_),
    .A2(_15645_),
    .A3(_16151_),
    .ZN(_16152_));
 NAND2_X2 _42858_ (.A1(_16144_),
    .A2(_16152_),
    .ZN(_16153_));
 OAI21_X1 _42859_ (.A(_16135_),
    .B1(_16153_),
    .B2(_15951_),
    .ZN(_05248_));
 NAND2_X1 _42860_ (.A1(_16117_),
    .A2(\icache.lce.lce_cmd_inst.data_r [424]),
    .ZN(_16154_));
 BUF_X16 _42861_ (.A(_15371_),
    .Z(_16155_));
 AND2_X1 _42862_ (.A1(_16155_),
    .A2(\icache.data_mems_6__data_mem.data_o [40]),
    .ZN(_16156_));
 AND2_X1 _42863_ (.A1(_15616_),
    .A2(\icache.data_mems_7__data_mem.data_o [40]),
    .ZN(_16157_));
 OAI21_X2 _42864_ (.A(_15433_),
    .B1(_16156_),
    .B2(_16157_),
    .ZN(_16158_));
 AND2_X1 _42865_ (.A1(_15736_),
    .A2(\icache.data_mems_4__data_mem.data_o [40]),
    .ZN(_16159_));
 AND2_X1 _42866_ (.A1(_15454_),
    .A2(\icache.data_mems_5__data_mem.data_o [40]),
    .ZN(_16160_));
 OAI21_X2 _42867_ (.A(_15370_),
    .B1(_16159_),
    .B2(_16160_),
    .ZN(_16161_));
 AOI21_X2 _42868_ (.A(_15431_),
    .B1(_16158_),
    .B2(_16161_),
    .ZN(_16162_));
 AND2_X1 _42869_ (.A1(_15736_),
    .A2(\icache.data_mems_2__data_mem.data_o [40]),
    .ZN(_16163_));
 AND2_X1 _42870_ (.A1(_15438_),
    .A2(\icache.data_mems_3__data_mem.data_o [40]),
    .ZN(_16164_));
 OAI21_X2 _42871_ (.A(_15450_),
    .B1(_16163_),
    .B2(_16164_),
    .ZN(_16165_));
 INV_X1 _42872_ (.A(\icache.data_mems_0__data_mem.data_o [40]),
    .ZN(_16166_));
 NAND2_X1 _42873_ (.A1(_15756_),
    .A2(_16166_),
    .ZN(_16167_));
 INV_X8 _42874_ (.A(\icache.data_mems_1__data_mem.data_o [40]),
    .ZN(_16168_));
 BUF_X16 _42875_ (.A(_15387_),
    .Z(_16169_));
 NAND2_X1 _42876_ (.A1(_16168_),
    .A2(_16169_),
    .ZN(_16170_));
 NAND3_X2 _42877_ (.A1(_16167_),
    .A2(_16170_),
    .A3(_15464_),
    .ZN(_16171_));
 AOI21_X2 _42878_ (.A(_15449_),
    .B1(_16165_),
    .B2(_16171_),
    .ZN(_16172_));
 NOR2_X4 _42879_ (.A1(_16162_),
    .A2(_16172_),
    .ZN(_16173_));
 BUF_X8 _42880_ (.A(_15351_),
    .Z(_16174_));
 OAI21_X1 _42881_ (.A(_16154_),
    .B1(_16173_),
    .B2(_16174_),
    .ZN(_05249_));
 NAND2_X1 _42882_ (.A1(_16117_),
    .A2(\icache.lce.lce_cmd_inst.data_r [425]),
    .ZN(_16175_));
 AND2_X1 _42883_ (.A1(_15548_),
    .A2(\icache.data_mems_4__data_mem.data_o [41]),
    .ZN(_16176_));
 AND2_X1 _42884_ (.A1(_15556_),
    .A2(\icache.data_mems_5__data_mem.data_o [41]),
    .ZN(_16177_));
 OAI21_X1 _42885_ (.A(_15660_),
    .B1(_16176_),
    .B2(_16177_),
    .ZN(_16178_));
 INV_X2 _42886_ (.A(\icache.data_mems_6__data_mem.data_o [41]),
    .ZN(_16179_));
 NAND2_X2 _42887_ (.A1(_15537_),
    .A2(_16179_),
    .ZN(_16180_));
 INV_X2 _42888_ (.A(\icache.data_mems_7__data_mem.data_o [41]),
    .ZN(_16181_));
 NAND2_X2 _42889_ (.A1(_16181_),
    .A2(_15810_),
    .ZN(_16182_));
 NAND3_X2 _42890_ (.A1(_16180_),
    .A2(_16182_),
    .A3(_15812_),
    .ZN(_16183_));
 AND3_X1 _42891_ (.A1(_16178_),
    .A2(_15655_),
    .A3(_16183_),
    .ZN(_16184_));
 OR2_X1 _42892_ (.A1(_15334_),
    .A2(\icache.data_mems_2__data_mem.data_o [41]),
    .ZN(_16185_));
 INV_X8 _42893_ (.A(\icache.data_mems_3__data_mem.data_o [41]),
    .ZN(_16186_));
 NAND2_X1 _42894_ (.A1(_16186_),
    .A2(_15776_),
    .ZN(_16187_));
 NAND2_X4 _42895_ (.A1(_16185_),
    .A2(_16187_),
    .ZN(_16188_));
 NAND2_X1 _42896_ (.A1(_16188_),
    .A2(_15545_),
    .ZN(_16189_));
 INV_X8 _42897_ (.A(\icache.data_mems_0__data_mem.data_o [41]),
    .ZN(_16190_));
 NAND2_X1 _42898_ (.A1(_15537_),
    .A2(_16190_),
    .ZN(_16191_));
 INV_X1 _42899_ (.A(\icache.data_mems_1__data_mem.data_o [41]),
    .ZN(_16192_));
 NAND2_X1 _42900_ (.A1(_16192_),
    .A2(_15541_),
    .ZN(_16193_));
 NAND2_X4 _42901_ (.A1(_16191_),
    .A2(_16193_),
    .ZN(_16194_));
 BUF_X16 _42902_ (.A(_15405_),
    .Z(_16195_));
 NAND2_X1 _42903_ (.A1(_16194_),
    .A2(_16195_),
    .ZN(_16196_));
 AOI21_X1 _42904_ (.A(_15670_),
    .B1(_16189_),
    .B2(_16196_),
    .ZN(_16197_));
 OR2_X4 _42905_ (.A1(_16184_),
    .A2(_16197_),
    .ZN(_16198_));
 OAI21_X1 _42906_ (.A(_16175_),
    .B1(_16198_),
    .B2(_16174_),
    .ZN(_05250_));
 NAND2_X1 _42907_ (.A1(_16117_),
    .A2(\icache.lce.lce_cmd_inst.data_r [426]),
    .ZN(_16199_));
 BUF_X16 _42908_ (.A(_15819_),
    .Z(_16200_));
 AND2_X1 _42909_ (.A1(_15636_),
    .A2(\icache.data_mems_0__data_mem.data_o [42]),
    .ZN(_16201_));
 AND2_X1 _42910_ (.A1(_15906_),
    .A2(\icache.data_mems_1__data_mem.data_o [42]),
    .ZN(_16202_));
 OAI21_X2 _42911_ (.A(_15853_),
    .B1(_16201_),
    .B2(_16202_),
    .ZN(_16203_));
 INV_X1 _42912_ (.A(\icache.data_mems_2__data_mem.data_o [42]),
    .ZN(_16204_));
 NOR2_X1 _42913_ (.A1(_16204_),
    .A2(_15436_),
    .ZN(_16205_));
 AND2_X1 _42914_ (.A1(_15375_),
    .A2(\icache.data_mems_3__data_mem.data_o [42]),
    .ZN(_16206_));
 OAI21_X2 _42915_ (.A(_15332_),
    .B1(_16205_),
    .B2(_16206_),
    .ZN(_16207_));
 AOI21_X2 _42916_ (.A(_16200_),
    .B1(_16203_),
    .B2(_16207_),
    .ZN(_16208_));
 BUF_X32 _42917_ (.A(_15331_),
    .Z(_16209_));
 INV_X8 _42918_ (.A(\icache.data_mems_6__data_mem.data_o [42]),
    .ZN(_16210_));
 NOR2_X1 _42919_ (.A1(_16210_),
    .A2(_15452_),
    .ZN(_16211_));
 AND2_X1 _42920_ (.A1(_15454_),
    .A2(\icache.data_mems_7__data_mem.data_o [42]),
    .ZN(_16212_));
 OAI21_X2 _42921_ (.A(_16209_),
    .B1(_16211_),
    .B2(_16212_),
    .ZN(_16213_));
 OR2_X1 _42922_ (.A1(_15457_),
    .A2(\icache.data_mems_4__data_mem.data_o [42]),
    .ZN(_16214_));
 INV_X2 _42923_ (.A(\icache.data_mems_5__data_mem.data_o [42]),
    .ZN(_16215_));
 NAND2_X1 _42924_ (.A1(_16215_),
    .A2(_16112_),
    .ZN(_16216_));
 BUF_X16 _42925_ (.A(_15463_),
    .Z(_16217_));
 NAND3_X2 _42926_ (.A1(_16214_),
    .A2(_16216_),
    .A3(_16217_),
    .ZN(_16218_));
 AOI21_X2 _42927_ (.A(_15329_),
    .B1(_16213_),
    .B2(_16218_),
    .ZN(_16219_));
 NOR2_X4 _42928_ (.A1(_16208_),
    .A2(_16219_),
    .ZN(_16220_));
 OAI21_X1 _42929_ (.A(_16199_),
    .B1(_16220_),
    .B2(_16174_),
    .ZN(_05251_));
 NAND2_X1 _42930_ (.A1(_16117_),
    .A2(\icache.lce.lce_cmd_inst.data_r [427]),
    .ZN(_16221_));
 BUF_X8 _42931_ (.A(_15371_),
    .Z(_16222_));
 AND2_X2 _42932_ (.A1(_16222_),
    .A2(\icache.data_mems_6__data_mem.data_o [43]),
    .ZN(_16223_));
 BUF_X8 _42933_ (.A(_15322_),
    .Z(_16224_));
 AND2_X2 _42934_ (.A1(_16224_),
    .A2(\icache.data_mems_7__data_mem.data_o [43]),
    .ZN(_16225_));
 BUF_X16 _42935_ (.A(_15341_),
    .Z(_16226_));
 BUF_X16 _42936_ (.A(_16226_),
    .Z(_16227_));
 NOR3_X4 _42937_ (.A1(_16223_),
    .A2(_16225_),
    .A3(_16227_),
    .ZN(_16228_));
 BUF_X16 _42938_ (.A(_15330_),
    .Z(_16229_));
 BUF_X16 _42939_ (.A(_16229_),
    .Z(_16230_));
 INV_X2 _42940_ (.A(\icache.data_mems_4__data_mem.data_o [43]),
    .ZN(_16231_));
 NAND2_X1 _42941_ (.A1(_15692_),
    .A2(_16231_),
    .ZN(_16232_));
 INV_X1 _42942_ (.A(\icache.data_mems_5__data_mem.data_o [43]),
    .ZN(_16233_));
 NAND2_X1 _42943_ (.A1(_16233_),
    .A2(_16008_),
    .ZN(_16234_));
 AOI21_X2 _42944_ (.A(_16230_),
    .B1(_16232_),
    .B2(_16234_),
    .ZN(_16235_));
 OAI21_X2 _42945_ (.A(_15905_),
    .B1(_16228_),
    .B2(_16235_),
    .ZN(_16236_));
 BUF_X16 _42946_ (.A(_15644_),
    .Z(_16237_));
 INV_X8 _42947_ (.A(\icache.data_mems_0__data_mem.data_o [43]),
    .ZN(_16238_));
 NAND2_X1 _42948_ (.A1(_16035_),
    .A2(_16238_),
    .ZN(_16239_));
 INV_X1 _42949_ (.A(\icache.data_mems_1__data_mem.data_o [43]),
    .ZN(_16240_));
 NAND2_X2 _42950_ (.A1(_16240_),
    .A2(_16018_),
    .ZN(_16241_));
 AOI21_X2 _42951_ (.A(_16014_),
    .B1(_16239_),
    .B2(_16241_),
    .ZN(_16242_));
 INV_X4 _42952_ (.A(\icache.data_mems_2__data_mem.data_o [43]),
    .ZN(_16243_));
 NAND2_X1 _42953_ (.A1(_15679_),
    .A2(_16243_),
    .ZN(_16244_));
 INV_X4 _42954_ (.A(\icache.data_mems_3__data_mem.data_o [43]),
    .ZN(_16245_));
 NAND2_X1 _42955_ (.A1(_16245_),
    .A2(_15922_),
    .ZN(_16246_));
 AOI21_X2 _42956_ (.A(_16021_),
    .B1(_16244_),
    .B2(_16246_),
    .ZN(_16247_));
 OAI21_X2 _42957_ (.A(_16237_),
    .B1(_16242_),
    .B2(_16247_),
    .ZN(_16248_));
 NAND2_X4 _42958_ (.A1(_16236_),
    .A2(_16248_),
    .ZN(_16249_));
 OAI21_X1 _42959_ (.A(_16221_),
    .B1(_16249_),
    .B2(_16174_),
    .ZN(_05252_));
 NAND2_X1 _42960_ (.A1(_16117_),
    .A2(\icache.lce.lce_cmd_inst.data_r [428]),
    .ZN(_16250_));
 OR2_X1 _42961_ (.A1(_15486_),
    .A2(\icache.data_mems_4__data_mem.data_o [44]),
    .ZN(_16251_));
 INV_X1 _42962_ (.A(\icache.data_mems_5__data_mem.data_o [44]),
    .ZN(_16252_));
 BUF_X16 _42963_ (.A(_15471_),
    .Z(_16253_));
 NAND2_X1 _42964_ (.A1(_16252_),
    .A2(_16253_),
    .ZN(_16254_));
 NAND2_X1 _42965_ (.A1(_16251_),
    .A2(_16254_),
    .ZN(_16255_));
 BUF_X16 _42966_ (.A(_15369_),
    .Z(_16256_));
 NAND2_X1 _42967_ (.A1(_16255_),
    .A2(_16256_),
    .ZN(_16257_));
 OR2_X1 _42968_ (.A1(_15486_),
    .A2(\icache.data_mems_6__data_mem.data_o [44]),
    .ZN(_16258_));
 INV_X8 _42969_ (.A(\icache.data_mems_7__data_mem.data_o [44]),
    .ZN(_16259_));
 NAND2_X1 _42970_ (.A1(_16259_),
    .A2(_16253_),
    .ZN(_16260_));
 NAND2_X2 _42971_ (.A1(_16258_),
    .A2(_16260_),
    .ZN(_16261_));
 BUF_X16 _42972_ (.A(_15497_),
    .Z(_16262_));
 NAND2_X1 _42973_ (.A1(_16261_),
    .A2(_16262_),
    .ZN(_16263_));
 NAND2_X1 _42974_ (.A1(_16257_),
    .A2(_16263_),
    .ZN(_16264_));
 BUF_X16 _42975_ (.A(_15502_),
    .Z(_16265_));
 BUF_X16 _42976_ (.A(_16265_),
    .Z(_16266_));
 NAND2_X1 _42977_ (.A1(_16264_),
    .A2(_16266_),
    .ZN(_16267_));
 OR2_X2 _42978_ (.A1(_16015_),
    .A2(\icache.data_mems_0__data_mem.data_o [44]),
    .ZN(_16268_));
 INV_X8 _42979_ (.A(\icache.data_mems_1__data_mem.data_o [44]),
    .ZN(_16269_));
 NAND2_X2 _42980_ (.A1(_16269_),
    .A2(_16018_),
    .ZN(_16270_));
 AOI21_X4 _42981_ (.A(_16014_),
    .B1(_16268_),
    .B2(_16270_),
    .ZN(_16271_));
 BUF_X16 _42982_ (.A(_15322_),
    .Z(_16272_));
 OR2_X2 _42983_ (.A1(_16272_),
    .A2(\icache.data_mems_2__data_mem.data_o [44]),
    .ZN(_16273_));
 INV_X8 _42984_ (.A(\icache.data_mems_3__data_mem.data_o [44]),
    .ZN(_16274_));
 NAND2_X2 _42985_ (.A1(_16274_),
    .A2(_15922_),
    .ZN(_16275_));
 AOI21_X4 _42986_ (.A(_16021_),
    .B1(_16273_),
    .B2(_16275_),
    .ZN(_16276_));
 OAI21_X4 _42987_ (.A(_16237_),
    .B1(_16271_),
    .B2(_16276_),
    .ZN(_16277_));
 NAND2_X2 _42988_ (.A1(_16267_),
    .A2(_16277_),
    .ZN(_16278_));
 OAI21_X1 _42989_ (.A(_16250_),
    .B1(_16278_),
    .B2(_16174_),
    .ZN(_05253_));
 NAND2_X1 _42990_ (.A1(_16117_),
    .A2(\icache.lce.lce_cmd_inst.data_r [429]),
    .ZN(_16279_));
 OR2_X1 _42991_ (.A1(_15387_),
    .A2(\icache.data_mems_4__data_mem.data_o [45]),
    .ZN(_16280_));
 NAND2_X1 _42992_ (.A1(_15517_),
    .A2(_15391_),
    .ZN(_16281_));
 NAND2_X1 _42993_ (.A1(_16280_),
    .A2(_16281_),
    .ZN(_16282_));
 NAND2_X1 _42994_ (.A1(_16282_),
    .A2(_15770_),
    .ZN(_16283_));
 NAND2_X1 _42995_ (.A1(_15772_),
    .A2(_15526_),
    .ZN(_16284_));
 NAND2_X1 _42996_ (.A1(_15524_),
    .A2(_15776_),
    .ZN(_16285_));
 NAND2_X2 _42997_ (.A1(_16284_),
    .A2(_16285_),
    .ZN(_16286_));
 NAND2_X1 _42998_ (.A1(_16286_),
    .A2(_15804_),
    .ZN(_16287_));
 AOI21_X1 _42999_ (.A(_15686_),
    .B1(_16283_),
    .B2(_16287_),
    .ZN(_16288_));
 NOR2_X2 _43000_ (.A1(_15510_),
    .A2(_15518_),
    .ZN(_16289_));
 AND2_X2 _43001_ (.A1(_15488_),
    .A2(\icache.data_mems_3__data_mem.data_o [45]),
    .ZN(_16290_));
 OAI21_X2 _43002_ (.A(_15664_),
    .B1(_16289_),
    .B2(_16290_),
    .ZN(_16291_));
 OR2_X2 _43003_ (.A1(_15700_),
    .A2(\icache.data_mems_0__data_mem.data_o [45]),
    .ZN(_16292_));
 NAND2_X2 _43004_ (.A1(_15504_),
    .A2(_15495_),
    .ZN(_16293_));
 NAND3_X4 _43005_ (.A1(_16292_),
    .A2(_16293_),
    .A3(_15586_),
    .ZN(_16294_));
 AND3_X1 _43006_ (.A1(_16291_),
    .A2(_15699_),
    .A3(_16294_),
    .ZN(_16295_));
 OR2_X2 _43007_ (.A1(_16288_),
    .A2(_16295_),
    .ZN(_16296_));
 OAI21_X1 _43008_ (.A(_16279_),
    .B1(_16296_),
    .B2(_16174_),
    .ZN(_05254_));
 NAND2_X1 _43009_ (.A1(_16117_),
    .A2(\icache.lce.lce_cmd_inst.data_r [430]),
    .ZN(_16297_));
 OR2_X1 _43010_ (.A1(_15387_),
    .A2(\icache.data_mems_0__data_mem.data_o [46]),
    .ZN(_16298_));
 NAND2_X1 _43011_ (.A1(_15532_),
    .A2(_15391_),
    .ZN(_16299_));
 NAND2_X4 _43012_ (.A1(_16298_),
    .A2(_16299_),
    .ZN(_16300_));
 NAND2_X1 _43013_ (.A1(_16300_),
    .A2(_15770_),
    .ZN(_16301_));
 NAND2_X1 _43014_ (.A1(_15398_),
    .A2(_15540_),
    .ZN(_16302_));
 NAND2_X2 _43015_ (.A1(_15538_),
    .A2(_15402_),
    .ZN(_16303_));
 NAND2_X2 _43016_ (.A1(_16302_),
    .A2(_16303_),
    .ZN(_16304_));
 NAND2_X1 _43017_ (.A1(_16304_),
    .A2(_15804_),
    .ZN(_16305_));
 AOI21_X1 _43018_ (.A(_16049_),
    .B1(_16301_),
    .B2(_16305_),
    .ZN(_16306_));
 BUF_X16 _43019_ (.A(_15483_),
    .Z(_16307_));
 NAND2_X2 _43020_ (.A1(_15772_),
    .A2(\icache.data_mems_6__data_mem.data_o [46]),
    .ZN(_16308_));
 NAND2_X2 _43021_ (.A1(_15338_),
    .A2(\icache.data_mems_7__data_mem.data_o [46]),
    .ZN(_16309_));
 AOI21_X2 _43022_ (.A(_16307_),
    .B1(_16308_),
    .B2(_16309_),
    .ZN(_16310_));
 NAND2_X1 _43023_ (.A1(_15772_),
    .A2(\icache.data_mems_4__data_mem.data_o [46]),
    .ZN(_16311_));
 NAND2_X1 _43024_ (.A1(_15338_),
    .A2(\icache.data_mems_5__data_mem.data_o [46]),
    .ZN(_16312_));
 AOI21_X2 _43025_ (.A(_15664_),
    .B1(_16311_),
    .B2(_16312_),
    .ZN(_16313_));
 BUF_X16 _43026_ (.A(_15313_),
    .Z(_16314_));
 NOR3_X1 _43027_ (.A1(_16310_),
    .A2(_16313_),
    .A3(_16314_),
    .ZN(_16315_));
 OR2_X2 _43028_ (.A1(_16306_),
    .A2(_16315_),
    .ZN(_16316_));
 OAI21_X1 _43029_ (.A(_16297_),
    .B1(_16316_),
    .B2(_16174_),
    .ZN(_05256_));
 NAND2_X1 _43030_ (.A1(_16117_),
    .A2(\icache.lce.lce_cmd_inst.data_r [431]),
    .ZN(_16317_));
 NOR2_X1 _43031_ (.A1(_15583_),
    .A2(_15359_),
    .ZN(_16318_));
 BUF_X16 _43032_ (.A(net1309),
    .Z(_16319_));
 AND2_X1 _43033_ (.A1(_16319_),
    .A2(\icache.data_mems_5__data_mem.data_o [47]),
    .ZN(_16320_));
 BUF_X16 _43034_ (.A(_15310_),
    .Z(_16321_));
 OR3_X1 _43035_ (.A1(_16318_),
    .A2(_16320_),
    .A3(_16321_),
    .ZN(_16322_));
 NAND2_X1 _43036_ (.A1(_15475_),
    .A2(\icache.data_mems_7__data_mem.data_o [47]),
    .ZN(_16323_));
 BUF_X16 _43037_ (.A(_15320_),
    .Z(_16324_));
 OAI211_X2 _43038_ (.A(_16323_),
    .B(_16324_),
    .C1(_15479_),
    .C2(_15591_),
    .ZN(_16325_));
 AOI21_X1 _43039_ (.A(_15686_),
    .B1(_16322_),
    .B2(_16325_),
    .ZN(_16326_));
 BUF_X16 _43040_ (.A(_15330_),
    .Z(_16327_));
 NOR2_X2 _43041_ (.A1(_15563_),
    .A2(_15518_),
    .ZN(_16328_));
 AND2_X1 _43042_ (.A1(_15488_),
    .A2(\icache.data_mems_3__data_mem.data_o [47]),
    .ZN(_16329_));
 OAI21_X1 _43043_ (.A(_16327_),
    .B1(_16328_),
    .B2(_16329_),
    .ZN(_16330_));
 NAND2_X2 _43044_ (.A1(_15523_),
    .A2(_15572_),
    .ZN(_16331_));
 NAND2_X2 _43045_ (.A1(_15570_),
    .A2(_15495_),
    .ZN(_16332_));
 NAND3_X2 _43046_ (.A1(_16331_),
    .A2(_16332_),
    .A3(_15586_),
    .ZN(_16333_));
 AND3_X1 _43047_ (.A1(_16330_),
    .A2(_15699_),
    .A3(_16333_),
    .ZN(_16334_));
 OR2_X4 _43048_ (.A1(_16326_),
    .A2(_16334_),
    .ZN(_16335_));
 OAI21_X1 _43049_ (.A(_16317_),
    .B1(_16335_),
    .B2(_16174_),
    .ZN(_05257_));
 BUF_X8 _43050_ (.A(_15601_),
    .Z(_16336_));
 NAND2_X1 _43051_ (.A1(_16336_),
    .A2(\icache.lce.lce_cmd_inst.data_r [432]),
    .ZN(_16337_));
 OR2_X1 _43052_ (.A1(_15751_),
    .A2(\icache.data_mems_6__data_mem.data_o [48]),
    .ZN(_16338_));
 NAND2_X1 _43053_ (.A1(_15623_),
    .A2(_16015_),
    .ZN(_16339_));
 NAND2_X2 _43054_ (.A1(_16338_),
    .A2(_16339_),
    .ZN(_16340_));
 BUF_X16 _43055_ (.A(_15331_),
    .Z(_16341_));
 NAND2_X1 _43056_ (.A1(_16340_),
    .A2(_16341_),
    .ZN(_16342_));
 BUF_X8 _43057_ (.A(_15548_),
    .Z(_16343_));
 NAND2_X1 _43058_ (.A1(_16343_),
    .A2(_15630_),
    .ZN(_16344_));
 NAND2_X1 _43059_ (.A1(_15628_),
    .A2(_16253_),
    .ZN(_16345_));
 NAND2_X1 _43060_ (.A1(_16344_),
    .A2(_16345_),
    .ZN(_16346_));
 BUF_X16 _43061_ (.A(_15586_),
    .Z(_16347_));
 NAND2_X1 _43062_ (.A1(_16346_),
    .A2(_16347_),
    .ZN(_16348_));
 NAND2_X1 _43063_ (.A1(_16342_),
    .A2(_16348_),
    .ZN(_16349_));
 NAND2_X1 _43064_ (.A1(_16349_),
    .A2(_16266_),
    .ZN(_16350_));
 NOR2_X4 _43065_ (.A1(_15605_),
    .A2(_16001_),
    .ZN(_16351_));
 AND2_X1 _43066_ (.A1(_15916_),
    .A2(\icache.data_mems_1__data_mem.data_o [48]),
    .ZN(_16352_));
 NOR3_X2 _43067_ (.A1(_16351_),
    .A2(_16352_),
    .A3(_15545_),
    .ZN(_16353_));
 NAND2_X1 _43068_ (.A1(_15679_),
    .A2(_15615_),
    .ZN(_16354_));
 NAND2_X2 _43069_ (.A1(_15613_),
    .A2(_15922_),
    .ZN(_16355_));
 AOI21_X2 _43070_ (.A(_16021_),
    .B1(_16354_),
    .B2(_16355_),
    .ZN(_16356_));
 OAI21_X2 _43071_ (.A(_16237_),
    .B1(_16353_),
    .B2(_16356_),
    .ZN(_16357_));
 NAND2_X4 _43072_ (.A1(_16350_),
    .A2(_16357_),
    .ZN(_16358_));
 OAI21_X1 _43073_ (.A(_16337_),
    .B1(_16358_),
    .B2(_16174_),
    .ZN(_05258_));
 NAND2_X1 _43074_ (.A1(_16336_),
    .A2(\icache.lce.lce_cmd_inst.data_r [433]),
    .ZN(_16359_));
 BUF_X16 _43075_ (.A(_15408_),
    .Z(_16360_));
 OR2_X1 _43076_ (.A1(_15317_),
    .A2(\icache.data_mems_4__data_mem.data_o [49]),
    .ZN(_16361_));
 NAND2_X1 _43077_ (.A1(_15651_),
    .A2(_15323_),
    .ZN(_16362_));
 AND3_X1 _43078_ (.A1(_16361_),
    .A2(_16362_),
    .A3(_15369_),
    .ZN(_16363_));
 NAND2_X2 _43079_ (.A1(_15736_),
    .A2(\icache.data_mems_6__data_mem.data_o [49]),
    .ZN(_16364_));
 NAND2_X2 _43080_ (.A1(_15916_),
    .A2(\icache.data_mems_7__data_mem.data_o [49]),
    .ZN(_16365_));
 AOI21_X2 _43081_ (.A(_16307_),
    .B1(_16364_),
    .B2(_16365_),
    .ZN(_16366_));
 OAI21_X1 _43082_ (.A(_16360_),
    .B1(_16363_),
    .B2(_16366_),
    .ZN(_16367_));
 OR2_X1 _43083_ (.A1(_15411_),
    .A2(\icache.data_mems_0__data_mem.data_o [49]),
    .ZN(_16368_));
 NAND2_X1 _43084_ (.A1(_15640_),
    .A2(_15323_),
    .ZN(_16369_));
 NAND2_X2 _43085_ (.A1(_16368_),
    .A2(_16369_),
    .ZN(_16370_));
 NAND2_X1 _43086_ (.A1(_16370_),
    .A2(_15406_),
    .ZN(_16371_));
 BUF_X8 _43087_ (.A(_15833_),
    .Z(_16372_));
 NAND2_X1 _43088_ (.A1(_16343_),
    .A2(\icache.data_mems_2__data_mem.data_o [49]),
    .ZN(_16373_));
 NAND2_X1 _43089_ (.A1(_16083_),
    .A2(\icache.data_mems_3__data_mem.data_o [49]),
    .ZN(_16374_));
 NAND3_X1 _43090_ (.A1(_16373_),
    .A2(_15321_),
    .A3(_16374_),
    .ZN(_16375_));
 NAND3_X1 _43091_ (.A1(_16371_),
    .A2(_16372_),
    .A3(_16375_),
    .ZN(_16376_));
 AND2_X1 _43092_ (.A1(_16367_),
    .A2(_16376_),
    .ZN(_16377_));
 OAI21_X1 _43093_ (.A(_16359_),
    .B1(_16377_),
    .B2(_16174_),
    .ZN(_05259_));
 NAND2_X1 _43094_ (.A1(_16336_),
    .A2(\icache.lce.lce_cmd_inst.data_r [434]),
    .ZN(_16378_));
 OR2_X1 _43095_ (.A1(_15876_),
    .A2(\icache.data_mems_6__data_mem.data_o [50]),
    .ZN(_16379_));
 NAND2_X1 _43096_ (.A1(_15665_),
    .A2(_15985_),
    .ZN(_16380_));
 AND3_X1 _43097_ (.A1(_16379_),
    .A2(_16380_),
    .A3(_15378_),
    .ZN(_16381_));
 NAND2_X1 _43098_ (.A1(_15772_),
    .A2(\icache.data_mems_4__data_mem.data_o [50]),
    .ZN(_16382_));
 NAND2_X1 _43099_ (.A1(_15338_),
    .A2(\icache.data_mems_5__data_mem.data_o [50]),
    .ZN(_16383_));
 AOI21_X1 _43100_ (.A(_15331_),
    .B1(_16382_),
    .B2(_16383_),
    .ZN(_16384_));
 OR3_X1 _43101_ (.A1(_16381_),
    .A2(_15734_),
    .A3(_16384_),
    .ZN(_16385_));
 BUF_X16 _43102_ (.A(_16307_),
    .Z(_16386_));
 NOR2_X2 _43103_ (.A1(_15675_),
    .A2(_15318_),
    .ZN(_16387_));
 AND2_X1 _43104_ (.A1(_15541_),
    .A2(\icache.data_mems_1__data_mem.data_o [50]),
    .ZN(_16388_));
 OAI21_X2 _43105_ (.A(_16386_),
    .B1(_16387_),
    .B2(_16388_),
    .ZN(_16389_));
 BUF_X16 _43106_ (.A(_15644_),
    .Z(_16390_));
 BUF_X16 _43107_ (.A(_15397_),
    .Z(_16391_));
 NAND2_X1 _43108_ (.A1(_16391_),
    .A2(_15680_),
    .ZN(_16392_));
 INV_X1 _43109_ (.A(\icache.data_mems_3__data_mem.data_o [50]),
    .ZN(_16393_));
 BUF_X16 _43110_ (.A(_15308_),
    .Z(_16394_));
 NAND2_X1 _43111_ (.A1(_16393_),
    .A2(_16394_),
    .ZN(_16395_));
 BUF_X16 _43112_ (.A(_15432_),
    .Z(_16396_));
 NAND3_X2 _43113_ (.A1(_16392_),
    .A2(_16395_),
    .A3(_16396_),
    .ZN(_16397_));
 NAND3_X2 _43114_ (.A1(_16389_),
    .A2(_16390_),
    .A3(_16397_),
    .ZN(_16398_));
 NAND2_X4 _43115_ (.A1(_16385_),
    .A2(_16398_),
    .ZN(_16399_));
 BUF_X8 _43116_ (.A(_15351_),
    .Z(_16400_));
 OAI21_X1 _43117_ (.A(_16378_),
    .B1(_16399_),
    .B2(_16400_),
    .ZN(_05260_));
 NAND2_X1 _43118_ (.A1(_16336_),
    .A2(\icache.lce.lce_cmd_inst.data_r [435]),
    .ZN(_16401_));
 NOR2_X1 _43119_ (.A1(_15702_),
    .A2(_15985_),
    .ZN(_16402_));
 AND2_X1 _43120_ (.A1(_15556_),
    .A2(\icache.data_mems_1__data_mem.data_o [51]),
    .ZN(_16403_));
 NOR2_X4 _43121_ (.A1(_16402_),
    .A2(_16403_),
    .ZN(_16404_));
 NOR2_X1 _43122_ (.A1(_16404_),
    .A2(_15425_),
    .ZN(_16405_));
 BUF_X16 _43123_ (.A(_15502_),
    .Z(_16406_));
 NAND2_X2 _43124_ (.A1(_16155_),
    .A2(\icache.data_mems_2__data_mem.data_o [51]),
    .ZN(_16407_));
 BUF_X16 _43125_ (.A(_15390_),
    .Z(_16408_));
 NAND2_X2 _43126_ (.A1(_16408_),
    .A2(\icache.data_mems_3__data_mem.data_o [51]),
    .ZN(_16409_));
 AOI21_X2 _43127_ (.A(_15660_),
    .B1(_16407_),
    .B2(_16409_),
    .ZN(_16410_));
 NOR3_X1 _43128_ (.A1(_16405_),
    .A2(_16406_),
    .A3(_16410_),
    .ZN(_16411_));
 NOR2_X1 _43129_ (.A1(_15693_),
    .A2(_15359_),
    .ZN(_16412_));
 AND2_X1 _43130_ (.A1(_15362_),
    .A2(\icache.data_mems_7__data_mem.data_o [51]),
    .ZN(_16413_));
 OR3_X2 _43131_ (.A1(_16412_),
    .A2(_16413_),
    .A3(_15483_),
    .ZN(_16414_));
 OR2_X1 _43132_ (.A1(_15550_),
    .A2(\icache.data_mems_4__data_mem.data_o [51]),
    .ZN(_16415_));
 NAND2_X1 _43133_ (.A1(_15687_),
    .A2(_15421_),
    .ZN(_16416_));
 NAND2_X1 _43134_ (.A1(_16415_),
    .A2(_16416_),
    .ZN(_16417_));
 BUF_X16 _43135_ (.A(_15483_),
    .Z(_16418_));
 NAND2_X1 _43136_ (.A1(_16417_),
    .A2(_16418_),
    .ZN(_16419_));
 AOI21_X1 _43137_ (.A(_15579_),
    .B1(_16414_),
    .B2(_16419_),
    .ZN(_16420_));
 OR2_X4 _43138_ (.A1(_16411_),
    .A2(_16420_),
    .ZN(_16421_));
 OAI21_X1 _43139_ (.A(_16401_),
    .B1(_16421_),
    .B2(_16400_),
    .ZN(_05261_));
 NAND2_X1 _43140_ (.A1(_16336_),
    .A2(\icache.lce.lce_cmd_inst.data_r [436]),
    .ZN(_16422_));
 NOR2_X1 _43141_ (.A1(_15722_),
    .A2(_15359_),
    .ZN(_16423_));
 AND2_X1 _43142_ (.A1(_16319_),
    .A2(\icache.data_mems_3__data_mem.data_o [52]),
    .ZN(_16424_));
 OR3_X1 _43143_ (.A1(_16423_),
    .A2(_16424_),
    .A3(_16053_),
    .ZN(_16425_));
 NAND2_X1 _43144_ (.A1(_16394_),
    .A2(\icache.data_mems_1__data_mem.data_o [52]),
    .ZN(_16426_));
 INV_X1 _43145_ (.A(\icache.data_mems_0__data_mem.data_o [52]),
    .ZN(_16427_));
 OAI211_X2 _43146_ (.A(_16426_),
    .B(_16056_),
    .C1(_15728_),
    .C2(_16427_),
    .ZN(_16428_));
 AOI21_X1 _43147_ (.A(_16049_),
    .B1(_16425_),
    .B2(_16428_),
    .ZN(_16429_));
 NAND2_X1 _43148_ (.A1(_15736_),
    .A2(\icache.data_mems_4__data_mem.data_o [52]),
    .ZN(_16430_));
 OAI211_X2 _43149_ (.A(_16430_),
    .B(_15727_),
    .C1(_15627_),
    .C2(_15713_),
    .ZN(_16431_));
 NAND2_X1 _43150_ (.A1(_16343_),
    .A2(\icache.data_mems_6__data_mem.data_o [52]),
    .ZN(_16432_));
 NAND2_X1 _43151_ (.A1(_16083_),
    .A2(\icache.data_mems_7__data_mem.data_o [52]),
    .ZN(_16433_));
 NAND3_X1 _43152_ (.A1(_16432_),
    .A2(_15321_),
    .A3(_16433_),
    .ZN(_16434_));
 AOI21_X1 _43153_ (.A(_15579_),
    .B1(_16431_),
    .B2(_16434_),
    .ZN(_16435_));
 OR2_X4 _43154_ (.A1(_16429_),
    .A2(_16435_),
    .ZN(_16436_));
 OAI21_X1 _43155_ (.A(_16422_),
    .B1(_16436_),
    .B2(_16400_),
    .ZN(_05262_));
 NAND2_X1 _43156_ (.A1(_16336_),
    .A2(\icache.lce.lce_cmd_inst.data_r [437]),
    .ZN(_16437_));
 BUF_X8 _43157_ (.A(_15833_),
    .Z(_16438_));
 NOR2_X2 _43158_ (.A1(_15554_),
    .A2(\icache.data_mems_3__data_mem.data_o [53]),
    .ZN(_16439_));
 AOI211_X2 _43159_ (.A(_15445_),
    .B(_16439_),
    .C1(_15721_),
    .C2(_15743_),
    .ZN(_16440_));
 NAND2_X2 _43160_ (.A1(_15836_),
    .A2(\icache.data_mems_0__data_mem.data_o [53]),
    .ZN(_16441_));
 NAND2_X2 _43161_ (.A1(_15511_),
    .A2(\icache.data_mems_1__data_mem.data_o [53]),
    .ZN(_16442_));
 AOI21_X1 _43162_ (.A(_15477_),
    .B1(_16441_),
    .B2(_16442_),
    .ZN(_16443_));
 OAI21_X1 _43163_ (.A(_16438_),
    .B1(_16440_),
    .B2(_16443_),
    .ZN(_16444_));
 NAND2_X1 _43164_ (.A1(_15569_),
    .A2(_15759_),
    .ZN(_16445_));
 NAND2_X1 _43165_ (.A1(_15757_),
    .A2(_15573_),
    .ZN(_16446_));
 NAND2_X1 _43166_ (.A1(_16445_),
    .A2(_16446_),
    .ZN(_16447_));
 NAND2_X1 _43167_ (.A1(_16447_),
    .A2(_15343_),
    .ZN(_16448_));
 NAND2_X1 _43168_ (.A1(_15736_),
    .A2(_15750_),
    .ZN(_16449_));
 NAND2_X1 _43169_ (.A1(_15748_),
    .A2(_15738_),
    .ZN(_16450_));
 NAND2_X2 _43170_ (.A1(_16449_),
    .A2(_16450_),
    .ZN(_16451_));
 NAND2_X1 _43171_ (.A1(_16451_),
    .A2(_16230_),
    .ZN(_16452_));
 NAND3_X1 _43172_ (.A1(_16448_),
    .A2(_16452_),
    .A3(_15849_),
    .ZN(_16453_));
 AND2_X4 _43173_ (.A1(_16444_),
    .A2(_16453_),
    .ZN(_16454_));
 OAI21_X1 _43174_ (.A(_16437_),
    .B1(_16454_),
    .B2(_16400_),
    .ZN(_05263_));
 NAND2_X1 _43175_ (.A1(_16336_),
    .A2(\icache.lce.lce_cmd_inst.data_r [438]),
    .ZN(_16455_));
 OR2_X1 _43176_ (.A1(_15317_),
    .A2(\icache.data_mems_0__data_mem.data_o [54]),
    .ZN(_16456_));
 NAND2_X1 _43177_ (.A1(_15787_),
    .A2(_15776_),
    .ZN(_16457_));
 NAND2_X4 _43178_ (.A1(_16456_),
    .A2(_16457_),
    .ZN(_16458_));
 NAND2_X1 _43179_ (.A1(_16458_),
    .A2(_16256_),
    .ZN(_16459_));
 OR2_X1 _43180_ (.A1(_15387_),
    .A2(\icache.data_mems_2__data_mem.data_o [54]),
    .ZN(_16460_));
 NAND2_X1 _43181_ (.A1(_15782_),
    .A2(_15391_),
    .ZN(_16461_));
 NAND2_X4 _43182_ (.A1(_16460_),
    .A2(_16461_),
    .ZN(_16462_));
 NAND2_X1 _43183_ (.A1(_16462_),
    .A2(_16262_),
    .ZN(_16463_));
 NAND2_X1 _43184_ (.A1(_16459_),
    .A2(_16463_),
    .ZN(_16464_));
 NAND2_X1 _43185_ (.A1(_16464_),
    .A2(_15580_),
    .ZN(_16465_));
 NOR2_X1 _43186_ (.A1(_15767_),
    .A2(_15518_),
    .ZN(_16466_));
 AND2_X1 _43187_ (.A1(_16061_),
    .A2(\icache.data_mems_5__data_mem.data_o [54]),
    .ZN(_16467_));
 NOR3_X2 _43188_ (.A1(_16466_),
    .A2(_16467_),
    .A3(_15779_),
    .ZN(_16468_));
 NAND2_X2 _43189_ (.A1(_15491_),
    .A2(_15775_),
    .ZN(_16469_));
 NAND2_X4 _43190_ (.A1(_15773_),
    .A2(_16067_),
    .ZN(_16470_));
 AOI21_X2 _43191_ (.A(_16021_),
    .B1(_16469_),
    .B2(_16470_),
    .ZN(_16471_));
 OAI21_X2 _43192_ (.A(_16013_),
    .B1(_16468_),
    .B2(_16471_),
    .ZN(_16472_));
 NAND2_X4 _43193_ (.A1(_16465_),
    .A2(_16472_),
    .ZN(_16473_));
 OAI21_X1 _43194_ (.A(_16455_),
    .B1(_16473_),
    .B2(_16400_),
    .ZN(_05264_));
 NAND2_X1 _43195_ (.A1(_16336_),
    .A2(\icache.lce.lce_cmd_inst.data_r [439]),
    .ZN(_16474_));
 NAND2_X2 _43196_ (.A1(_15674_),
    .A2(_15816_),
    .ZN(_16475_));
 NAND2_X2 _43197_ (.A1(_15814_),
    .A2(_15986_),
    .ZN(_16476_));
 AOI21_X2 _43198_ (.A(_15567_),
    .B1(_16475_),
    .B2(_16476_),
    .ZN(_16477_));
 NAND2_X2 _43199_ (.A1(_15627_),
    .A2(_15809_),
    .ZN(_16478_));
 NAND2_X4 _43200_ (.A1(_15807_),
    .A2(_15461_),
    .ZN(_16479_));
 AOI21_X2 _43201_ (.A(_16005_),
    .B1(_16478_),
    .B2(_16479_),
    .ZN(_16480_));
 OAI21_X2 _43202_ (.A(_15905_),
    .B1(_16477_),
    .B2(_16480_),
    .ZN(_16481_));
 NOR2_X4 _43203_ (.A1(_15795_),
    .A2(_16001_),
    .ZN(_16482_));
 AND2_X1 _43204_ (.A1(_15906_),
    .A2(\icache.data_mems_1__data_mem.data_o [55]),
    .ZN(_16483_));
 OAI21_X2 _43205_ (.A(_16386_),
    .B1(_16482_),
    .B2(_16483_),
    .ZN(_16484_));
 NAND2_X2 _43206_ (.A1(_16035_),
    .A2(_15801_),
    .ZN(_16485_));
 NAND2_X2 _43207_ (.A1(_15799_),
    .A2(_15728_),
    .ZN(_16486_));
 NAND3_X2 _43208_ (.A1(_16485_),
    .A2(_16486_),
    .A3(_16396_),
    .ZN(_16487_));
 NAND3_X2 _43209_ (.A1(_16484_),
    .A2(_16390_),
    .A3(_16487_),
    .ZN(_16488_));
 NAND2_X4 _43210_ (.A1(_16481_),
    .A2(_16488_),
    .ZN(_16489_));
 OAI21_X1 _43211_ (.A(_16474_),
    .B1(_16489_),
    .B2(_16400_),
    .ZN(_05265_));
 NAND2_X1 _43212_ (.A1(_16336_),
    .A2(\icache.lce.lce_cmd_inst.data_r [440]),
    .ZN(_16490_));
 NAND2_X1 _43213_ (.A1(_15772_),
    .A2(_15839_),
    .ZN(_16491_));
 NAND2_X1 _43214_ (.A1(_15837_),
    .A2(_15955_),
    .ZN(_16492_));
 NAND2_X2 _43215_ (.A1(_16491_),
    .A2(_16492_),
    .ZN(_16493_));
 NAND2_X1 _43216_ (.A1(_16493_),
    .A2(_15610_),
    .ZN(_16494_));
 NAND2_X1 _43217_ (.A1(_15612_),
    .A2(_15845_),
    .ZN(_16495_));
 NAND2_X1 _43218_ (.A1(_15843_),
    .A2(_15616_),
    .ZN(_16496_));
 NAND2_X2 _43219_ (.A1(_16495_),
    .A2(_16496_),
    .ZN(_16497_));
 NAND2_X1 _43220_ (.A1(_16497_),
    .A2(_15619_),
    .ZN(_16498_));
 AND3_X1 _43221_ (.A1(_16494_),
    .A2(_16498_),
    .A3(_15940_),
    .ZN(_16499_));
 NOR2_X4 _43222_ (.A1(_15829_),
    .A2(_15533_),
    .ZN(_16500_));
 AND2_X2 _43223_ (.A1(_15784_),
    .A2(\icache.data_mems_3__data_mem.data_o [56]),
    .ZN(_16501_));
 OAI21_X4 _43224_ (.A(_16209_),
    .B1(_16500_),
    .B2(_16501_),
    .ZN(_16502_));
 NOR2_X4 _43225_ (.A1(_15824_),
    .A2(_15518_),
    .ZN(_16503_));
 AND2_X1 _43226_ (.A1(_15488_),
    .A2(\icache.data_mems_1__data_mem.data_o [56]),
    .ZN(_16504_));
 OAI21_X2 _43227_ (.A(_15553_),
    .B1(_16503_),
    .B2(_16504_),
    .ZN(_16505_));
 AOI21_X2 _43228_ (.A(_15449_),
    .B1(_16502_),
    .B2(_16505_),
    .ZN(_16506_));
 NOR2_X4 _43229_ (.A1(_16499_),
    .A2(_16506_),
    .ZN(_16507_));
 OAI21_X1 _43230_ (.A(_16490_),
    .B1(_16507_),
    .B2(_16400_),
    .ZN(_05267_));
 NAND2_X1 _43231_ (.A1(_16336_),
    .A2(\icache.lce.lce_cmd_inst.data_r [441]),
    .ZN(_16508_));
 NOR2_X1 _43232_ (.A1(_15858_),
    .A2(_15985_),
    .ZN(_16509_));
 AND2_X1 _43233_ (.A1(_15556_),
    .A2(\icache.data_mems_7__data_mem.data_o [57]),
    .ZN(_16510_));
 NOR2_X2 _43234_ (.A1(_16509_),
    .A2(_16510_),
    .ZN(_16511_));
 BUF_X16 _43235_ (.A(_16226_),
    .Z(_16512_));
 NOR2_X1 _43236_ (.A1(_16511_),
    .A2(_16512_),
    .ZN(_16513_));
 NAND2_X1 _43237_ (.A1(_16155_),
    .A2(\icache.data_mems_4__data_mem.data_o [57]),
    .ZN(_16514_));
 NAND2_X1 _43238_ (.A1(_16408_),
    .A2(\icache.data_mems_5__data_mem.data_o [57]),
    .ZN(_16515_));
 AOI21_X1 _43239_ (.A(_15477_),
    .B1(_16514_),
    .B2(_16515_),
    .ZN(_16516_));
 OAI21_X1 _43240_ (.A(_16360_),
    .B1(_16513_),
    .B2(_16516_),
    .ZN(_16517_));
 OR2_X1 _43241_ (.A1(_15550_),
    .A2(\icache.data_mems_0__data_mem.data_o [57]),
    .ZN(_16518_));
 NAND2_X1 _43242_ (.A1(_15867_),
    .A2(_15421_),
    .ZN(_16519_));
 NAND2_X2 _43243_ (.A1(_16518_),
    .A2(_16519_),
    .ZN(_16520_));
 NAND2_X1 _43244_ (.A1(_16520_),
    .A2(_15343_),
    .ZN(_16521_));
 OR2_X1 _43245_ (.A1(_15411_),
    .A2(\icache.data_mems_2__data_mem.data_o [57]),
    .ZN(_16522_));
 NAND2_X1 _43246_ (.A1(_15863_),
    .A2(_15323_),
    .ZN(_16523_));
 NAND2_X4 _43247_ (.A1(_16522_),
    .A2(_16523_),
    .ZN(_16524_));
 NAND2_X1 _43248_ (.A1(_16524_),
    .A2(_16230_),
    .ZN(_16525_));
 NAND3_X1 _43249_ (.A1(_16521_),
    .A2(_16525_),
    .A3(_15315_),
    .ZN(_16526_));
 AND2_X4 _43250_ (.A1(_16517_),
    .A2(_16526_),
    .ZN(_16527_));
 OAI21_X1 _43251_ (.A(_16508_),
    .B1(_16527_),
    .B2(_16400_),
    .ZN(_05268_));
 BUF_X16 _43252_ (.A(_15601_),
    .Z(_16528_));
 NAND2_X1 _43253_ (.A1(_16528_),
    .A2(\icache.lce.lce_cmd_inst.data_r [442]),
    .ZN(_16529_));
 NAND2_X1 _43254_ (.A1(_15398_),
    .A2(_15887_),
    .ZN(_16530_));
 NAND2_X1 _43255_ (.A1(_15885_),
    .A2(_15402_),
    .ZN(_16531_));
 NAND2_X2 _43256_ (.A1(_16530_),
    .A2(_16531_),
    .ZN(_16532_));
 NAND2_X1 _43257_ (.A1(_16532_),
    .A2(_16256_),
    .ZN(_16533_));
 NAND2_X1 _43258_ (.A1(_16155_),
    .A2(_15893_),
    .ZN(_16534_));
 NAND2_X1 _43259_ (.A1(_15891_),
    .A2(_15391_),
    .ZN(_16535_));
 NAND2_X2 _43260_ (.A1(_16534_),
    .A2(_16535_),
    .ZN(_16536_));
 NAND2_X1 _43261_ (.A1(_16536_),
    .A2(_16262_),
    .ZN(_16537_));
 NAND2_X1 _43262_ (.A1(_16533_),
    .A2(_16537_),
    .ZN(_16538_));
 NAND2_X1 _43263_ (.A1(_16538_),
    .A2(_16266_),
    .ZN(_16539_));
 NAND2_X1 _43264_ (.A1(_16155_),
    .A2(\icache.data_mems_2__data_mem.data_o [58]),
    .ZN(_16540_));
 BUF_X16 _43265_ (.A(_15320_),
    .Z(_16541_));
 NAND2_X1 _43266_ (.A1(_15606_),
    .A2(\icache.data_mems_3__data_mem.data_o [58]),
    .ZN(_16542_));
 AND3_X1 _43267_ (.A1(_16540_),
    .A2(_16541_),
    .A3(_16542_),
    .ZN(_16543_));
 BUF_X16 _43268_ (.A(_15394_),
    .Z(_16544_));
 OR2_X1 _43269_ (.A1(_15876_),
    .A2(\icache.data_mems_0__data_mem.data_o [58]),
    .ZN(_16545_));
 NAND2_X1 _43270_ (.A1(_15879_),
    .A2(_15985_),
    .ZN(_16546_));
 AOI21_X2 _43271_ (.A(_16544_),
    .B1(_16545_),
    .B2(_16546_),
    .ZN(_16547_));
 OAI21_X2 _43272_ (.A(_16237_),
    .B1(_16543_),
    .B2(_16547_),
    .ZN(_16548_));
 NAND2_X4 _43273_ (.A1(_16539_),
    .A2(_16548_),
    .ZN(_16549_));
 OAI21_X1 _43274_ (.A(_16529_),
    .B1(_16549_),
    .B2(_16400_),
    .ZN(_05269_));
 NAND2_X1 _43275_ (.A1(_16528_),
    .A2(\icache.lce.lce_cmd_inst.data_r [443]),
    .ZN(_16550_));
 OR2_X1 _43276_ (.A1(_15435_),
    .A2(\icache.data_mems_0__data_mem.data_o [59]),
    .ZN(_16551_));
 INV_X1 _43277_ (.A(\icache.data_mems_1__data_mem.data_o [59]),
    .ZN(_16552_));
 NAND2_X1 _43278_ (.A1(_16552_),
    .A2(_15606_),
    .ZN(_16553_));
 NAND2_X1 _43279_ (.A1(_16551_),
    .A2(_16553_),
    .ZN(_16554_));
 NAND2_X1 _43280_ (.A1(_16554_),
    .A2(_15610_),
    .ZN(_16555_));
 INV_X8 _43281_ (.A(\icache.data_mems_2__data_mem.data_o [59]),
    .ZN(_16556_));
 NAND2_X1 _43282_ (.A1(_15612_),
    .A2(_16556_),
    .ZN(_16557_));
 INV_X1 _43283_ (.A(\icache.data_mems_3__data_mem.data_o [59]),
    .ZN(_16558_));
 NAND2_X1 _43284_ (.A1(_16558_),
    .A2(_15616_),
    .ZN(_16559_));
 NAND2_X1 _43285_ (.A1(_16557_),
    .A2(_16559_),
    .ZN(_16560_));
 NAND2_X1 _43286_ (.A1(_16560_),
    .A2(_15619_),
    .ZN(_16561_));
 BUF_X16 _43287_ (.A(_15314_),
    .Z(_16562_));
 AND3_X1 _43288_ (.A1(_16555_),
    .A2(_16561_),
    .A3(_16562_),
    .ZN(_16563_));
 BUF_X16 _43289_ (.A(_15328_),
    .Z(_16564_));
 INV_X1 _43290_ (.A(\icache.data_mems_6__data_mem.data_o [59]),
    .ZN(_16565_));
 NOR2_X1 _43291_ (.A1(_16565_),
    .A2(_15478_),
    .ZN(_16566_));
 AND2_X1 _43292_ (.A1(_15876_),
    .A2(\icache.data_mems_7__data_mem.data_o [59]),
    .ZN(_16567_));
 OAI21_X2 _43293_ (.A(_16209_),
    .B1(_16566_),
    .B2(_16567_),
    .ZN(_16568_));
 INV_X1 _43294_ (.A(\icache.data_mems_4__data_mem.data_o [59]),
    .ZN(_16569_));
 NOR2_X1 _43295_ (.A1(_16569_),
    .A2(_15751_),
    .ZN(_16570_));
 AND2_X1 _43296_ (.A1(_15700_),
    .A2(\icache.data_mems_5__data_mem.data_o [59]),
    .ZN(_16571_));
 OAI21_X2 _43297_ (.A(_15553_),
    .B1(_16570_),
    .B2(_16571_),
    .ZN(_16572_));
 AOI21_X2 _43298_ (.A(_16564_),
    .B1(_16568_),
    .B2(_16572_),
    .ZN(_16573_));
 NOR2_X4 _43299_ (.A1(_16563_),
    .A2(_16573_),
    .ZN(_16574_));
 OAI21_X1 _43300_ (.A(_16550_),
    .B1(_16574_),
    .B2(_16400_),
    .ZN(_05270_));
 NAND2_X1 _43301_ (.A1(_16528_),
    .A2(\icache.lce.lce_cmd_inst.data_r [444]),
    .ZN(_16575_));
 OR2_X2 _43302_ (.A1(_16015_),
    .A2(\icache.data_mems_4__data_mem.data_o [60]),
    .ZN(_16576_));
 NAND2_X2 _43303_ (.A1(_15485_),
    .A2(_16018_),
    .ZN(_16577_));
 BUF_X16 _43304_ (.A(_15586_),
    .Z(_16578_));
 NAND3_X2 _43305_ (.A1(_16576_),
    .A2(_16577_),
    .A3(_16578_),
    .ZN(_16579_));
 BUF_X8 _43306_ (.A(_15554_),
    .Z(_16580_));
 NAND2_X2 _43307_ (.A1(_16580_),
    .A2(_15494_),
    .ZN(_16581_));
 NAND2_X2 _43308_ (.A1(_15492_),
    .A2(_15922_),
    .ZN(_16582_));
 BUF_X16 _43309_ (.A(_16229_),
    .Z(_16583_));
 NAND3_X2 _43310_ (.A1(_16581_),
    .A2(_16582_),
    .A3(_16583_),
    .ZN(_16584_));
 AOI21_X2 _43311_ (.A(_15431_),
    .B1(_16579_),
    .B2(_16584_),
    .ZN(_16585_));
 OR2_X2 _43312_ (.A1(_16015_),
    .A2(\icache.data_mems_0__data_mem.data_o [60]),
    .ZN(_16586_));
 NAND2_X2 _43313_ (.A1(_15469_),
    .A2(_16018_),
    .ZN(_16587_));
 NAND3_X2 _43314_ (.A1(_16586_),
    .A2(_16587_),
    .A3(_16578_),
    .ZN(_16588_));
 INV_X1 _43315_ (.A(\icache.data_mems_2__data_mem.data_o [60]),
    .ZN(_16589_));
 NAND2_X2 _43316_ (.A1(_16580_),
    .A2(_16589_),
    .ZN(_16590_));
 NAND2_X2 _43317_ (.A1(_15480_),
    .A2(_15922_),
    .ZN(_16591_));
 NAND3_X2 _43318_ (.A1(_16590_),
    .A2(_16591_),
    .A3(_16583_),
    .ZN(_16592_));
 AOI21_X2 _43319_ (.A(_15449_),
    .B1(_16588_),
    .B2(_16592_),
    .ZN(_16593_));
 NOR2_X4 _43320_ (.A1(_16585_),
    .A2(_16593_),
    .ZN(_16594_));
 BUF_X8 _43321_ (.A(_15351_),
    .Z(_16595_));
 OAI21_X1 _43322_ (.A(_16575_),
    .B1(_16594_),
    .B2(_16595_),
    .ZN(_05271_));
 NAND2_X1 _43323_ (.A1(_16528_),
    .A2(\icache.lce.lce_cmd_inst.data_r [445]),
    .ZN(_16596_));
 NOR2_X1 _43324_ (.A1(_15442_),
    .A2(_15505_),
    .ZN(_16597_));
 AND2_X1 _43325_ (.A1(_15390_),
    .A2(\icache.data_mems_5__data_mem.data_o [61]),
    .ZN(_16598_));
 OR3_X2 _43326_ (.A1(_16597_),
    .A2(_16598_),
    .A3(_16321_),
    .ZN(_16599_));
 OR2_X1 _43327_ (.A1(_15411_),
    .A2(\icache.data_mems_6__data_mem.data_o [61]),
    .ZN(_16600_));
 NAND2_X1 _43328_ (.A1(_15434_),
    .A2(_15511_),
    .ZN(_16601_));
 NAND2_X1 _43329_ (.A1(_16600_),
    .A2(_16601_),
    .ZN(_16602_));
 NAND2_X1 _43330_ (.A1(_16602_),
    .A2(_15514_),
    .ZN(_16603_));
 AOI21_X1 _43331_ (.A(_15686_),
    .B1(_16599_),
    .B2(_16603_),
    .ZN(_16604_));
 NOR2_X1 _43332_ (.A1(_15459_),
    .A2(_15518_),
    .ZN(_16605_));
 AND2_X1 _43333_ (.A1(_16061_),
    .A2(\icache.data_mems_1__data_mem.data_o [61]),
    .ZN(_16606_));
 OAI21_X1 _43334_ (.A(_15484_),
    .B1(_16605_),
    .B2(_16606_),
    .ZN(_16607_));
 OR2_X1 _43335_ (.A1(_15700_),
    .A2(\icache.data_mems_2__data_mem.data_o [61]),
    .ZN(_16608_));
 NAND2_X2 _43336_ (.A1(_15451_),
    .A2(_16067_),
    .ZN(_16609_));
 NAND3_X2 _43337_ (.A1(_16608_),
    .A2(_16609_),
    .A3(_15378_),
    .ZN(_16610_));
 AND3_X1 _43338_ (.A1(_16607_),
    .A2(_15430_),
    .A3(_16610_),
    .ZN(_16611_));
 OR2_X2 _43339_ (.A1(_16604_),
    .A2(_16611_),
    .ZN(_16612_));
 OAI21_X1 _43340_ (.A(_16596_),
    .B1(_16612_),
    .B2(_16595_),
    .ZN(_05272_));
 NAND2_X1 _43341_ (.A1(_16528_),
    .A2(\icache.lce.lce_cmd_inst.data_r [446]),
    .ZN(_16613_));
 NOR2_X4 _43342_ (.A1(_15413_),
    .A2(_15443_),
    .ZN(_16614_));
 AND2_X1 _43343_ (.A1(_15738_),
    .A2(\icache.data_mems_1__data_mem.data_o [62]),
    .ZN(_16615_));
 NOR3_X2 _43344_ (.A1(_16614_),
    .A2(_16615_),
    .A3(_15740_),
    .ZN(_16616_));
 NAND2_X4 _43345_ (.A1(_15747_),
    .A2(_15420_),
    .ZN(_16617_));
 NAND2_X2 _43346_ (.A1(_15418_),
    .A2(_15461_),
    .ZN(_16618_));
 AOI21_X2 _43347_ (.A(_16005_),
    .B1(_16617_),
    .B2(_16618_),
    .ZN(_16619_));
 OAI21_X2 _43348_ (.A(_15735_),
    .B1(_16616_),
    .B2(_16619_),
    .ZN(_16620_));
 BUF_X16 _43349_ (.A(_15678_),
    .Z(_16621_));
 NOR2_X2 _43350_ (.A1(_15389_),
    .A2(_15436_),
    .ZN(_16622_));
 AND2_X1 _43351_ (.A1(_15438_),
    .A2(\icache.data_mems_7__data_mem.data_o [62]),
    .ZN(_16623_));
 OAI21_X2 _43352_ (.A(_16621_),
    .B1(_16622_),
    .B2(_16623_),
    .ZN(_16624_));
 NAND2_X2 _43353_ (.A1(_15756_),
    .A2(_15401_),
    .ZN(_16625_));
 NAND2_X2 _43354_ (.A1(_15399_),
    .A2(_16169_),
    .ZN(_16626_));
 NAND3_X2 _43355_ (.A1(_16625_),
    .A2(_16626_),
    .A3(_15853_),
    .ZN(_16627_));
 NAND3_X2 _43356_ (.A1(_16624_),
    .A2(_16143_),
    .A3(_16627_),
    .ZN(_16628_));
 NAND2_X4 _43357_ (.A1(_16620_),
    .A2(_16628_),
    .ZN(_16629_));
 OAI21_X1 _43358_ (.A(_16613_),
    .B1(_16629_),
    .B2(_16595_),
    .ZN(_05273_));
 NAND2_X1 _43359_ (.A1(_16528_),
    .A2(\icache.lce.lce_cmd_inst.data_r [447]),
    .ZN(_16630_));
 BUF_X8 _43360_ (.A(_15408_),
    .Z(_16631_));
 OR2_X1 _43361_ (.A1(_15550_),
    .A2(\icache.data_mems_4__data_mem.data_o [63]),
    .ZN(_16632_));
 NAND2_X1 _43362_ (.A1(_15358_),
    .A2(_15478_),
    .ZN(_16633_));
 BUF_X16 _43363_ (.A(_15341_),
    .Z(_16634_));
 AND3_X1 _43364_ (.A1(_16632_),
    .A2(_16633_),
    .A3(_16634_),
    .ZN(_16635_));
 NAND2_X1 _43365_ (.A1(_15836_),
    .A2(\icache.data_mems_6__data_mem.data_o [63]),
    .ZN(_16636_));
 NAND2_X1 _43366_ (.A1(_15511_),
    .A2(\icache.data_mems_7__data_mem.data_o [63]),
    .ZN(_16637_));
 AOI21_X1 _43367_ (.A(_16056_),
    .B1(_16636_),
    .B2(_16637_),
    .ZN(_16638_));
 OAI21_X1 _43368_ (.A(_16631_),
    .B1(_16635_),
    .B2(_16638_),
    .ZN(_16639_));
 BUF_X16 _43369_ (.A(_15314_),
    .Z(_16640_));
 OR2_X1 _43370_ (.A1(_15334_),
    .A2(\icache.data_mems_2__data_mem.data_o [63]),
    .ZN(_16641_));
 NAND2_X1 _43371_ (.A1(_15380_),
    .A2(_15955_),
    .ZN(_16642_));
 BUF_X16 _43372_ (.A(_15330_),
    .Z(_16643_));
 AND3_X1 _43373_ (.A1(_16641_),
    .A2(_16642_),
    .A3(_16643_),
    .ZN(_16644_));
 NAND2_X1 _43374_ (.A1(_16391_),
    .A2(\icache.data_mems_0__data_mem.data_o [63]),
    .ZN(_16645_));
 NAND2_X1 _43375_ (.A1(_15475_),
    .A2(\icache.data_mems_1__data_mem.data_o [63]),
    .ZN(_16646_));
 AOI21_X1 _43376_ (.A(_16324_),
    .B1(_16645_),
    .B2(_16646_),
    .ZN(_16647_));
 OAI21_X1 _43377_ (.A(_16640_),
    .B1(_16644_),
    .B2(_16647_),
    .ZN(_16648_));
 AND2_X4 _43378_ (.A1(_16639_),
    .A2(_16648_),
    .ZN(_16649_));
 OAI21_X1 _43379_ (.A(_16630_),
    .B1(_16649_),
    .B2(_16595_),
    .ZN(_05274_));
 NAND2_X1 _43380_ (.A1(_16528_),
    .A2(\icache.lce.lce_cmd_inst.data_r [448]),
    .ZN(_16650_));
 OR2_X1 _43381_ (.A1(_15784_),
    .A2(\icache.data_mems_3__data_mem.data_o [0]),
    .ZN(_16651_));
 NAND2_X1 _43382_ (.A1(_15344_),
    .A2(_15486_),
    .ZN(_16652_));
 NAND3_X2 _43383_ (.A1(_16651_),
    .A2(_16652_),
    .A3(_15432_),
    .ZN(_16653_));
 OR2_X1 _43384_ (.A1(\icache.data_mems_1__data_mem.data_o [0]),
    .A2(_15374_),
    .ZN(_16654_));
 NAND2_X1 _43385_ (.A1(_15333_),
    .A2(_15317_),
    .ZN(_16655_));
 NAND3_X2 _43386_ (.A1(_16654_),
    .A2(_16655_),
    .A3(_15484_),
    .ZN(_16656_));
 AOI21_X2 _43387_ (.A(_16200_),
    .B1(_16653_),
    .B2(_16656_),
    .ZN(_16657_));
 NAND2_X1 _43388_ (.A1(_15398_),
    .A2(\icache.data_mems_7__data_mem.data_o [0]),
    .ZN(_16658_));
 NAND2_X1 _43389_ (.A1(_15955_),
    .A2(\icache.data_mems_6__data_mem.data_o [0]),
    .ZN(_16659_));
 NAND3_X1 _43390_ (.A1(_16658_),
    .A2(_16541_),
    .A3(_16659_),
    .ZN(_16660_));
 NAND2_X1 _43391_ (.A1(_16253_),
    .A2(\icache.data_mems_4__data_mem.data_o [0]),
    .ZN(_16661_));
 INV_X1 _43392_ (.A(\icache.data_mems_5__data_mem.data_o [0]),
    .ZN(_16662_));
 OAI211_X2 _43393_ (.A(_16661_),
    .B(_16307_),
    .C1(_15909_),
    .C2(_16662_),
    .ZN(_16663_));
 AND3_X1 _43394_ (.A1(_16660_),
    .A2(_16265_),
    .A3(_16663_),
    .ZN(_16664_));
 NOR2_X4 _43395_ (.A1(_16657_),
    .A2(_16664_),
    .ZN(_16665_));
 OAI21_X1 _43396_ (.A(_16650_),
    .B1(_16665_),
    .B2(_16595_),
    .ZN(_05275_));
 NAND2_X1 _43397_ (.A1(_16528_),
    .A2(\icache.lce.lce_cmd_inst.data_r [449]),
    .ZN(_16666_));
 INV_X2 _43398_ (.A(\icache.data_mems_5__data_mem.data_o [1]),
    .ZN(_16667_));
 NOR2_X1 _43399_ (.A1(_16667_),
    .A2(_15533_),
    .ZN(_16668_));
 AND2_X1 _43400_ (.A1(_15308_),
    .A2(\icache.data_mems_4__data_mem.data_o [1]),
    .ZN(_16669_));
 OR3_X1 _43401_ (.A1(_16668_),
    .A2(_16669_),
    .A3(_15424_),
    .ZN(_16670_));
 NAND2_X1 _43402_ (.A1(_15318_),
    .A2(\icache.data_mems_6__data_mem.data_o [1]),
    .ZN(_16671_));
 INV_X1 _43403_ (.A(\icache.data_mems_7__data_mem.data_o [1]),
    .ZN(_16672_));
 OAI211_X4 _43404_ (.A(_16671_),
    .B(_15321_),
    .C1(_15479_),
    .C2(_16672_),
    .ZN(_16673_));
 AND3_X1 _43405_ (.A1(_16670_),
    .A2(_16033_),
    .A3(_16673_),
    .ZN(_16674_));
 AND2_X1 _43406_ (.A1(_15306_),
    .A2(\icache.data_mems_3__data_mem.data_o [1]),
    .ZN(_16675_));
 AND2_X1 _43407_ (.A1(_16319_),
    .A2(\icache.data_mems_2__data_mem.data_o [1]),
    .ZN(_16676_));
 OAI21_X2 _43408_ (.A(_16209_),
    .B1(_16675_),
    .B2(_16676_),
    .ZN(_16677_));
 INV_X1 _43409_ (.A(\icache.data_mems_1__data_mem.data_o [1]),
    .ZN(_16678_));
 NOR2_X2 _43410_ (.A1(_16678_),
    .A2(_15714_),
    .ZN(_16679_));
 AND2_X1 _43411_ (.A1(_15322_),
    .A2(\icache.data_mems_0__data_mem.data_o [1]),
    .ZN(_16680_));
 OAI21_X4 _43412_ (.A(_15553_),
    .B1(_16679_),
    .B2(_16680_),
    .ZN(_16681_));
 AOI21_X2 _43413_ (.A(_15449_),
    .B1(_16677_),
    .B2(_16681_),
    .ZN(_16682_));
 NOR2_X4 _43414_ (.A1(_16674_),
    .A2(_16682_),
    .ZN(_16683_));
 OAI21_X1 _43415_ (.A(_16666_),
    .B1(_16683_),
    .B2(_16595_),
    .ZN(_05276_));
 NAND2_X1 _43416_ (.A1(_16528_),
    .A2(\icache.lce.lce_cmd_inst.data_r [450]),
    .ZN(_16684_));
 INV_X4 _43417_ (.A(\icache.data_mems_3__data_mem.data_o [2]),
    .ZN(_16685_));
 NOR2_X1 _43418_ (.A1(_16685_),
    .A2(_15359_),
    .ZN(_16686_));
 AND2_X1 _43419_ (.A1(_16319_),
    .A2(\icache.data_mems_2__data_mem.data_o [2]),
    .ZN(_16687_));
 OR3_X1 _43420_ (.A1(_16686_),
    .A2(_16687_),
    .A3(_16053_),
    .ZN(_16688_));
 NAND2_X1 _43421_ (.A1(_15636_),
    .A2(\icache.data_mems_1__data_mem.data_o [2]),
    .ZN(_16689_));
 INV_X8 _43422_ (.A(\icache.data_mems_0__data_mem.data_o [2]),
    .ZN(_16690_));
 OAI211_X2 _43423_ (.A(_16689_),
    .B(_16056_),
    .C1(_15692_),
    .C2(_16690_),
    .ZN(_16691_));
 AND3_X1 _43424_ (.A1(_16688_),
    .A2(_15474_),
    .A3(_16691_),
    .ZN(_16692_));
 INV_X4 _43425_ (.A(\icache.data_mems_7__data_mem.data_o [2]),
    .ZN(_16693_));
 NOR2_X1 _43426_ (.A1(_16693_),
    .A2(_15518_),
    .ZN(_16694_));
 AND2_X1 _43427_ (.A1(_16061_),
    .A2(\icache.data_mems_6__data_mem.data_o [2]),
    .ZN(_16695_));
 OAI21_X1 _43428_ (.A(_16327_),
    .B1(_16694_),
    .B2(_16695_),
    .ZN(_16696_));
 OR2_X1 _43429_ (.A1(_15700_),
    .A2(\icache.data_mems_5__data_mem.data_o [2]),
    .ZN(_16697_));
 INV_X1 _43430_ (.A(\icache.data_mems_4__data_mem.data_o [2]),
    .ZN(_16698_));
 NAND2_X1 _43431_ (.A1(_16698_),
    .A2(_16067_),
    .ZN(_16699_));
 NAND3_X1 _43432_ (.A1(_16697_),
    .A2(_16699_),
    .A3(_15342_),
    .ZN(_16700_));
 AOI21_X2 _43433_ (.A(_16564_),
    .B1(_16696_),
    .B2(_16700_),
    .ZN(_16701_));
 NOR2_X4 _43434_ (.A1(_16692_),
    .A2(_16701_),
    .ZN(_16702_));
 OAI21_X1 _43435_ (.A(_16684_),
    .B1(_16702_),
    .B2(_16595_),
    .ZN(_05278_));
 NAND2_X1 _43436_ (.A1(_16528_),
    .A2(\icache.lce.lce_cmd_inst.data_r [451]),
    .ZN(_16703_));
 INV_X1 _43437_ (.A(\icache.data_mems_5__data_mem.data_o [3]),
    .ZN(_16704_));
 NOR2_X4 _43438_ (.A1(_16704_),
    .A2(_15505_),
    .ZN(_16705_));
 AND2_X1 _43439_ (.A1(_15390_),
    .A2(\icache.data_mems_4__data_mem.data_o [3]),
    .ZN(_16706_));
 OR3_X1 _43440_ (.A1(_16705_),
    .A2(_16706_),
    .A3(_16321_),
    .ZN(_16707_));
 OR2_X1 _43441_ (.A1(_15411_),
    .A2(\icache.data_mems_7__data_mem.data_o [3]),
    .ZN(_16708_));
 INV_X4 _43442_ (.A(\icache.data_mems_6__data_mem.data_o [3]),
    .ZN(_16709_));
 NAND2_X1 _43443_ (.A1(_16709_),
    .A2(_15511_),
    .ZN(_16710_));
 NAND2_X2 _43444_ (.A1(_16708_),
    .A2(_16710_),
    .ZN(_16711_));
 NAND2_X1 _43445_ (.A1(_16711_),
    .A2(_15514_),
    .ZN(_16712_));
 AND3_X1 _43446_ (.A1(_16707_),
    .A2(_16033_),
    .A3(_16712_),
    .ZN(_16713_));
 BUF_X16 _43447_ (.A(_15367_),
    .Z(_16714_));
 AND2_X1 _43448_ (.A1(_15548_),
    .A2(\icache.data_mems_3__data_mem.data_o [3]),
    .ZN(_16715_));
 AND2_X2 _43449_ (.A1(_15488_),
    .A2(\icache.data_mems_2__data_mem.data_o [3]),
    .ZN(_16716_));
 OAI21_X1 _43450_ (.A(_16327_),
    .B1(_16715_),
    .B2(_16716_),
    .ZN(_16717_));
 INV_X2 _43451_ (.A(\icache.data_mems_1__data_mem.data_o [3]),
    .ZN(_16718_));
 NOR2_X2 _43452_ (.A1(_16718_),
    .A2(_15359_),
    .ZN(_16719_));
 AND2_X1 _43453_ (.A1(_15308_),
    .A2(\icache.data_mems_0__data_mem.data_o [3]),
    .ZN(_16720_));
 OAI21_X2 _43454_ (.A(_15445_),
    .B1(_16719_),
    .B2(_16720_),
    .ZN(_16721_));
 AOI21_X1 _43455_ (.A(_16714_),
    .B1(_16717_),
    .B2(_16721_),
    .ZN(_16722_));
 NOR2_X2 _43456_ (.A1(_16713_),
    .A2(_16722_),
    .ZN(_16723_));
 OAI21_X1 _43457_ (.A(_16703_),
    .B1(_16723_),
    .B2(_16595_),
    .ZN(_05279_));
 BUF_X16 _43458_ (.A(_15301_),
    .Z(_16724_));
 BUF_X8 _43459_ (.A(_16724_),
    .Z(_16725_));
 NAND2_X1 _43460_ (.A1(_16725_),
    .A2(\icache.lce.lce_cmd_inst.data_r [452]),
    .ZN(_16726_));
 INV_X4 _43461_ (.A(\icache.data_mems_7__data_mem.data_o [4]),
    .ZN(_16727_));
 NOR2_X2 _43462_ (.A1(_16727_),
    .A2(_16001_),
    .ZN(_16728_));
 AND2_X1 _43463_ (.A1(_16224_),
    .A2(\icache.data_mems_6__data_mem.data_o [4]),
    .ZN(_16729_));
 OAI21_X2 _43464_ (.A(_15433_),
    .B1(_16728_),
    .B2(_16729_),
    .ZN(_16730_));
 OR2_X1 _43465_ (.A1(_15906_),
    .A2(\icache.data_mems_5__data_mem.data_o [4]),
    .ZN(_16731_));
 INV_X1 _43466_ (.A(\icache.data_mems_4__data_mem.data_o [4]),
    .ZN(_16732_));
 NAND2_X2 _43467_ (.A1(_16732_),
    .A2(_16008_),
    .ZN(_16733_));
 NAND3_X2 _43468_ (.A1(_16731_),
    .A2(_16733_),
    .A3(_15446_),
    .ZN(_16734_));
 NAND3_X2 _43469_ (.A1(_16730_),
    .A2(_15905_),
    .A3(_16734_),
    .ZN(_16735_));
 OR2_X1 _43470_ (.A1(_16083_),
    .A2(\icache.data_mems_3__data_mem.data_o [4]),
    .ZN(_16736_));
 INV_X8 _43471_ (.A(\icache.data_mems_2__data_mem.data_o [4]),
    .ZN(_16737_));
 NAND2_X2 _43472_ (.A1(_16737_),
    .A2(_15986_),
    .ZN(_16738_));
 NAND3_X2 _43473_ (.A1(_16736_),
    .A2(_16738_),
    .A3(_15988_),
    .ZN(_16739_));
 INV_X1 _43474_ (.A(\icache.data_mems_1__data_mem.data_o [4]),
    .ZN(_16740_));
 NAND2_X1 _43475_ (.A1(_16580_),
    .A2(_16740_),
    .ZN(_16741_));
 INV_X2 _43476_ (.A(\icache.data_mems_0__data_mem.data_o [4]),
    .ZN(_16742_));
 NAND2_X1 _43477_ (.A1(_16742_),
    .A2(_15922_),
    .ZN(_16743_));
 NAND3_X2 _43478_ (.A1(_16741_),
    .A2(_16743_),
    .A3(_15994_),
    .ZN(_16744_));
 NAND3_X2 _43479_ (.A1(_16739_),
    .A2(_16744_),
    .A3(_15996_),
    .ZN(_16745_));
 NAND2_X4 _43480_ (.A1(_16735_),
    .A2(_16745_),
    .ZN(_16746_));
 OAI21_X1 _43481_ (.A(_16726_),
    .B1(_16746_),
    .B2(_16595_),
    .ZN(_05280_));
 NAND2_X1 _43482_ (.A1(_16725_),
    .A2(\icache.lce.lce_cmd_inst.data_r [453]),
    .ZN(_16747_));
 AND2_X1 _43483_ (.A1(_15306_),
    .A2(\icache.data_mems_5__data_mem.data_o [5]),
    .ZN(_16748_));
 AND2_X1 _43484_ (.A1(_15390_),
    .A2(\icache.data_mems_4__data_mem.data_o [5]),
    .ZN(_16749_));
 OR3_X2 _43485_ (.A1(_16748_),
    .A2(_16749_),
    .A3(_16321_),
    .ZN(_16750_));
 INV_X1 _43486_ (.A(\icache.data_mems_7__data_mem.data_o [5]),
    .ZN(_16751_));
 NAND2_X1 _43487_ (.A1(_15836_),
    .A2(_16751_),
    .ZN(_16752_));
 INV_X1 _43488_ (.A(\icache.data_mems_6__data_mem.data_o [5]),
    .ZN(_16753_));
 NAND2_X1 _43489_ (.A1(_16753_),
    .A2(_15511_),
    .ZN(_16754_));
 NAND2_X2 _43490_ (.A1(_16752_),
    .A2(_16754_),
    .ZN(_16755_));
 NAND2_X1 _43491_ (.A1(_16755_),
    .A2(_15514_),
    .ZN(_16756_));
 AOI21_X2 _43492_ (.A(_15686_),
    .B1(_16750_),
    .B2(_16756_),
    .ZN(_16757_));
 AND2_X1 _43493_ (.A1(_15548_),
    .A2(\icache.data_mems_3__data_mem.data_o [5]),
    .ZN(_16758_));
 AND2_X1 _43494_ (.A1(_16061_),
    .A2(\icache.data_mems_2__data_mem.data_o [5]),
    .ZN(_16759_));
 OAI21_X1 _43495_ (.A(_16327_),
    .B1(_16758_),
    .B2(_16759_),
    .ZN(_16760_));
 OR2_X1 _43496_ (.A1(_15700_),
    .A2(\icache.data_mems_1__data_mem.data_o [5]),
    .ZN(_16761_));
 INV_X8 _43497_ (.A(\icache.data_mems_0__data_mem.data_o [5]),
    .ZN(_16762_));
 NAND2_X1 _43498_ (.A1(_16762_),
    .A2(_15495_),
    .ZN(_16763_));
 NAND3_X1 _43499_ (.A1(_16761_),
    .A2(_16763_),
    .A3(_15342_),
    .ZN(_16764_));
 AND3_X1 _43500_ (.A1(_16760_),
    .A2(_15430_),
    .A3(_16764_),
    .ZN(_16765_));
 OR2_X4 _43501_ (.A1(_16757_),
    .A2(_16765_),
    .ZN(_16766_));
 OAI21_X1 _43502_ (.A(_16747_),
    .B1(_16766_),
    .B2(_16595_),
    .ZN(_05281_));
 NAND2_X1 _43503_ (.A1(_16725_),
    .A2(\icache.lce.lce_cmd_inst.data_r [454]),
    .ZN(_16767_));
 AND2_X1 _43504_ (.A1(_15554_),
    .A2(\icache.data_mems_5__data_mem.data_o [6]),
    .ZN(_16768_));
 AND2_X1 _43505_ (.A1(_15876_),
    .A2(\icache.data_mems_4__data_mem.data_o [6]),
    .ZN(_16769_));
 OR3_X1 _43506_ (.A1(_16768_),
    .A2(_16769_),
    .A3(_15394_),
    .ZN(_16770_));
 AND2_X1 _43507_ (.A1(_15548_),
    .A2(\icache.data_mems_7__data_mem.data_o [6]),
    .ZN(_16771_));
 AND2_X1 _43508_ (.A1(_15784_),
    .A2(\icache.data_mems_6__data_mem.data_o [6]),
    .ZN(_16772_));
 OR3_X1 _43509_ (.A1(_16771_),
    .A2(_16772_),
    .A3(_15405_),
    .ZN(_16773_));
 NAND2_X2 _43510_ (.A1(_16770_),
    .A2(_16773_),
    .ZN(_16774_));
 NAND2_X2 _43511_ (.A1(_16774_),
    .A2(_16266_),
    .ZN(_16775_));
 AND2_X1 _43512_ (.A1(_15372_),
    .A2(\icache.data_mems_1__data_mem.data_o [6]),
    .ZN(_16776_));
 AND2_X1 _43513_ (.A1(_15916_),
    .A2(\icache.data_mems_0__data_mem.data_o [6]),
    .ZN(_16777_));
 NOR3_X1 _43514_ (.A1(_16776_),
    .A2(_16777_),
    .A3(_15779_),
    .ZN(_16778_));
 OR2_X1 _43515_ (.A1(_16272_),
    .A2(\icache.data_mems_3__data_mem.data_o [6]),
    .ZN(_16779_));
 INV_X8 _43516_ (.A(\icache.data_mems_2__data_mem.data_o [6]),
    .ZN(_16780_));
 NAND2_X4 _43517_ (.A1(_16780_),
    .A2(_15922_),
    .ZN(_16781_));
 AOI21_X2 _43518_ (.A(_16021_),
    .B1(_16779_),
    .B2(_16781_),
    .ZN(_16782_));
 OAI21_X1 _43519_ (.A(_16237_),
    .B1(_16778_),
    .B2(_16782_),
    .ZN(_16783_));
 NAND2_X2 _43520_ (.A1(_16775_),
    .A2(_16783_),
    .ZN(_16784_));
 BUF_X16 _43521_ (.A(_15302_),
    .Z(_16785_));
 BUF_X4 _43522_ (.A(_16785_),
    .Z(_16786_));
 OAI21_X1 _43523_ (.A(_16767_),
    .B1(_16784_),
    .B2(_16786_),
    .ZN(_05282_));
 NAND2_X1 _43524_ (.A1(_16725_),
    .A2(\icache.lce.lce_cmd_inst.data_r [455]),
    .ZN(_16787_));
 INV_X1 _43525_ (.A(\icache.data_mems_5__data_mem.data_o [7]),
    .ZN(_16788_));
 NOR2_X2 _43526_ (.A1(_16788_),
    .A2(_16001_),
    .ZN(_16789_));
 AND2_X1 _43527_ (.A1(_16224_),
    .A2(\icache.data_mems_4__data_mem.data_o [7]),
    .ZN(_16790_));
 OAI21_X2 _43528_ (.A(_15853_),
    .B1(_16789_),
    .B2(_16790_),
    .ZN(_16791_));
 OR2_X1 _43529_ (.A1(_15906_),
    .A2(\icache.data_mems_7__data_mem.data_o [7]),
    .ZN(_16792_));
 INV_X4 _43530_ (.A(\icache.data_mems_6__data_mem.data_o [7]),
    .ZN(_16793_));
 NAND2_X1 _43531_ (.A1(_16793_),
    .A2(_16008_),
    .ZN(_16794_));
 NAND3_X1 _43532_ (.A1(_16792_),
    .A2(_16794_),
    .A3(_15860_),
    .ZN(_16795_));
 AOI21_X1 _43533_ (.A(_15431_),
    .B1(_16791_),
    .B2(_16795_),
    .ZN(_16796_));
 INV_X1 _43534_ (.A(\icache.data_mems_3__data_mem.data_o [7]),
    .ZN(_16797_));
 NAND2_X1 _43535_ (.A1(_16035_),
    .A2(_16797_),
    .ZN(_16798_));
 INV_X16 _43536_ (.A(\icache.data_mems_2__data_mem.data_o [7]),
    .ZN(_16799_));
 NAND2_X2 _43537_ (.A1(_16799_),
    .A2(_16018_),
    .ZN(_16800_));
 NAND3_X2 _43538_ (.A1(_16798_),
    .A2(_16800_),
    .A3(_15911_),
    .ZN(_16801_));
 INV_X1 _43539_ (.A(\icache.data_mems_1__data_mem.data_o [7]),
    .ZN(_16802_));
 NAND2_X1 _43540_ (.A1(_16580_),
    .A2(_16802_),
    .ZN(_16803_));
 INV_X4 _43541_ (.A(\icache.data_mems_0__data_mem.data_o [7]),
    .ZN(_16804_));
 BUF_X8 _43542_ (.A(_15460_),
    .Z(_16805_));
 NAND2_X1 _43543_ (.A1(_16804_),
    .A2(_16805_),
    .ZN(_16806_));
 NAND3_X2 _43544_ (.A1(_16803_),
    .A2(_16806_),
    .A3(_16217_),
    .ZN(_16807_));
 AOI21_X1 _43545_ (.A(_16714_),
    .B1(_16801_),
    .B2(_16807_),
    .ZN(_16808_));
 NOR2_X2 _43546_ (.A1(_16796_),
    .A2(_16808_),
    .ZN(_16809_));
 OAI21_X1 _43547_ (.A(_16787_),
    .B1(_16809_),
    .B2(_16786_),
    .ZN(_05283_));
 NAND2_X1 _43548_ (.A1(_16725_),
    .A2(\icache.lce.lce_cmd_inst.data_r [456]),
    .ZN(_16810_));
 AND2_X1 _43549_ (.A1(_15671_),
    .A2(\icache.data_mems_1__data_mem.data_o [8]),
    .ZN(_16811_));
 AND2_X1 _43550_ (.A1(_16224_),
    .A2(\icache.data_mems_0__data_mem.data_o [8]),
    .ZN(_16812_));
 NOR3_X2 _43551_ (.A1(_16811_),
    .A2(_16812_),
    .A3(_15740_),
    .ZN(_16813_));
 INV_X1 _43552_ (.A(\icache.data_mems_3__data_mem.data_o [8]),
    .ZN(_16814_));
 NAND2_X2 _43553_ (.A1(_15692_),
    .A2(_16814_),
    .ZN(_16815_));
 INV_X8 _43554_ (.A(\icache.data_mems_2__data_mem.data_o [8]),
    .ZN(_16816_));
 NAND2_X4 _43555_ (.A1(_16816_),
    .A2(_16008_),
    .ZN(_16817_));
 AOI21_X4 _43556_ (.A(_16005_),
    .B1(_16815_),
    .B2(_16817_),
    .ZN(_16818_));
 OAI21_X2 _43557_ (.A(_15735_),
    .B1(_16813_),
    .B2(_16818_),
    .ZN(_16819_));
 AND2_X1 _43558_ (.A1(_15671_),
    .A2(\icache.data_mems_5__data_mem.data_o [8]),
    .ZN(_16820_));
 AND2_X1 _43559_ (.A1(_16224_),
    .A2(\icache.data_mems_4__data_mem.data_o [8]),
    .ZN(_16821_));
 OAI21_X2 _43560_ (.A(_16386_),
    .B1(_16820_),
    .B2(_16821_),
    .ZN(_16822_));
 BUF_X16 _43561_ (.A(_16012_),
    .Z(_16823_));
 OR2_X1 _43562_ (.A1(_15906_),
    .A2(\icache.data_mems_7__data_mem.data_o [8]),
    .ZN(_16824_));
 INV_X4 _43563_ (.A(\icache.data_mems_6__data_mem.data_o [8]),
    .ZN(_16825_));
 NAND2_X2 _43564_ (.A1(_16825_),
    .A2(_16008_),
    .ZN(_16826_));
 NAND3_X2 _43565_ (.A1(_16824_),
    .A2(_16826_),
    .A3(_16396_),
    .ZN(_16827_));
 NAND3_X2 _43566_ (.A1(_16822_),
    .A2(_16823_),
    .A3(_16827_),
    .ZN(_16828_));
 NAND2_X4 _43567_ (.A1(_16819_),
    .A2(_16828_),
    .ZN(_16829_));
 OAI21_X1 _43568_ (.A(_16810_),
    .B1(_16829_),
    .B2(_16786_),
    .ZN(_05284_));
 NAND2_X1 _43569_ (.A1(_16725_),
    .A2(\icache.lce.lce_cmd_inst.data_r [457]),
    .ZN(_16830_));
 INV_X1 _43570_ (.A(\icache.data_mems_7__data_mem.data_o [9]),
    .ZN(_16831_));
 NOR2_X2 _43571_ (.A1(_16831_),
    .A2(_15318_),
    .ZN(_16832_));
 AND2_X1 _43572_ (.A1(_15616_),
    .A2(\icache.data_mems_6__data_mem.data_o [9]),
    .ZN(_16833_));
 OAI21_X2 _43573_ (.A(_15433_),
    .B1(_16832_),
    .B2(_16833_),
    .ZN(_16834_));
 INV_X4 _43574_ (.A(\icache.data_mems_5__data_mem.data_o [9]),
    .ZN(_16835_));
 NOR2_X2 _43575_ (.A1(_16835_),
    .A2(_15452_),
    .ZN(_16836_));
 AND2_X2 _43576_ (.A1(_15738_),
    .A2(\icache.data_mems_4__data_mem.data_o [9]),
    .ZN(_16837_));
 OAI21_X4 _43577_ (.A(_15370_),
    .B1(_16836_),
    .B2(_16837_),
    .ZN(_16838_));
 NAND3_X1 _43578_ (.A1(_16834_),
    .A2(_16838_),
    .A3(_16143_),
    .ZN(_16839_));
 INV_X1 _43579_ (.A(\icache.data_mems_3__data_mem.data_o [9]),
    .ZN(_16840_));
 NAND2_X1 _43580_ (.A1(_15747_),
    .A2(_16840_),
    .ZN(_16841_));
 INV_X16 _43581_ (.A(\icache.data_mems_2__data_mem.data_o [9]),
    .ZN(_16842_));
 NAND2_X2 _43582_ (.A1(_16842_),
    .A2(_15752_),
    .ZN(_16843_));
 NAND3_X2 _43583_ (.A1(_16841_),
    .A2(_16843_),
    .A3(_15988_),
    .ZN(_16844_));
 INV_X1 _43584_ (.A(\icache.data_mems_1__data_mem.data_o [9]),
    .ZN(_16845_));
 NAND2_X1 _43585_ (.A1(_15756_),
    .A2(_16845_),
    .ZN(_16846_));
 INV_X4 _43586_ (.A(\icache.data_mems_0__data_mem.data_o [9]),
    .ZN(_16847_));
 NAND2_X2 _43587_ (.A1(_16847_),
    .A2(_16169_),
    .ZN(_16848_));
 NAND3_X2 _43588_ (.A1(_16846_),
    .A2(_16848_),
    .A3(_15994_),
    .ZN(_16849_));
 NAND3_X1 _43589_ (.A1(_16844_),
    .A2(_16849_),
    .A3(_15996_),
    .ZN(_16850_));
 NAND2_X2 _43590_ (.A1(_16839_),
    .A2(_16850_),
    .ZN(_16851_));
 OAI21_X1 _43591_ (.A(_16830_),
    .B1(_16851_),
    .B2(_16786_),
    .ZN(_05285_));
 NAND2_X1 _43592_ (.A1(_16725_),
    .A2(\icache.lce.lce_cmd_inst.data_r [458]),
    .ZN(_16852_));
 OR2_X1 _43593_ (.A1(_15435_),
    .A2(\icache.data_mems_3__data_mem.data_o [10]),
    .ZN(_16853_));
 INV_X8 _43594_ (.A(\icache.data_mems_2__data_mem.data_o [10]),
    .ZN(_16854_));
 NAND2_X1 _43595_ (.A1(_16854_),
    .A2(_15606_),
    .ZN(_16855_));
 NAND2_X1 _43596_ (.A1(_16853_),
    .A2(_16855_),
    .ZN(_16856_));
 NAND2_X1 _43597_ (.A1(_16856_),
    .A2(_16230_),
    .ZN(_16857_));
 INV_X1 _43598_ (.A(\icache.data_mems_1__data_mem.data_o [10]),
    .ZN(_16858_));
 NAND2_X1 _43599_ (.A1(_15612_),
    .A2(_16858_),
    .ZN(_16859_));
 INV_X1 _43600_ (.A(\icache.data_mems_0__data_mem.data_o [10]),
    .ZN(_16860_));
 NAND2_X1 _43601_ (.A1(_16860_),
    .A2(_15616_),
    .ZN(_16861_));
 NAND2_X1 _43602_ (.A1(_16859_),
    .A2(_16861_),
    .ZN(_16862_));
 NAND2_X1 _43603_ (.A1(_16862_),
    .A2(_16512_),
    .ZN(_16863_));
 AND3_X1 _43604_ (.A1(_16857_),
    .A2(_16863_),
    .A3(_16562_),
    .ZN(_16864_));
 BUF_X16 _43605_ (.A(_15369_),
    .Z(_16865_));
 INV_X4 _43606_ (.A(\icache.data_mems_5__data_mem.data_o [10]),
    .ZN(_16866_));
 BUF_X16 _43607_ (.A(_15435_),
    .Z(_16867_));
 NOR2_X2 _43608_ (.A1(_16866_),
    .A2(_16867_),
    .ZN(_16868_));
 AND2_X1 _43609_ (.A1(_15916_),
    .A2(\icache.data_mems_4__data_mem.data_o [10]),
    .ZN(_16869_));
 OAI21_X2 _43610_ (.A(_16865_),
    .B1(_16868_),
    .B2(_16869_),
    .ZN(_16870_));
 OR2_X1 _43611_ (.A1(_16272_),
    .A2(\icache.data_mems_7__data_mem.data_o [10]),
    .ZN(_16871_));
 INV_X4 _43612_ (.A(\icache.data_mems_6__data_mem.data_o [10]),
    .ZN(_16872_));
 NAND2_X1 _43613_ (.A1(_16872_),
    .A2(_16805_),
    .ZN(_16873_));
 NAND3_X2 _43614_ (.A1(_16871_),
    .A2(_16873_),
    .A3(_16583_),
    .ZN(_16874_));
 AOI21_X2 _43615_ (.A(_16564_),
    .B1(_16870_),
    .B2(_16874_),
    .ZN(_16875_));
 NOR2_X4 _43616_ (.A1(_16864_),
    .A2(_16875_),
    .ZN(_16876_));
 OAI21_X1 _43617_ (.A(_16852_),
    .B1(_16876_),
    .B2(_16786_),
    .ZN(_05286_));
 NAND2_X1 _43618_ (.A1(_16725_),
    .A2(\icache.lce.lce_cmd_inst.data_r [459]),
    .ZN(_16877_));
 INV_X4 _43619_ (.A(\icache.data_mems_5__data_mem.data_o [11]),
    .ZN(_16878_));
 NOR2_X1 _43620_ (.A1(_16878_),
    .A2(_15533_),
    .ZN(_16879_));
 AND2_X1 _43621_ (.A1(_15390_),
    .A2(\icache.data_mems_4__data_mem.data_o [11]),
    .ZN(_16880_));
 OR3_X2 _43622_ (.A1(_16879_),
    .A2(_16880_),
    .A3(_15424_),
    .ZN(_16881_));
 NAND2_X1 _43623_ (.A1(_16394_),
    .A2(\icache.data_mems_6__data_mem.data_o [11]),
    .ZN(_16882_));
 INV_X1 _43624_ (.A(\icache.data_mems_7__data_mem.data_o [11]),
    .ZN(_16883_));
 OAI211_X4 _43625_ (.A(_16882_),
    .B(_15321_),
    .C1(_15479_),
    .C2(_16883_),
    .ZN(_16884_));
 AND3_X1 _43626_ (.A1(_16881_),
    .A2(_16033_),
    .A3(_16884_),
    .ZN(_16885_));
 AND2_X1 _43627_ (.A1(_15372_),
    .A2(\icache.data_mems_1__data_mem.data_o [11]),
    .ZN(_16886_));
 AND2_X1 _43628_ (.A1(_15438_),
    .A2(\icache.data_mems_0__data_mem.data_o [11]),
    .ZN(_16887_));
 OAI21_X1 _43629_ (.A(_16865_),
    .B1(_16886_),
    .B2(_16887_),
    .ZN(_16888_));
 INV_X2 _43630_ (.A(\icache.data_mems_3__data_mem.data_o [11]),
    .ZN(_16889_));
 NAND2_X1 _43631_ (.A1(_15756_),
    .A2(_16889_),
    .ZN(_16890_));
 INV_X8 _43632_ (.A(\icache.data_mems_2__data_mem.data_o [11]),
    .ZN(_16891_));
 NAND2_X4 _43633_ (.A1(_16891_),
    .A2(_16169_),
    .ZN(_16892_));
 NAND3_X2 _43634_ (.A1(_16890_),
    .A2(_16892_),
    .A3(_16583_),
    .ZN(_16893_));
 AOI21_X1 _43635_ (.A(_16714_),
    .B1(_16888_),
    .B2(_16893_),
    .ZN(_16894_));
 NOR2_X2 _43636_ (.A1(_16885_),
    .A2(_16894_),
    .ZN(_16895_));
 OAI21_X1 _43637_ (.A(_16877_),
    .B1(_16895_),
    .B2(_16786_),
    .ZN(_05287_));
 NAND2_X1 _43638_ (.A1(_16725_),
    .A2(\icache.lce.lce_cmd_inst.data_r [460]),
    .ZN(_16896_));
 AND2_X2 _43639_ (.A1(_15397_),
    .A2(\icache.data_mems_5__data_mem.data_o [12]),
    .ZN(_16897_));
 AND2_X1 _43640_ (.A1(_16319_),
    .A2(\icache.data_mems_4__data_mem.data_o [12]),
    .ZN(_16898_));
 OR3_X1 _43641_ (.A1(_16897_),
    .A2(_16898_),
    .A3(_16321_),
    .ZN(_16899_));
 NAND2_X1 _43642_ (.A1(_15636_),
    .A2(\icache.data_mems_7__data_mem.data_o [12]),
    .ZN(_16900_));
 INV_X8 _43643_ (.A(\icache.data_mems_6__data_mem.data_o [12]),
    .ZN(_16901_));
 OAI211_X4 _43644_ (.A(_16900_),
    .B(_16324_),
    .C1(_15692_),
    .C2(_16901_),
    .ZN(_16902_));
 AND3_X1 _43645_ (.A1(_16899_),
    .A2(_16033_),
    .A3(_16902_),
    .ZN(_16903_));
 AND2_X1 _43646_ (.A1(_15306_),
    .A2(\icache.data_mems_3__data_mem.data_o [12]),
    .ZN(_16904_));
 AND2_X1 _43647_ (.A1(_16061_),
    .A2(\icache.data_mems_2__data_mem.data_o [12]),
    .ZN(_16905_));
 OAI21_X1 _43648_ (.A(_16327_),
    .B1(_16904_),
    .B2(_16905_),
    .ZN(_16906_));
 INV_X1 _43649_ (.A(\icache.data_mems_1__data_mem.data_o [12]),
    .ZN(_16907_));
 NAND2_X2 _43650_ (.A1(_15491_),
    .A2(_16907_),
    .ZN(_16908_));
 INV_X8 _43651_ (.A(\icache.data_mems_0__data_mem.data_o [12]),
    .ZN(_16909_));
 NAND2_X1 _43652_ (.A1(_16909_),
    .A2(_16067_),
    .ZN(_16910_));
 NAND3_X1 _43653_ (.A1(_16908_),
    .A2(_16910_),
    .A3(_15342_),
    .ZN(_16911_));
 AOI21_X1 _43654_ (.A(_16714_),
    .B1(_16906_),
    .B2(_16911_),
    .ZN(_16912_));
 NOR2_X2 _43655_ (.A1(_16903_),
    .A2(_16912_),
    .ZN(_16913_));
 OAI21_X1 _43656_ (.A(_16896_),
    .B1(_16913_),
    .B2(_16786_),
    .ZN(_05289_));
 NAND2_X1 _43657_ (.A1(_16725_),
    .A2(\icache.lce.lce_cmd_inst.data_r [461]),
    .ZN(_16914_));
 AND2_X1 _43658_ (.A1(_16222_),
    .A2(\icache.data_mems_3__data_mem.data_o [13]),
    .ZN(_16915_));
 AND2_X2 _43659_ (.A1(_16224_),
    .A2(\icache.data_mems_2__data_mem.data_o [13]),
    .ZN(_16916_));
 OAI21_X1 _43660_ (.A(_15708_),
    .B1(_16915_),
    .B2(_16916_),
    .ZN(_16917_));
 INV_X1 _43661_ (.A(\icache.data_mems_1__data_mem.data_o [13]),
    .ZN(_16918_));
 NAND2_X1 _43662_ (.A1(_15692_),
    .A2(_16918_),
    .ZN(_16919_));
 INV_X8 _43663_ (.A(\icache.data_mems_0__data_mem.data_o [13]),
    .ZN(_16920_));
 NAND2_X2 _43664_ (.A1(_16920_),
    .A2(_16008_),
    .ZN(_16921_));
 NAND3_X2 _43665_ (.A1(_16919_),
    .A2(_16921_),
    .A3(_15446_),
    .ZN(_16922_));
 AOI21_X1 _43666_ (.A(_16200_),
    .B1(_16917_),
    .B2(_16922_),
    .ZN(_16923_));
 INV_X8 _43667_ (.A(\icache.data_mems_7__data_mem.data_o [13]),
    .ZN(_16924_));
 NOR2_X2 _43668_ (.A1(_16924_),
    .A2(_15436_),
    .ZN(_16925_));
 AND2_X1 _43669_ (.A1(_15454_),
    .A2(\icache.data_mems_6__data_mem.data_o [13]),
    .ZN(_16926_));
 OAI21_X1 _43670_ (.A(_16209_),
    .B1(_16925_),
    .B2(_16926_),
    .ZN(_16927_));
 INV_X2 _43671_ (.A(\icache.data_mems_5__data_mem.data_o [13]),
    .ZN(_16928_));
 NAND2_X1 _43672_ (.A1(_15627_),
    .A2(_16928_),
    .ZN(_16929_));
 INV_X2 _43673_ (.A(\icache.data_mems_4__data_mem.data_o [13]),
    .ZN(_16930_));
 NAND2_X1 _43674_ (.A1(_16930_),
    .A2(_15461_),
    .ZN(_16931_));
 NAND3_X1 _43675_ (.A1(_16929_),
    .A2(_16931_),
    .A3(_16217_),
    .ZN(_16932_));
 AOI21_X1 _43676_ (.A(_16564_),
    .B1(_16927_),
    .B2(_16932_),
    .ZN(_16933_));
 NOR2_X2 _43677_ (.A1(_16923_),
    .A2(_16933_),
    .ZN(_16934_));
 OAI21_X1 _43678_ (.A(_16914_),
    .B1(_16934_),
    .B2(_16786_),
    .ZN(_05290_));
 BUF_X4 _43679_ (.A(_16724_),
    .Z(_16935_));
 NAND2_X1 _43680_ (.A1(_16935_),
    .A2(\icache.lce.lce_cmd_inst.data_r [462]),
    .ZN(_16936_));
 AND2_X1 _43681_ (.A1(_15548_),
    .A2(\icache.data_mems_1__data_mem.data_o [14]),
    .ZN(_16937_));
 AND2_X1 _43682_ (.A1(_15876_),
    .A2(\icache.data_mems_0__data_mem.data_o [14]),
    .ZN(_16938_));
 OR3_X1 _43683_ (.A1(_16937_),
    .A2(_16938_),
    .A3(_15394_),
    .ZN(_16939_));
 INV_X1 _43684_ (.A(\icache.data_mems_3__data_mem.data_o [14]),
    .ZN(_16940_));
 NOR2_X4 _43685_ (.A1(_16940_),
    .A2(_15751_),
    .ZN(_16941_));
 AND2_X2 _43686_ (.A1(_15784_),
    .A2(\icache.data_mems_2__data_mem.data_o [14]),
    .ZN(_16942_));
 OR3_X1 _43687_ (.A1(_16941_),
    .A2(_16942_),
    .A3(_15405_),
    .ZN(_16943_));
 NAND2_X1 _43688_ (.A1(_16939_),
    .A2(_16943_),
    .ZN(_16944_));
 NAND2_X1 _43689_ (.A1(_16944_),
    .A2(_15580_),
    .ZN(_16945_));
 AND2_X1 _43690_ (.A1(_15372_),
    .A2(\icache.data_mems_7__data_mem.data_o [14]),
    .ZN(_16946_));
 AND2_X1 _43691_ (.A1(_15616_),
    .A2(\icache.data_mems_6__data_mem.data_o [14]),
    .ZN(_16947_));
 OAI21_X1 _43692_ (.A(_16621_),
    .B1(_16946_),
    .B2(_16947_),
    .ZN(_16948_));
 OR2_X2 _43693_ (.A1(_15776_),
    .A2(\icache.data_mems_5__data_mem.data_o [14]),
    .ZN(_16949_));
 INV_X4 _43694_ (.A(\icache.data_mems_4__data_mem.data_o [14]),
    .ZN(_16950_));
 NAND2_X2 _43695_ (.A1(_16950_),
    .A2(_16169_),
    .ZN(_16951_));
 NAND3_X4 _43696_ (.A1(_16949_),
    .A2(_16951_),
    .A3(_15901_),
    .ZN(_16952_));
 NAND3_X1 _43697_ (.A1(_16948_),
    .A2(_16823_),
    .A3(_16952_),
    .ZN(_16953_));
 NAND2_X2 _43698_ (.A1(_16945_),
    .A2(_16953_),
    .ZN(_16954_));
 OAI21_X1 _43699_ (.A(_16936_),
    .B1(_16954_),
    .B2(_16786_),
    .ZN(_05291_));
 NAND2_X1 _43700_ (.A1(_16935_),
    .A2(\icache.lce.lce_cmd_inst.data_r [463]),
    .ZN(_16955_));
 BUF_X16 _43701_ (.A(_15819_),
    .Z(_16956_));
 INV_X8 _43702_ (.A(\icache.data_mems_3__data_mem.data_o [15]),
    .ZN(_16957_));
 NOR2_X1 _43703_ (.A1(_16957_),
    .A2(_15359_),
    .ZN(_16958_));
 AND2_X1 _43704_ (.A1(_16319_),
    .A2(\icache.data_mems_2__data_mem.data_o [15]),
    .ZN(_16959_));
 OAI21_X2 _43705_ (.A(_15708_),
    .B1(_16958_),
    .B2(_16959_),
    .ZN(_16960_));
 INV_X1 _43706_ (.A(\icache.data_mems_1__data_mem.data_o [15]),
    .ZN(_16961_));
 NOR2_X2 _43707_ (.A1(_16961_),
    .A2(_15334_),
    .ZN(_16962_));
 AND2_X1 _43708_ (.A1(_15322_),
    .A2(\icache.data_mems_0__data_mem.data_o [15]),
    .ZN(_16963_));
 OAI21_X4 _43709_ (.A(_15712_),
    .B1(_16962_),
    .B2(_16963_),
    .ZN(_16964_));
 AOI21_X2 _43710_ (.A(_16956_),
    .B1(_16960_),
    .B2(_16964_),
    .ZN(_16965_));
 INV_X2 _43711_ (.A(\icache.data_mems_5__data_mem.data_o [15]),
    .ZN(_16966_));
 NOR2_X1 _43712_ (.A1(_16966_),
    .A2(_15518_),
    .ZN(_16967_));
 AND2_X1 _43713_ (.A1(_16061_),
    .A2(\icache.data_mems_4__data_mem.data_o [15]),
    .ZN(_16968_));
 OAI21_X2 _43714_ (.A(_16865_),
    .B1(_16967_),
    .B2(_16968_),
    .ZN(_16969_));
 INV_X1 _43715_ (.A(\icache.data_mems_7__data_mem.data_o [15]),
    .ZN(_16970_));
 NAND2_X1 _43716_ (.A1(_15523_),
    .A2(_16970_),
    .ZN(_16971_));
 INV_X4 _43717_ (.A(\icache.data_mems_6__data_mem.data_o [15]),
    .ZN(_16972_));
 NAND2_X1 _43718_ (.A1(_16972_),
    .A2(_15495_),
    .ZN(_16973_));
 NAND3_X2 _43719_ (.A1(_16971_),
    .A2(_16973_),
    .A3(_16583_),
    .ZN(_16974_));
 AOI21_X2 _43720_ (.A(_16564_),
    .B1(_16969_),
    .B2(_16974_),
    .ZN(_16975_));
 NOR2_X4 _43721_ (.A1(_16965_),
    .A2(_16975_),
    .ZN(_16976_));
 OAI21_X1 _43722_ (.A(_16955_),
    .B1(_16976_),
    .B2(_16786_),
    .ZN(_05292_));
 NAND2_X1 _43723_ (.A1(_16935_),
    .A2(\icache.lce.lce_cmd_inst.data_r [464]),
    .ZN(_16977_));
 AND2_X1 _43724_ (.A1(_16222_),
    .A2(\icache.data_mems_5__data_mem.data_o [16]),
    .ZN(_16978_));
 AND2_X1 _43725_ (.A1(_16224_),
    .A2(\icache.data_mems_4__data_mem.data_o [16]),
    .ZN(_16979_));
 OAI21_X1 _43726_ (.A(_15853_),
    .B1(_16978_),
    .B2(_16979_),
    .ZN(_16980_));
 INV_X1 _43727_ (.A(\icache.data_mems_7__data_mem.data_o [16]),
    .ZN(_16981_));
 NAND2_X1 _43728_ (.A1(_15692_),
    .A2(_16981_),
    .ZN(_16982_));
 INV_X8 _43729_ (.A(\icache.data_mems_6__data_mem.data_o [16]),
    .ZN(_16983_));
 NAND2_X1 _43730_ (.A1(_16983_),
    .A2(_16008_),
    .ZN(_16984_));
 NAND3_X1 _43731_ (.A1(_16982_),
    .A2(_16984_),
    .A3(_15860_),
    .ZN(_16985_));
 AOI21_X1 _43732_ (.A(_15431_),
    .B1(_16980_),
    .B2(_16985_),
    .ZN(_16986_));
 INV_X2 _43733_ (.A(\icache.data_mems_1__data_mem.data_o [16]),
    .ZN(_16987_));
 NOR2_X1 _43734_ (.A1(_16987_),
    .A2(_16867_),
    .ZN(_16988_));
 AND2_X1 _43735_ (.A1(_15916_),
    .A2(\icache.data_mems_0__data_mem.data_o [16]),
    .ZN(_16989_));
 OAI21_X1 _43736_ (.A(_16865_),
    .B1(_16988_),
    .B2(_16989_),
    .ZN(_16990_));
 OR2_X1 _43737_ (.A1(_16272_),
    .A2(\icache.data_mems_3__data_mem.data_o [16]),
    .ZN(_16991_));
 INV_X16 _43738_ (.A(\icache.data_mems_2__data_mem.data_o [16]),
    .ZN(_16992_));
 NAND2_X2 _43739_ (.A1(_16992_),
    .A2(_16805_),
    .ZN(_16993_));
 NAND3_X1 _43740_ (.A1(_16991_),
    .A2(_16993_),
    .A3(_16583_),
    .ZN(_16994_));
 AOI21_X1 _43741_ (.A(_16714_),
    .B1(_16990_),
    .B2(_16994_),
    .ZN(_16995_));
 NOR2_X2 _43742_ (.A1(_16986_),
    .A2(_16995_),
    .ZN(_16996_));
 BUF_X8 _43743_ (.A(_16785_),
    .Z(_16997_));
 OAI21_X1 _43744_ (.A(_16977_),
    .B1(_16996_),
    .B2(_16997_),
    .ZN(_05293_));
 NAND2_X1 _43745_ (.A1(_16935_),
    .A2(\icache.lce.lce_cmd_inst.data_r [465]),
    .ZN(_16998_));
 OR2_X1 _43746_ (.A1(_15387_),
    .A2(\icache.data_mems_3__data_mem.data_o [17]),
    .ZN(_16999_));
 INV_X8 _43747_ (.A(\icache.data_mems_2__data_mem.data_o [17]),
    .ZN(_17000_));
 NAND2_X1 _43748_ (.A1(_17000_),
    .A2(_15391_),
    .ZN(_17001_));
 NAND2_X4 _43749_ (.A1(_16999_),
    .A2(_17001_),
    .ZN(_17002_));
 NAND2_X1 _43750_ (.A1(_17002_),
    .A2(_16341_),
    .ZN(_17003_));
 INV_X1 _43751_ (.A(\icache.data_mems_1__data_mem.data_o [17]),
    .ZN(_17004_));
 NAND2_X1 _43752_ (.A1(_15398_),
    .A2(_17004_),
    .ZN(_17005_));
 INV_X8 _43753_ (.A(\icache.data_mems_0__data_mem.data_o [17]),
    .ZN(_17006_));
 NAND2_X1 _43754_ (.A1(_17006_),
    .A2(_15955_),
    .ZN(_17007_));
 NAND2_X1 _43755_ (.A1(_17005_),
    .A2(_17007_),
    .ZN(_17008_));
 NAND2_X1 _43756_ (.A1(_17008_),
    .A2(_16347_),
    .ZN(_17009_));
 NAND2_X4 _43757_ (.A1(_17003_),
    .A2(_17009_),
    .ZN(_17010_));
 NAND2_X1 _43758_ (.A1(_17010_),
    .A2(_15580_),
    .ZN(_17011_));
 INV_X2 _43759_ (.A(\icache.data_mems_5__data_mem.data_o [17]),
    .ZN(_17012_));
 NOR2_X2 _43760_ (.A1(_17012_),
    .A2(_15505_),
    .ZN(_17013_));
 AND2_X1 _43761_ (.A1(_16061_),
    .A2(\icache.data_mems_4__data_mem.data_o [17]),
    .ZN(_17014_));
 NOR3_X2 _43762_ (.A1(_17013_),
    .A2(_17014_),
    .A3(_15779_),
    .ZN(_17015_));
 BUF_X16 _43763_ (.A(_15609_),
    .Z(_17016_));
 OR2_X1 _43764_ (.A1(_15700_),
    .A2(\icache.data_mems_7__data_mem.data_o [17]),
    .ZN(_17017_));
 INV_X4 _43765_ (.A(\icache.data_mems_6__data_mem.data_o [17]),
    .ZN(_17018_));
 NAND2_X1 _43766_ (.A1(_17018_),
    .A2(_16067_),
    .ZN(_17019_));
 AOI21_X2 _43767_ (.A(_17016_),
    .B1(_17017_),
    .B2(_17019_),
    .ZN(_17020_));
 OAI21_X2 _43768_ (.A(_16013_),
    .B1(_17015_),
    .B2(_17020_),
    .ZN(_17021_));
 NAND2_X2 _43769_ (.A1(_17011_),
    .A2(_17021_),
    .ZN(_17022_));
 OAI21_X1 _43770_ (.A(_16998_),
    .B1(_17022_),
    .B2(_16997_),
    .ZN(_05294_));
 NAND2_X1 _43771_ (.A1(_16935_),
    .A2(\icache.lce.lce_cmd_inst.data_r [466]),
    .ZN(_17023_));
 AND2_X1 _43772_ (.A1(_16222_),
    .A2(\icache.data_mems_7__data_mem.data_o [18]),
    .ZN(_17024_));
 AND2_X1 _43773_ (.A1(_16224_),
    .A2(\icache.data_mems_6__data_mem.data_o [18]),
    .ZN(_17025_));
 OAI21_X1 _43774_ (.A(_15708_),
    .B1(_17024_),
    .B2(_17025_),
    .ZN(_17026_));
 INV_X1 _43775_ (.A(\icache.data_mems_5__data_mem.data_o [18]),
    .ZN(_17027_));
 NAND2_X2 _43776_ (.A1(_15692_),
    .A2(_17027_),
    .ZN(_17028_));
 INV_X1 _43777_ (.A(\icache.data_mems_4__data_mem.data_o [18]),
    .ZN(_17029_));
 NAND2_X4 _43778_ (.A1(_17029_),
    .A2(_16008_),
    .ZN(_17030_));
 NAND3_X4 _43779_ (.A1(_17028_),
    .A2(_17030_),
    .A3(_15446_),
    .ZN(_17031_));
 AOI21_X1 _43780_ (.A(_15431_),
    .B1(_17026_),
    .B2(_17031_),
    .ZN(_17032_));
 INV_X8 _43781_ (.A(\icache.data_mems_3__data_mem.data_o [18]),
    .ZN(_17033_));
 NOR2_X2 _43782_ (.A1(_17033_),
    .A2(_16867_),
    .ZN(_17034_));
 AND2_X1 _43783_ (.A1(_15454_),
    .A2(\icache.data_mems_2__data_mem.data_o [18]),
    .ZN(_17035_));
 OAI21_X2 _43784_ (.A(_16209_),
    .B1(_17034_),
    .B2(_17035_),
    .ZN(_17036_));
 INV_X1 _43785_ (.A(\icache.data_mems_1__data_mem.data_o [18]),
    .ZN(_17037_));
 NAND2_X1 _43786_ (.A1(_15627_),
    .A2(_17037_),
    .ZN(_17038_));
 INV_X1 _43787_ (.A(\icache.data_mems_0__data_mem.data_o [18]),
    .ZN(_17039_));
 NAND2_X1 _43788_ (.A1(_17039_),
    .A2(_15461_),
    .ZN(_17040_));
 NAND3_X1 _43789_ (.A1(_17038_),
    .A2(_17040_),
    .A3(_16217_),
    .ZN(_17041_));
 AOI21_X2 _43790_ (.A(_16714_),
    .B1(_17036_),
    .B2(_17041_),
    .ZN(_17042_));
 NOR2_X2 _43791_ (.A1(_17032_),
    .A2(_17042_),
    .ZN(_17043_));
 OAI21_X1 _43792_ (.A(_17023_),
    .B1(_17043_),
    .B2(_16997_),
    .ZN(_05295_));
 NAND2_X1 _43793_ (.A1(_16935_),
    .A2(\icache.lce.lce_cmd_inst.data_r [467]),
    .ZN(_17044_));
 AND2_X1 _43794_ (.A1(_16222_),
    .A2(\icache.data_mems_1__data_mem.data_o [19]),
    .ZN(_17045_));
 AND2_X1 _43795_ (.A1(_16224_),
    .A2(\icache.data_mems_0__data_mem.data_o [19]),
    .ZN(_17046_));
 OAI21_X2 _43796_ (.A(_15853_),
    .B1(_17045_),
    .B2(_17046_),
    .ZN(_17047_));
 OR2_X1 _43797_ (.A1(_15906_),
    .A2(\icache.data_mems_3__data_mem.data_o [19]),
    .ZN(_17048_));
 INV_X16 _43798_ (.A(\icache.data_mems_2__data_mem.data_o [19]),
    .ZN(_17049_));
 NAND2_X4 _43799_ (.A1(_17049_),
    .A2(_16008_),
    .ZN(_17050_));
 NAND3_X2 _43800_ (.A1(_17048_),
    .A2(_17050_),
    .A3(_15911_),
    .ZN(_17051_));
 AOI21_X2 _43801_ (.A(_16956_),
    .B1(_17047_),
    .B2(_17051_),
    .ZN(_17052_));
 INV_X1 _43802_ (.A(\icache.data_mems_7__data_mem.data_o [19]),
    .ZN(_17053_));
 NAND2_X1 _43803_ (.A1(_15674_),
    .A2(_17053_),
    .ZN(_17054_));
 INV_X4 _43804_ (.A(\icache.data_mems_6__data_mem.data_o [19]),
    .ZN(_17055_));
 NAND2_X1 _43805_ (.A1(_17055_),
    .A2(_16018_),
    .ZN(_17056_));
 NAND3_X1 _43806_ (.A1(_17054_),
    .A2(_17056_),
    .A3(_15911_),
    .ZN(_17057_));
 INV_X1 _43807_ (.A(\icache.data_mems_5__data_mem.data_o [19]),
    .ZN(_17058_));
 NAND2_X1 _43808_ (.A1(_16580_),
    .A2(_17058_),
    .ZN(_17059_));
 INV_X1 _43809_ (.A(\icache.data_mems_4__data_mem.data_o [19]),
    .ZN(_17060_));
 NAND2_X1 _43810_ (.A1(_17060_),
    .A2(_16805_),
    .ZN(_17061_));
 NAND3_X1 _43811_ (.A1(_17059_),
    .A2(_17061_),
    .A3(_16217_),
    .ZN(_17062_));
 AOI21_X1 _43812_ (.A(_16564_),
    .B1(_17057_),
    .B2(_17062_),
    .ZN(_17063_));
 NOR2_X2 _43813_ (.A1(_17052_),
    .A2(_17063_),
    .ZN(_17064_));
 OAI21_X1 _43814_ (.A(_17044_),
    .B1(_17064_),
    .B2(_16997_),
    .ZN(_05296_));
 NAND2_X1 _43815_ (.A1(_16935_),
    .A2(\icache.lce.lce_cmd_inst.data_r [468]),
    .ZN(_17065_));
 AND2_X1 _43816_ (.A1(_15397_),
    .A2(\icache.data_mems_3__data_mem.data_o [20]),
    .ZN(_17066_));
 AND2_X1 _43817_ (.A1(_16319_),
    .A2(\icache.data_mems_2__data_mem.data_o [20]),
    .ZN(_17067_));
 BUF_X16 _43818_ (.A(net1304),
    .Z(_17068_));
 OR3_X1 _43819_ (.A1(_17066_),
    .A2(_17067_),
    .A3(_17068_),
    .ZN(_17069_));
 NAND2_X1 _43820_ (.A1(_16222_),
    .A2(\icache.data_mems_1__data_mem.data_o [20]),
    .ZN(_17070_));
 INV_X1 _43821_ (.A(\icache.data_mems_0__data_mem.data_o [20]),
    .ZN(_17071_));
 OAI211_X2 _43822_ (.A(_17070_),
    .B(_16056_),
    .C1(_15747_),
    .C2(_17071_),
    .ZN(_17072_));
 AOI21_X1 _43823_ (.A(_16049_),
    .B1(_17069_),
    .B2(_17072_),
    .ZN(_17073_));
 OR2_X1 _43824_ (.A1(_15411_),
    .A2(\icache.data_mems_5__data_mem.data_o [20]),
    .ZN(_17074_));
 INV_X1 _43825_ (.A(\icache.data_mems_4__data_mem.data_o [20]),
    .ZN(_17075_));
 NAND2_X1 _43826_ (.A1(_17075_),
    .A2(_15323_),
    .ZN(_17076_));
 NAND2_X2 _43827_ (.A1(_17074_),
    .A2(_17076_),
    .ZN(_17077_));
 NAND2_X1 _43828_ (.A1(_17077_),
    .A2(_16195_),
    .ZN(_17078_));
 INV_X1 _43829_ (.A(\icache.data_mems_7__data_mem.data_o [20]),
    .ZN(_17079_));
 NAND2_X1 _43830_ (.A1(_15417_),
    .A2(_17079_),
    .ZN(_17080_));
 INV_X1 _43831_ (.A(\icache.data_mems_6__data_mem.data_o [20]),
    .ZN(_17081_));
 NAND2_X1 _43832_ (.A1(_17081_),
    .A2(_15421_),
    .ZN(_17082_));
 NAND2_X1 _43833_ (.A1(_17080_),
    .A2(_17082_),
    .ZN(_17083_));
 NAND2_X1 _43834_ (.A1(_17083_),
    .A2(_16541_),
    .ZN(_17084_));
 AOI21_X1 _43835_ (.A(_15579_),
    .B1(_17078_),
    .B2(_17084_),
    .ZN(_17085_));
 OR2_X4 _43836_ (.A1(_17073_),
    .A2(_17085_),
    .ZN(_17086_));
 OAI21_X1 _43837_ (.A(_17065_),
    .B1(_17086_),
    .B2(_16997_),
    .ZN(_05297_));
 NAND2_X1 _43838_ (.A1(_16935_),
    .A2(\icache.lce.lce_cmd_inst.data_r [469]),
    .ZN(_17087_));
 INV_X2 _43839_ (.A(\icache.data_mems_5__data_mem.data_o [21]),
    .ZN(_17088_));
 NOR2_X1 _43840_ (.A1(_17088_),
    .A2(_15810_),
    .ZN(_17089_));
 AND2_X1 _43841_ (.A1(_15550_),
    .A2(\icache.data_mems_4__data_mem.data_o [21]),
    .ZN(_17090_));
 OR3_X2 _43842_ (.A1(_17089_),
    .A2(_17090_),
    .A3(_15394_),
    .ZN(_17091_));
 OR2_X1 _43843_ (.A1(_15486_),
    .A2(\icache.data_mems_7__data_mem.data_o [21]),
    .ZN(_17092_));
 INV_X4 _43844_ (.A(\icache.data_mems_6__data_mem.data_o [21]),
    .ZN(_17093_));
 NAND2_X1 _43845_ (.A1(_17093_),
    .A2(_16253_),
    .ZN(_17094_));
 NAND2_X2 _43846_ (.A1(_17092_),
    .A2(_17094_),
    .ZN(_17095_));
 NAND2_X1 _43847_ (.A1(_17095_),
    .A2(_16262_),
    .ZN(_17096_));
 NAND2_X4 _43848_ (.A1(_17091_),
    .A2(_17096_),
    .ZN(_17097_));
 NAND2_X1 _43849_ (.A1(_17097_),
    .A2(_16266_),
    .ZN(_17098_));
 AND2_X2 _43850_ (.A1(_16391_),
    .A2(\icache.data_mems_3__data_mem.data_o [21]),
    .ZN(_17099_));
 AND2_X2 _43851_ (.A1(_16394_),
    .A2(\icache.data_mems_2__data_mem.data_o [21]),
    .ZN(_17100_));
 OAI21_X1 _43852_ (.A(_16621_),
    .B1(_17099_),
    .B2(_17100_),
    .ZN(_17101_));
 OR2_X1 _43853_ (.A1(_15318_),
    .A2(\icache.data_mems_1__data_mem.data_o [21]),
    .ZN(_17102_));
 INV_X8 _43854_ (.A(\icache.data_mems_0__data_mem.data_o [21]),
    .ZN(_17103_));
 NAND2_X2 _43855_ (.A1(_17103_),
    .A2(_15324_),
    .ZN(_17104_));
 NAND3_X1 _43856_ (.A1(_17102_),
    .A2(_17104_),
    .A3(_15901_),
    .ZN(_17105_));
 NAND3_X1 _43857_ (.A1(_17101_),
    .A2(_16390_),
    .A3(_17105_),
    .ZN(_17106_));
 NAND2_X2 _43858_ (.A1(_17098_),
    .A2(_17106_),
    .ZN(_17107_));
 OAI21_X1 _43859_ (.A(_17087_),
    .B1(_17107_),
    .B2(_16997_),
    .ZN(_05298_));
 NAND2_X1 _43860_ (.A1(_16935_),
    .A2(\icache.lce.lce_cmd_inst.data_r [470]),
    .ZN(_17108_));
 AND2_X1 _43861_ (.A1(_15569_),
    .A2(\icache.data_mems_3__data_mem.data_o [22]),
    .ZN(_17109_));
 AND2_X2 _43862_ (.A1(_15375_),
    .A2(\icache.data_mems_2__data_mem.data_o [22]),
    .ZN(_17110_));
 OAI21_X2 _43863_ (.A(_15708_),
    .B1(_17109_),
    .B2(_17110_),
    .ZN(_17111_));
 AND2_X1 _43864_ (.A1(_15569_),
    .A2(\icache.data_mems_1__data_mem.data_o [22]),
    .ZN(_17112_));
 AND2_X1 _43865_ (.A1(_16272_),
    .A2(\icache.data_mems_0__data_mem.data_o [22]),
    .ZN(_17113_));
 OAI21_X2 _43866_ (.A(_15712_),
    .B1(_17112_),
    .B2(_17113_),
    .ZN(_17114_));
 AOI21_X2 _43867_ (.A(_16956_),
    .B1(_17111_),
    .B2(_17114_),
    .ZN(_17115_));
 INV_X8 _43868_ (.A(\icache.data_mems_7__data_mem.data_o [22]),
    .ZN(_17116_));
 NOR2_X2 _43869_ (.A1(_17116_),
    .A2(_15318_),
    .ZN(_17117_));
 AND2_X2 _43870_ (.A1(_15616_),
    .A2(\icache.data_mems_6__data_mem.data_o [22]),
    .ZN(_17118_));
 OAI21_X1 _43871_ (.A(_16209_),
    .B1(_17117_),
    .B2(_17118_),
    .ZN(_17119_));
 INV_X1 _43872_ (.A(\icache.data_mems_5__data_mem.data_o [22]),
    .ZN(_17120_));
 NOR2_X2 _43873_ (.A1(_17120_),
    .A2(_15335_),
    .ZN(_17121_));
 AND2_X2 _43874_ (.A1(_15346_),
    .A2(\icache.data_mems_4__data_mem.data_o [22]),
    .ZN(_17122_));
 OAI21_X2 _43875_ (.A(_15553_),
    .B1(_17121_),
    .B2(_17122_),
    .ZN(_17123_));
 AOI21_X1 _43876_ (.A(_16564_),
    .B1(_17119_),
    .B2(_17123_),
    .ZN(_17124_));
 NOR2_X2 _43877_ (.A1(_17115_),
    .A2(_17124_),
    .ZN(_17125_));
 OAI21_X1 _43878_ (.A(_17108_),
    .B1(_17125_),
    .B2(_16997_),
    .ZN(_05300_));
 NAND2_X1 _43879_ (.A1(_16935_),
    .A2(\icache.lce.lce_cmd_inst.data_r [471]),
    .ZN(_17126_));
 AND2_X1 _43880_ (.A1(_15554_),
    .A2(\icache.data_mems_7__data_mem.data_o [23]),
    .ZN(_17127_));
 AND2_X1 _43881_ (.A1(_15550_),
    .A2(\icache.data_mems_6__data_mem.data_o [23]),
    .ZN(_17128_));
 OR3_X4 _43882_ (.A1(_17127_),
    .A2(_17128_),
    .A3(_15609_),
    .ZN(_17129_));
 INV_X1 _43883_ (.A(\icache.data_mems_5__data_mem.data_o [23]),
    .ZN(_17130_));
 NAND2_X1 _43884_ (.A1(_16343_),
    .A2(_17130_),
    .ZN(_17131_));
 INV_X1 _43885_ (.A(\icache.data_mems_4__data_mem.data_o [23]),
    .ZN(_17132_));
 NAND2_X1 _43886_ (.A1(_17132_),
    .A2(_15564_),
    .ZN(_17133_));
 NAND2_X1 _43887_ (.A1(_17131_),
    .A2(_17133_),
    .ZN(_17134_));
 NAND2_X1 _43888_ (.A1(_17134_),
    .A2(_16347_),
    .ZN(_17135_));
 NAND2_X4 _43889_ (.A1(_17129_),
    .A2(_17135_),
    .ZN(_17136_));
 NAND2_X1 _43890_ (.A1(_17136_),
    .A2(_16266_),
    .ZN(_17137_));
 OR2_X1 _43891_ (.A1(_16015_),
    .A2(\icache.data_mems_1__data_mem.data_o [23]),
    .ZN(_17138_));
 INV_X8 _43892_ (.A(\icache.data_mems_0__data_mem.data_o [23]),
    .ZN(_17139_));
 NAND2_X1 _43893_ (.A1(_17139_),
    .A2(_16018_),
    .ZN(_17140_));
 NAND3_X1 _43894_ (.A1(_17138_),
    .A2(_17140_),
    .A3(_15761_),
    .ZN(_17141_));
 INV_X1 _43895_ (.A(\icache.data_mems_3__data_mem.data_o [23]),
    .ZN(_17142_));
 NAND2_X1 _43896_ (.A1(_16580_),
    .A2(_17142_),
    .ZN(_17143_));
 INV_X16 _43897_ (.A(\icache.data_mems_2__data_mem.data_o [23]),
    .ZN(_17144_));
 NAND2_X2 _43898_ (.A1(_17144_),
    .A2(_16805_),
    .ZN(_17145_));
 NAND3_X1 _43899_ (.A1(_17143_),
    .A2(_17145_),
    .A3(_15754_),
    .ZN(_17146_));
 NAND3_X1 _43900_ (.A1(_17141_),
    .A2(_17146_),
    .A3(_15996_),
    .ZN(_17147_));
 NAND2_X2 _43901_ (.A1(_17137_),
    .A2(_17147_),
    .ZN(_17148_));
 OAI21_X1 _43902_ (.A(_17126_),
    .B1(_17148_),
    .B2(_16997_),
    .ZN(_05301_));
 BUF_X4 _43903_ (.A(_16724_),
    .Z(_17149_));
 NAND2_X1 _43904_ (.A1(_17149_),
    .A2(\icache.lce.lce_cmd_inst.data_r [472]),
    .ZN(_17150_));
 INV_X1 _43905_ (.A(\icache.data_mems_1__data_mem.data_o [24]),
    .ZN(_17151_));
 NAND2_X1 _43906_ (.A1(_15721_),
    .A2(_17151_),
    .ZN(_17152_));
 INV_X8 _43907_ (.A(\icache.data_mems_0__data_mem.data_o [24]),
    .ZN(_17153_));
 NAND2_X1 _43908_ (.A1(_17153_),
    .A2(_15479_),
    .ZN(_17154_));
 AOI21_X1 _43909_ (.A(_15567_),
    .B1(_17152_),
    .B2(_17154_),
    .ZN(_17155_));
 INV_X1 _43910_ (.A(\icache.data_mems_3__data_mem.data_o [24]),
    .ZN(_17156_));
 NAND2_X1 _43911_ (.A1(_15692_),
    .A2(_17156_),
    .ZN(_17157_));
 INV_X16 _43912_ (.A(\icache.data_mems_2__data_mem.data_o [24]),
    .ZN(_17158_));
 NAND2_X2 _43913_ (.A1(_17158_),
    .A2(_15752_),
    .ZN(_17159_));
 AOI21_X1 _43914_ (.A(_16005_),
    .B1(_17157_),
    .B2(_17159_),
    .ZN(_17160_));
 OAI21_X1 _43915_ (.A(_15735_),
    .B1(_17155_),
    .B2(_17160_),
    .ZN(_17161_));
 OR2_X1 _43916_ (.A1(_15967_),
    .A2(\icache.data_mems_7__data_mem.data_o [24]),
    .ZN(_17162_));
 INV_X8 _43917_ (.A(\icache.data_mems_6__data_mem.data_o [24]),
    .ZN(_17163_));
 NAND2_X2 _43918_ (.A1(_17163_),
    .A2(_15479_),
    .ZN(_17164_));
 NAND3_X2 _43919_ (.A1(_17162_),
    .A2(_17164_),
    .A3(_15754_),
    .ZN(_17165_));
 OR2_X1 _43920_ (.A1(_15906_),
    .A2(\icache.data_mems_5__data_mem.data_o [24]),
    .ZN(_17166_));
 INV_X1 _43921_ (.A(\icache.data_mems_4__data_mem.data_o [24]),
    .ZN(_17167_));
 NAND2_X1 _43922_ (.A1(_17167_),
    .A2(_15752_),
    .ZN(_17168_));
 NAND3_X1 _43923_ (.A1(_17166_),
    .A2(_17168_),
    .A3(_15761_),
    .ZN(_17169_));
 NAND3_X1 _43924_ (.A1(_17165_),
    .A2(_17169_),
    .A3(_15656_),
    .ZN(_17170_));
 NAND2_X2 _43925_ (.A1(_17161_),
    .A2(_17170_),
    .ZN(_17171_));
 OAI21_X1 _43926_ (.A(_17150_),
    .B1(_17171_),
    .B2(_16997_),
    .ZN(_05302_));
 NAND2_X1 _43927_ (.A1(_17149_),
    .A2(\icache.lce.lce_cmd_inst.data_r [473]),
    .ZN(_17172_));
 OR2_X1 _43928_ (.A1(_15751_),
    .A2(\icache.data_mems_7__data_mem.data_o [25]),
    .ZN(_17173_));
 INV_X4 _43929_ (.A(\icache.data_mems_6__data_mem.data_o [25]),
    .ZN(_17174_));
 NAND2_X1 _43930_ (.A1(_17174_),
    .A2(_16015_),
    .ZN(_17175_));
 NAND2_X1 _43931_ (.A1(_17173_),
    .A2(_17175_),
    .ZN(_17176_));
 NAND2_X1 _43932_ (.A1(_17176_),
    .A2(_16341_),
    .ZN(_17177_));
 INV_X1 _43933_ (.A(\icache.data_mems_5__data_mem.data_o [25]),
    .ZN(_17178_));
 NAND2_X1 _43934_ (.A1(_16343_),
    .A2(_17178_),
    .ZN(_17179_));
 INV_X1 _43935_ (.A(\icache.data_mems_4__data_mem.data_o [25]),
    .ZN(_17180_));
 NAND2_X1 _43936_ (.A1(_17180_),
    .A2(_15564_),
    .ZN(_17181_));
 NAND2_X1 _43937_ (.A1(_17179_),
    .A2(_17181_),
    .ZN(_17182_));
 NAND2_X1 _43938_ (.A1(_17182_),
    .A2(_16347_),
    .ZN(_17183_));
 NAND2_X2 _43939_ (.A1(_17177_),
    .A2(_17183_),
    .ZN(_17184_));
 NAND2_X1 _43940_ (.A1(_17184_),
    .A2(_16266_),
    .ZN(_17185_));
 INV_X1 _43941_ (.A(\icache.data_mems_1__data_mem.data_o [25]),
    .ZN(_17186_));
 NOR2_X1 _43942_ (.A1(_17186_),
    .A2(_16001_),
    .ZN(_17187_));
 AND2_X1 _43943_ (.A1(_15916_),
    .A2(\icache.data_mems_0__data_mem.data_o [25]),
    .ZN(_17188_));
 NOR3_X2 _43944_ (.A1(_17187_),
    .A2(_17188_),
    .A3(_15779_),
    .ZN(_17189_));
 OR2_X1 _43945_ (.A1(_16272_),
    .A2(\icache.data_mems_3__data_mem.data_o [25]),
    .ZN(_17190_));
 INV_X8 _43946_ (.A(\icache.data_mems_2__data_mem.data_o [25]),
    .ZN(_17191_));
 NAND2_X2 _43947_ (.A1(_17191_),
    .A2(_16805_),
    .ZN(_17192_));
 AOI21_X1 _43948_ (.A(_17016_),
    .B1(_17190_),
    .B2(_17192_),
    .ZN(_17193_));
 OAI21_X1 _43949_ (.A(_16237_),
    .B1(_17189_),
    .B2(_17193_),
    .ZN(_17194_));
 NAND2_X2 _43950_ (.A1(_17185_),
    .A2(_17194_),
    .ZN(_17195_));
 OAI21_X1 _43951_ (.A(_17172_),
    .B1(_17195_),
    .B2(_16997_),
    .ZN(_05303_));
 NAND2_X1 _43952_ (.A1(_17149_),
    .A2(\icache.lce.lce_cmd_inst.data_r [474]),
    .ZN(_17196_));
 AND2_X1 _43953_ (.A1(_15397_),
    .A2(\icache.data_mems_7__data_mem.data_o [26]),
    .ZN(_17197_));
 AND2_X1 _43954_ (.A1(_16319_),
    .A2(\icache.data_mems_6__data_mem.data_o [26]),
    .ZN(_17198_));
 OR3_X1 _43955_ (.A1(_17197_),
    .A2(_17198_),
    .A3(_17068_),
    .ZN(_17199_));
 NAND2_X1 _43956_ (.A1(_16394_),
    .A2(\icache.data_mems_4__data_mem.data_o [26]),
    .ZN(_17200_));
 INV_X2 _43957_ (.A(\icache.data_mems_5__data_mem.data_o [26]),
    .ZN(_17201_));
 OAI211_X2 _43958_ (.A(_17200_),
    .B(_16056_),
    .C1(_15728_),
    .C2(_17201_),
    .ZN(_17202_));
 NAND3_X1 _43959_ (.A1(_17199_),
    .A2(_16360_),
    .A3(_17202_),
    .ZN(_17203_));
 OR2_X1 _43960_ (.A1(_15411_),
    .A2(\icache.data_mems_3__data_mem.data_o [26]),
    .ZN(_17204_));
 INV_X8 _43961_ (.A(\icache.data_mems_2__data_mem.data_o [26]),
    .ZN(_17205_));
 NAND2_X1 _43962_ (.A1(_17205_),
    .A2(_15323_),
    .ZN(_17206_));
 NAND2_X2 _43963_ (.A1(_17204_),
    .A2(_17206_),
    .ZN(_17207_));
 NAND2_X1 _43964_ (.A1(_17207_),
    .A2(_15514_),
    .ZN(_17208_));
 INV_X1 _43965_ (.A(\icache.data_mems_1__data_mem.data_o [26]),
    .ZN(_17209_));
 NAND2_X1 _43966_ (.A1(_15417_),
    .A2(_17209_),
    .ZN(_17210_));
 INV_X1 _43967_ (.A(\icache.data_mems_0__data_mem.data_o [26]),
    .ZN(_17211_));
 NAND2_X1 _43968_ (.A1(_17211_),
    .A2(_15421_),
    .ZN(_17212_));
 NAND2_X1 _43969_ (.A1(_17210_),
    .A2(_17212_),
    .ZN(_17213_));
 NAND2_X1 _43970_ (.A1(_17213_),
    .A2(_16418_),
    .ZN(_17214_));
 NAND3_X1 _43971_ (.A1(_17208_),
    .A2(_17214_),
    .A3(_15315_),
    .ZN(_17215_));
 AND2_X4 _43972_ (.A1(_17203_),
    .A2(_17215_),
    .ZN(_17216_));
 BUF_X8 _43973_ (.A(_16785_),
    .Z(_17217_));
 OAI21_X1 _43974_ (.A(_17196_),
    .B1(_17216_),
    .B2(_17217_),
    .ZN(_05304_));
 NAND2_X1 _43975_ (.A1(_17149_),
    .A2(\icache.lce.lce_cmd_inst.data_r [475]),
    .ZN(_17218_));
 INV_X8 _43976_ (.A(\icache.data_mems_7__data_mem.data_o [27]),
    .ZN(_17219_));
 NOR2_X1 _43977_ (.A1(_17219_),
    .A2(_16001_),
    .ZN(_17220_));
 AND2_X1 _43978_ (.A1(_16224_),
    .A2(\icache.data_mems_6__data_mem.data_o [27]),
    .ZN(_17221_));
 OAI21_X2 _43979_ (.A(_15433_),
    .B1(_17220_),
    .B2(_17221_),
    .ZN(_17222_));
 OR2_X1 _43980_ (.A1(_15573_),
    .A2(\icache.data_mems_5__data_mem.data_o [27]),
    .ZN(_17223_));
 INV_X1 _43981_ (.A(\icache.data_mems_4__data_mem.data_o [27]),
    .ZN(_17224_));
 NAND2_X2 _43982_ (.A1(_17224_),
    .A2(_15752_),
    .ZN(_17225_));
 NAND3_X2 _43983_ (.A1(_17223_),
    .A2(_17225_),
    .A3(_15446_),
    .ZN(_17226_));
 AOI21_X1 _43984_ (.A(_15431_),
    .B1(_17222_),
    .B2(_17226_),
    .ZN(_17227_));
 BUF_X16 _43985_ (.A(_15369_),
    .Z(_17228_));
 INV_X1 _43986_ (.A(\icache.data_mems_1__data_mem.data_o [27]),
    .ZN(_17229_));
 NOR2_X1 _43987_ (.A1(_17229_),
    .A2(_15452_),
    .ZN(_17230_));
 AND2_X1 _43988_ (.A1(_15738_),
    .A2(\icache.data_mems_0__data_mem.data_o [27]),
    .ZN(_17231_));
 OAI21_X2 _43989_ (.A(_17228_),
    .B1(_17230_),
    .B2(_17231_),
    .ZN(_17232_));
 OR2_X1 _43990_ (.A1(_15457_),
    .A2(\icache.data_mems_3__data_mem.data_o [27]),
    .ZN(_17233_));
 INV_X8 _43991_ (.A(\icache.data_mems_2__data_mem.data_o [27]),
    .ZN(_17234_));
 NAND2_X2 _43992_ (.A1(_17234_),
    .A2(_16112_),
    .ZN(_17235_));
 BUF_X16 _43993_ (.A(_16229_),
    .Z(_17236_));
 NAND3_X2 _43994_ (.A1(_17233_),
    .A2(_17235_),
    .A3(_17236_),
    .ZN(_17237_));
 AOI21_X1 _43995_ (.A(_16714_),
    .B1(_17232_),
    .B2(_17237_),
    .ZN(_17238_));
 NOR2_X2 _43996_ (.A1(_17227_),
    .A2(_17238_),
    .ZN(_17239_));
 OAI21_X1 _43997_ (.A(_17218_),
    .B1(_17239_),
    .B2(_17217_),
    .ZN(_05305_));
 NAND2_X1 _43998_ (.A1(_17149_),
    .A2(\icache.lce.lce_cmd_inst.data_r [476]),
    .ZN(_17240_));
 AND2_X1 _43999_ (.A1(_16222_),
    .A2(\icache.data_mems_1__data_mem.data_o [28]),
    .ZN(_17241_));
 AND2_X1 _44000_ (.A1(_16253_),
    .A2(\icache.data_mems_0__data_mem.data_o [28]),
    .ZN(_17242_));
 OAI21_X2 _44001_ (.A(_15853_),
    .B1(_17241_),
    .B2(_17242_),
    .ZN(_17243_));
 INV_X1 _44002_ (.A(\icache.data_mems_3__data_mem.data_o [28]),
    .ZN(_17244_));
 NAND2_X2 _44003_ (.A1(_16035_),
    .A2(_17244_),
    .ZN(_17245_));
 INV_X8 _44004_ (.A(\icache.data_mems_2__data_mem.data_o [28]),
    .ZN(_17246_));
 NAND2_X2 _44005_ (.A1(_17246_),
    .A2(_15728_),
    .ZN(_17247_));
 NAND3_X2 _44006_ (.A1(_17245_),
    .A2(_17247_),
    .A3(_15911_),
    .ZN(_17248_));
 AOI21_X1 _44007_ (.A(_16956_),
    .B1(_17243_),
    .B2(_17248_),
    .ZN(_17249_));
 INV_X2 _44008_ (.A(\icache.data_mems_7__data_mem.data_o [28]),
    .ZN(_17250_));
 NOR2_X1 _44009_ (.A1(_17250_),
    .A2(_15335_),
    .ZN(_17251_));
 AND2_X1 _44010_ (.A1(_15346_),
    .A2(\icache.data_mems_6__data_mem.data_o [28]),
    .ZN(_17252_));
 OAI21_X2 _44011_ (.A(_16209_),
    .B1(_17251_),
    .B2(_17252_),
    .ZN(_17253_));
 INV_X1 _44012_ (.A(\icache.data_mems_5__data_mem.data_o [28]),
    .ZN(_17254_));
 NOR2_X1 _44013_ (.A1(_17254_),
    .A2(_15335_),
    .ZN(_17255_));
 AND2_X1 _44014_ (.A1(_15346_),
    .A2(\icache.data_mems_4__data_mem.data_o [28]),
    .ZN(_17256_));
 OAI21_X2 _44015_ (.A(_15553_),
    .B1(_17255_),
    .B2(_17256_),
    .ZN(_17257_));
 AOI21_X1 _44016_ (.A(_16564_),
    .B1(_17253_),
    .B2(_17257_),
    .ZN(_17258_));
 NOR2_X2 _44017_ (.A1(_17249_),
    .A2(_17258_),
    .ZN(_17259_));
 OAI21_X1 _44018_ (.A(_17240_),
    .B1(_17259_),
    .B2(_17217_),
    .ZN(_05306_));
 NAND2_X1 _44019_ (.A1(_17149_),
    .A2(\icache.lce.lce_cmd_inst.data_r [477]),
    .ZN(_17260_));
 NOR2_X1 _44020_ (.A1(_15908_),
    .A2(_15985_),
    .ZN(_17261_));
 AND2_X1 _44021_ (.A1(_15556_),
    .A2(\icache.data_mems_6__data_mem.data_o [29]),
    .ZN(_17262_));
 NOR2_X1 _44022_ (.A1(_17261_),
    .A2(_17262_),
    .ZN(_17263_));
 BUF_X16 _44023_ (.A(_16053_),
    .Z(_17264_));
 NOR2_X1 _44024_ (.A1(_17263_),
    .A2(_17264_),
    .ZN(_17265_));
 NAND2_X1 _44025_ (.A1(_15612_),
    .A2(\icache.data_mems_5__data_mem.data_o [29]),
    .ZN(_17266_));
 NAND2_X1 _44026_ (.A1(_16408_),
    .A2(\icache.data_mems_4__data_mem.data_o [29]),
    .ZN(_17267_));
 AOI21_X1 _44027_ (.A(_15432_),
    .B1(_17266_),
    .B2(_17267_),
    .ZN(_17268_));
 OAI21_X1 _44028_ (.A(_16631_),
    .B1(_17265_),
    .B2(_17268_),
    .ZN(_17269_));
 OR2_X1 _44029_ (.A1(_15411_),
    .A2(\icache.data_mems_3__data_mem.data_o [29]),
    .ZN(_17270_));
 NAND2_X1 _44030_ (.A1(_15914_),
    .A2(_15323_),
    .ZN(_17271_));
 NAND2_X1 _44031_ (.A1(_17270_),
    .A2(_17271_),
    .ZN(_17272_));
 BUF_X16 _44032_ (.A(_15311_),
    .Z(_17273_));
 NAND2_X1 _44033_ (.A1(_17272_),
    .A2(_17273_),
    .ZN(_17274_));
 NAND2_X1 _44034_ (.A1(_15417_),
    .A2(_15921_),
    .ZN(_17275_));
 NAND2_X1 _44035_ (.A1(_15919_),
    .A2(_15421_),
    .ZN(_17276_));
 NAND2_X1 _44036_ (.A1(_17275_),
    .A2(_17276_),
    .ZN(_17277_));
 NAND2_X1 _44037_ (.A1(_17277_),
    .A2(_16418_),
    .ZN(_17278_));
 NAND3_X1 _44038_ (.A1(_17274_),
    .A2(_17278_),
    .A3(_15315_),
    .ZN(_17279_));
 AND2_X4 _44039_ (.A1(_17269_),
    .A2(_17279_),
    .ZN(_17280_));
 OAI21_X1 _44040_ (.A(_17260_),
    .B1(_17280_),
    .B2(_17217_),
    .ZN(_05307_));
 NAND2_X1 _44041_ (.A1(_17149_),
    .A2(\icache.lce.lce_cmd_inst.data_r [478]),
    .ZN(_17281_));
 NOR2_X1 _44042_ (.A1(_15946_),
    .A2(_15460_),
    .ZN(_17282_));
 AND2_X1 _44043_ (.A1(_15876_),
    .A2(\icache.data_mems_0__data_mem.data_o [30]),
    .ZN(_17283_));
 NOR2_X2 _44044_ (.A1(_17282_),
    .A2(_17283_),
    .ZN(_17284_));
 NOR2_X1 _44045_ (.A1(_17284_),
    .A2(_15938_),
    .ZN(_17285_));
 NAND2_X2 _44046_ (.A1(_15836_),
    .A2(\icache.data_mems_3__data_mem.data_o [30]),
    .ZN(_17286_));
 NAND2_X2 _44047_ (.A1(_15511_),
    .A2(\icache.data_mems_2__data_mem.data_o [30]),
    .ZN(_17287_));
 AOI21_X2 _44048_ (.A(_15727_),
    .B1(_17286_),
    .B2(_17287_),
    .ZN(_17288_));
 NOR2_X4 _44049_ (.A1(_17285_),
    .A2(_17288_),
    .ZN(_17289_));
 NOR2_X1 _44050_ (.A1(_17289_),
    .A2(_16200_),
    .ZN(_17290_));
 NOR2_X4 _44051_ (.A1(_15935_),
    .A2(_16867_),
    .ZN(_17291_));
 AND2_X1 _44052_ (.A1(_15454_),
    .A2(\icache.data_mems_6__data_mem.data_o [30]),
    .ZN(_17292_));
 OAI21_X2 _44053_ (.A(_16209_),
    .B1(_17291_),
    .B2(_17292_),
    .ZN(_17293_));
 NOR2_X1 _44054_ (.A1(_15929_),
    .A2(_15335_),
    .ZN(_17294_));
 AND2_X1 _44055_ (.A1(_15346_),
    .A2(\icache.data_mems_4__data_mem.data_o [30]),
    .ZN(_17295_));
 OAI21_X2 _44056_ (.A(_15553_),
    .B1(_17294_),
    .B2(_17295_),
    .ZN(_17296_));
 AOI21_X1 _44057_ (.A(_16564_),
    .B1(_17293_),
    .B2(_17296_),
    .ZN(_17297_));
 NOR2_X2 _44058_ (.A1(_17290_),
    .A2(_17297_),
    .ZN(_17298_));
 OAI21_X1 _44059_ (.A(_17281_),
    .B1(_17298_),
    .B2(_17217_),
    .ZN(_05308_));
 NAND2_X1 _44060_ (.A1(_17149_),
    .A2(\icache.lce.lce_cmd_inst.data_r [479]),
    .ZN(_17299_));
 BUF_X16 _44061_ (.A(_15328_),
    .Z(_17300_));
 NOR2_X1 _44062_ (.A1(_15954_),
    .A2(_15452_),
    .ZN(_17301_));
 AND2_X1 _44063_ (.A1(_15738_),
    .A2(\icache.data_mems_4__data_mem.data_o [31]),
    .ZN(_17302_));
 OAI21_X2 _44064_ (.A(_15901_),
    .B1(_17301_),
    .B2(_17302_),
    .ZN(_17303_));
 NAND2_X1 _44065_ (.A1(_15627_),
    .A2(_15960_),
    .ZN(_17304_));
 NAND2_X2 _44066_ (.A1(_15958_),
    .A2(_16112_),
    .ZN(_17305_));
 NAND3_X2 _44067_ (.A1(_17304_),
    .A2(_17305_),
    .A3(_15911_),
    .ZN(_17306_));
 AOI21_X2 _44068_ (.A(_17300_),
    .B1(_17303_),
    .B2(_17306_),
    .ZN(_17307_));
 BUF_X16 _44069_ (.A(_15445_),
    .Z(_17308_));
 NOR2_X2 _44070_ (.A1(_15965_),
    .A2(_15452_),
    .ZN(_17309_));
 AND2_X1 _44071_ (.A1(_15738_),
    .A2(\icache.data_mems_0__data_mem.data_o [31]),
    .ZN(_17310_));
 OAI21_X2 _44072_ (.A(_17308_),
    .B1(_17309_),
    .B2(_17310_),
    .ZN(_17311_));
 INV_X1 _44073_ (.A(\icache.data_mems_3__data_mem.data_o [31]),
    .ZN(_17312_));
 NAND2_X2 _44074_ (.A1(_15627_),
    .A2(_17312_),
    .ZN(_17313_));
 NAND2_X1 _44075_ (.A1(_15969_),
    .A2(_16112_),
    .ZN(_17314_));
 NAND3_X2 _44076_ (.A1(_17313_),
    .A2(_17314_),
    .A3(_17236_),
    .ZN(_17315_));
 AOI21_X2 _44077_ (.A(_16714_),
    .B1(_17311_),
    .B2(_17315_),
    .ZN(_17316_));
 NOR2_X4 _44078_ (.A1(_17307_),
    .A2(_17316_),
    .ZN(_17317_));
 OAI21_X1 _44079_ (.A(_17299_),
    .B1(_17317_),
    .B2(_17217_),
    .ZN(_05309_));
 NAND2_X1 _44080_ (.A1(_17149_),
    .A2(\icache.lce.lce_cmd_inst.data_r [480]),
    .ZN(_17318_));
 NOR2_X1 _44081_ (.A1(_15978_),
    .A2(_15985_),
    .ZN(_17319_));
 AND2_X1 _44082_ (.A1(_15550_),
    .A2(\icache.data_mems_4__data_mem.data_o [32]),
    .ZN(_17320_));
 NOR2_X1 _44083_ (.A1(_17319_),
    .A2(_17320_),
    .ZN(_17321_));
 NOR2_X1 _44084_ (.A1(_17321_),
    .A2(_15425_),
    .ZN(_17322_));
 NAND2_X1 _44085_ (.A1(_15612_),
    .A2(\icache.data_mems_7__data_mem.data_o [32]),
    .ZN(_17323_));
 NAND2_X1 _44086_ (.A1(_16408_),
    .A2(\icache.data_mems_6__data_mem.data_o [32]),
    .ZN(_17324_));
 AOI21_X1 _44087_ (.A(_15660_),
    .B1(_17323_),
    .B2(_17324_),
    .ZN(_17325_));
 NOR3_X1 _44088_ (.A1(_17322_),
    .A2(_15724_),
    .A3(_17325_),
    .ZN(_17326_));
 NAND2_X1 _44089_ (.A1(_15417_),
    .A2(_15992_),
    .ZN(_17327_));
 NAND2_X1 _44090_ (.A1(_15990_),
    .A2(_15421_),
    .ZN(_17328_));
 NAND2_X2 _44091_ (.A1(_17327_),
    .A2(_17328_),
    .ZN(_17329_));
 NAND2_X1 _44092_ (.A1(_17329_),
    .A2(_16195_),
    .ZN(_17330_));
 NAND2_X1 _44093_ (.A1(_15417_),
    .A2(_15984_),
    .ZN(_17331_));
 NAND2_X1 _44094_ (.A1(_15982_),
    .A2(_15478_),
    .ZN(_17332_));
 NAND2_X2 _44095_ (.A1(_17331_),
    .A2(_17332_),
    .ZN(_17333_));
 NAND2_X1 _44096_ (.A1(_17333_),
    .A2(_16541_),
    .ZN(_17334_));
 AOI21_X1 _44097_ (.A(_15670_),
    .B1(_17330_),
    .B2(_17334_),
    .ZN(_17335_));
 OR2_X2 _44098_ (.A1(_17326_),
    .A2(_17335_),
    .ZN(_17336_));
 OAI21_X1 _44099_ (.A(_17318_),
    .B1(_17336_),
    .B2(_17217_),
    .ZN(_05311_));
 NAND2_X1 _44100_ (.A1(_17149_),
    .A2(\icache.lce.lce_cmd_inst.data_r [481]),
    .ZN(_17337_));
 NOR2_X1 _44101_ (.A1(_16007_),
    .A2(_15505_),
    .ZN(_17338_));
 AND2_X1 _44102_ (.A1(_15390_),
    .A2(\icache.data_mems_2__data_mem.data_o [33]),
    .ZN(_17339_));
 OR3_X2 _44103_ (.A1(_17338_),
    .A2(_17339_),
    .A3(_16053_),
    .ZN(_17340_));
 OR2_X1 _44104_ (.A1(_15411_),
    .A2(\icache.data_mems_1__data_mem.data_o [33]),
    .ZN(_17341_));
 NAND2_X1 _44105_ (.A1(_16000_),
    .A2(_15511_),
    .ZN(_17342_));
 NAND2_X1 _44106_ (.A1(_17341_),
    .A2(_17342_),
    .ZN(_17343_));
 NAND2_X1 _44107_ (.A1(_17343_),
    .A2(_15406_),
    .ZN(_17344_));
 AOI21_X2 _44108_ (.A(_16049_),
    .B1(_17340_),
    .B2(_17344_),
    .ZN(_17345_));
 NOR2_X1 _44109_ (.A1(_16017_),
    .A2(_15518_),
    .ZN(_17346_));
 AND2_X1 _44110_ (.A1(_16061_),
    .A2(\icache.data_mems_4__data_mem.data_o [33]),
    .ZN(_17347_));
 OAI21_X1 _44111_ (.A(_15484_),
    .B1(_17346_),
    .B2(_17347_),
    .ZN(_17348_));
 NAND2_X1 _44112_ (.A1(_15523_),
    .A2(_16024_),
    .ZN(_17349_));
 NAND2_X1 _44113_ (.A1(_16022_),
    .A2(_15495_),
    .ZN(_17350_));
 NAND3_X1 _44114_ (.A1(_17349_),
    .A2(_17350_),
    .A3(_15378_),
    .ZN(_17351_));
 AND3_X1 _44115_ (.A1(_17348_),
    .A2(_15522_),
    .A3(_17351_),
    .ZN(_17352_));
 OR2_X4 _44116_ (.A1(_17345_),
    .A2(_17352_),
    .ZN(_17353_));
 OAI21_X1 _44117_ (.A(_17337_),
    .B1(_17353_),
    .B2(_17217_),
    .ZN(_05312_));
 BUF_X8 _44118_ (.A(_16724_),
    .Z(_17354_));
 NAND2_X1 _44119_ (.A1(_17354_),
    .A2(\icache.lce.lce_cmd_inst.data_r [482]),
    .ZN(_17355_));
 NOR2_X1 _44120_ (.A1(_15523_),
    .A2(\icache.data_mems_6__data_mem.data_o [34]),
    .ZN(_17356_));
 AOI211_X2 _44121_ (.A(_15463_),
    .B(_17356_),
    .C1(_15679_),
    .C2(_16036_),
    .ZN(_17357_));
 NAND2_X1 _44122_ (.A1(_15612_),
    .A2(\icache.data_mems_5__data_mem.data_o [34]),
    .ZN(_17358_));
 NAND2_X1 _44123_ (.A1(_15346_),
    .A2(\icache.data_mems_4__data_mem.data_o [34]),
    .ZN(_17359_));
 AOI21_X1 _44124_ (.A(_16643_),
    .B1(_17358_),
    .B2(_17359_),
    .ZN(_17360_));
 NOR3_X1 _44125_ (.A1(_17357_),
    .A2(_15724_),
    .A3(_17360_),
    .ZN(_17361_));
 NAND2_X1 _44126_ (.A1(_16343_),
    .A2(\icache.data_mems_3__data_mem.data_o [34]),
    .ZN(_17362_));
 OAI211_X2 _44127_ (.A(_17362_),
    .B(_15678_),
    .C1(_15679_),
    .C2(_16042_),
    .ZN(_17363_));
 NAND2_X1 _44128_ (.A1(_15736_),
    .A2(\icache.data_mems_1__data_mem.data_o [34]),
    .ZN(_17364_));
 NAND2_X1 _44129_ (.A1(_15916_),
    .A2(\icache.data_mems_0__data_mem.data_o [34]),
    .ZN(_17365_));
 NAND3_X2 _44130_ (.A1(_17364_),
    .A2(_15673_),
    .A3(_17365_),
    .ZN(_17366_));
 AOI21_X1 _44131_ (.A(_15670_),
    .B1(_17363_),
    .B2(_17366_),
    .ZN(_17367_));
 OR2_X4 _44132_ (.A1(_17361_),
    .A2(_17367_),
    .ZN(_17368_));
 OAI21_X1 _44133_ (.A(_17355_),
    .B1(_17368_),
    .B2(_17217_),
    .ZN(_05313_));
 NAND2_X1 _44134_ (.A1(_17354_),
    .A2(\icache.lce.lce_cmd_inst.data_r [483]),
    .ZN(_17369_));
 OR2_X1 _44135_ (.A1(_15714_),
    .A2(\icache.data_mems_3__data_mem.data_o [35]),
    .ZN(_17370_));
 NAND2_X1 _44136_ (.A1(_16050_),
    .A2(_16408_),
    .ZN(_17371_));
 NAND2_X2 _44137_ (.A1(_17370_),
    .A2(_17371_),
    .ZN(_17372_));
 NAND2_X1 _44138_ (.A1(_17372_),
    .A2(_16341_),
    .ZN(_17373_));
 NAND2_X1 _44139_ (.A1(_15398_),
    .A2(_16057_),
    .ZN(_17374_));
 INV_X1 _44140_ (.A(\icache.data_mems_0__data_mem.data_o [35]),
    .ZN(_17375_));
 NAND2_X1 _44141_ (.A1(_17375_),
    .A2(_15402_),
    .ZN(_17376_));
 NAND2_X4 _44142_ (.A1(_17374_),
    .A2(_17376_),
    .ZN(_17377_));
 NAND2_X1 _44143_ (.A1(_17377_),
    .A2(_16347_),
    .ZN(_17378_));
 NAND2_X1 _44144_ (.A1(_17373_),
    .A2(_17378_),
    .ZN(_17379_));
 NAND2_X1 _44145_ (.A1(_17379_),
    .A2(_15580_),
    .ZN(_17380_));
 NAND2_X1 _44146_ (.A1(_15491_),
    .A2(_16066_),
    .ZN(_17381_));
 NAND2_X1 _44147_ (.A1(_16064_),
    .A2(_15985_),
    .ZN(_17382_));
 AND3_X1 _44148_ (.A1(_17381_),
    .A2(_17382_),
    .A3(_15463_),
    .ZN(_17383_));
 NAND2_X2 _44149_ (.A1(_15772_),
    .A2(\icache.data_mems_7__data_mem.data_o [35]),
    .ZN(_17384_));
 NAND2_X2 _44150_ (.A1(_15338_),
    .A2(\icache.data_mems_6__data_mem.data_o [35]),
    .ZN(_17385_));
 AOI21_X2 _44151_ (.A(_15484_),
    .B1(_17384_),
    .B2(_17385_),
    .ZN(_17386_));
 OR3_X2 _44152_ (.A1(_17383_),
    .A2(_17386_),
    .A3(_15699_),
    .ZN(_17387_));
 NAND2_X4 _44153_ (.A1(_17380_),
    .A2(_17387_),
    .ZN(_17388_));
 OAI21_X1 _44154_ (.A(_17369_),
    .B1(_17388_),
    .B2(_17217_),
    .ZN(_05314_));
 NAND2_X1 _44155_ (.A1(_17354_),
    .A2(\icache.lce.lce_cmd_inst.data_r [484]),
    .ZN(_17389_));
 NOR2_X1 _44156_ (.A1(_16074_),
    .A2(_15359_),
    .ZN(_17390_));
 AND2_X1 _44157_ (.A1(_16319_),
    .A2(\icache.data_mems_0__data_mem.data_o [36]),
    .ZN(_17391_));
 OR3_X2 _44158_ (.A1(_17390_),
    .A2(_17391_),
    .A3(_16321_),
    .ZN(_17392_));
 NAND2_X1 _44159_ (.A1(_15475_),
    .A2(\icache.data_mems_2__data_mem.data_o [36]),
    .ZN(_17393_));
 OAI211_X2 _44160_ (.A(_17393_),
    .B(_16324_),
    .C1(_15479_),
    .C2(_16079_),
    .ZN(_17394_));
 AND3_X1 _44161_ (.A1(_17392_),
    .A2(_15474_),
    .A3(_17394_),
    .ZN(_17395_));
 NOR2_X1 _44162_ (.A1(_16085_),
    .A2(_15505_),
    .ZN(_17396_));
 AND2_X1 _44163_ (.A1(_15700_),
    .A2(\icache.data_mems_6__data_mem.data_o [36]),
    .ZN(_17397_));
 OAI21_X2 _44164_ (.A(_16327_),
    .B1(_17396_),
    .B2(_17397_),
    .ZN(_17398_));
 NAND2_X1 _44165_ (.A1(_15491_),
    .A2(_16090_),
    .ZN(_17399_));
 NAND2_X1 _44166_ (.A1(_16088_),
    .A2(_16067_),
    .ZN(_17400_));
 NAND3_X1 _44167_ (.A1(_17399_),
    .A2(_17400_),
    .A3(_15342_),
    .ZN(_17401_));
 AOI21_X2 _44168_ (.A(_16564_),
    .B1(_17398_),
    .B2(_17401_),
    .ZN(_17402_));
 NOR2_X4 _44169_ (.A1(_17395_),
    .A2(_17402_),
    .ZN(_17403_));
 BUF_X8 _44170_ (.A(_16785_),
    .Z(_17404_));
 OAI21_X1 _44171_ (.A(_17389_),
    .B1(_17403_),
    .B2(_17404_),
    .ZN(_05315_));
 NAND2_X1 _44172_ (.A1(_17354_),
    .A2(\icache.lce.lce_cmd_inst.data_r [485]),
    .ZN(_17405_));
 OR2_X2 _44173_ (.A1(_15460_),
    .A2(\icache.data_mems_3__data_mem.data_o [37]),
    .ZN(_17406_));
 NAND2_X1 _44174_ (.A1(_16105_),
    .A2(_16253_),
    .ZN(_17407_));
 NAND2_X1 _44175_ (.A1(_17406_),
    .A2(_17407_),
    .ZN(_17408_));
 NAND2_X1 _44176_ (.A1(_17408_),
    .A2(_15911_),
    .ZN(_17409_));
 NAND2_X1 _44177_ (.A1(_15569_),
    .A2(_16111_),
    .ZN(_17410_));
 NAND2_X1 _44178_ (.A1(_16109_),
    .A2(_15573_),
    .ZN(_17411_));
 NAND2_X2 _44179_ (.A1(_17410_),
    .A2(_17411_),
    .ZN(_17412_));
 NAND2_X1 _44180_ (.A1(_17412_),
    .A2(_15576_),
    .ZN(_17413_));
 NAND3_X1 _44181_ (.A1(_17409_),
    .A2(_17413_),
    .A3(_15834_),
    .ZN(_17414_));
 BUF_X8 _44182_ (.A(_15408_),
    .Z(_17415_));
 OR2_X1 _44183_ (.A1(_15334_),
    .A2(\icache.data_mems_7__data_mem.data_o [37]),
    .ZN(_17416_));
 NAND2_X1 _44184_ (.A1(_16100_),
    .A2(_15955_),
    .ZN(_17417_));
 AND3_X1 _44185_ (.A1(_17416_),
    .A2(_17417_),
    .A3(_16643_),
    .ZN(_17418_));
 NAND2_X1 _44186_ (.A1(_16391_),
    .A2(\icache.data_mems_5__data_mem.data_o [37]),
    .ZN(_17419_));
 NAND2_X1 _44187_ (.A1(_15475_),
    .A2(\icache.data_mems_4__data_mem.data_o [37]),
    .ZN(_17420_));
 AOI21_X1 _44188_ (.A(_16324_),
    .B1(_17419_),
    .B2(_17420_),
    .ZN(_17421_));
 OAI21_X1 _44189_ (.A(_17415_),
    .B1(_17418_),
    .B2(_17421_),
    .ZN(_17422_));
 AND2_X2 _44190_ (.A1(_17414_),
    .A2(_17422_),
    .ZN(_17423_));
 OAI21_X1 _44191_ (.A(_17405_),
    .B1(_17423_),
    .B2(_17404_),
    .ZN(_05316_));
 NAND2_X1 _44192_ (.A1(_17354_),
    .A2(\icache.lce.lce_cmd_inst.data_r [486]),
    .ZN(_17424_));
 NOR2_X1 _44193_ (.A1(_16123_),
    .A2(_15985_),
    .ZN(_17425_));
 AND2_X1 _44194_ (.A1(_15550_),
    .A2(\icache.data_mems_6__data_mem.data_o [38]),
    .ZN(_17426_));
 NOR2_X2 _44195_ (.A1(_17425_),
    .A2(_17426_),
    .ZN(_17427_));
 NOR2_X1 _44196_ (.A1(_17427_),
    .A2(_17264_),
    .ZN(_17428_));
 NAND2_X1 _44197_ (.A1(_15612_),
    .A2(\icache.data_mems_5__data_mem.data_o [38]),
    .ZN(_17429_));
 NAND2_X1 _44198_ (.A1(_16408_),
    .A2(\icache.data_mems_4__data_mem.data_o [38]),
    .ZN(_17430_));
 AOI21_X2 _44199_ (.A(_16643_),
    .B1(_17429_),
    .B2(_17430_),
    .ZN(_17431_));
 NOR3_X1 _44200_ (.A1(_17428_),
    .A2(_15724_),
    .A3(_17431_),
    .ZN(_17432_));
 OR2_X1 _44201_ (.A1(_15556_),
    .A2(\icache.data_mems_1__data_mem.data_o [38]),
    .ZN(_17433_));
 NAND2_X1 _44202_ (.A1(_16129_),
    .A2(_15323_),
    .ZN(_17434_));
 NAND2_X4 _44203_ (.A1(_17433_),
    .A2(_17434_),
    .ZN(_17435_));
 NAND2_X1 _44204_ (.A1(_17435_),
    .A2(_16195_),
    .ZN(_17436_));
 NAND2_X1 _44205_ (.A1(_16343_),
    .A2(\icache.data_mems_3__data_mem.data_o [38]),
    .ZN(_17437_));
 NAND2_X1 _44206_ (.A1(_16083_),
    .A2(\icache.data_mems_2__data_mem.data_o [38]),
    .ZN(_17438_));
 NAND3_X1 _44207_ (.A1(_17437_),
    .A2(_15321_),
    .A3(_17438_),
    .ZN(_17439_));
 AOI21_X1 _44208_ (.A(_15670_),
    .B1(_17436_),
    .B2(_17439_),
    .ZN(_17440_));
 OR2_X2 _44209_ (.A1(_17432_),
    .A2(_17440_),
    .ZN(_17441_));
 OAI21_X1 _44210_ (.A(_17424_),
    .B1(_17441_),
    .B2(_17404_),
    .ZN(_05317_));
 NAND2_X1 _44211_ (.A1(_17354_),
    .A2(\icache.lce.lce_cmd_inst.data_r [487]),
    .ZN(_17442_));
 NOR2_X1 _44212_ (.A1(_15537_),
    .A2(\icache.data_mems_0__data_mem.data_o [39]),
    .ZN(_17443_));
 AOI211_X2 _44213_ (.A(_15497_),
    .B(_17443_),
    .C1(_16035_),
    .C2(_16149_),
    .ZN(_17444_));
 NAND2_X1 _44214_ (.A1(_15719_),
    .A2(\icache.data_mems_3__data_mem.data_o [39]),
    .ZN(_17445_));
 NAND2_X1 _44215_ (.A1(_15967_),
    .A2(\icache.data_mems_2__data_mem.data_o [39]),
    .ZN(_17446_));
 AOI21_X1 _44216_ (.A(_15673_),
    .B1(_17445_),
    .B2(_17446_),
    .ZN(_17447_));
 OAI21_X1 _44217_ (.A(_16438_),
    .B1(_17444_),
    .B2(_17447_),
    .ZN(_17448_));
 OR2_X1 _44218_ (.A1(_15714_),
    .A2(\icache.data_mems_5__data_mem.data_o [39]),
    .ZN(_17449_));
 NAND2_X1 _44219_ (.A1(_16139_),
    .A2(_16408_),
    .ZN(_17450_));
 NAND2_X1 _44220_ (.A1(_17449_),
    .A2(_17450_),
    .ZN(_17451_));
 NAND2_X1 _44221_ (.A1(_17451_),
    .A2(_15343_),
    .ZN(_17452_));
 NAND2_X1 _44222_ (.A1(_16391_),
    .A2(\icache.data_mems_7__data_mem.data_o [39]),
    .ZN(_17453_));
 NAND2_X2 _44223_ (.A1(_16394_),
    .A2(\icache.data_mems_6__data_mem.data_o [39]),
    .ZN(_17454_));
 NAND3_X2 _44224_ (.A1(_17453_),
    .A2(_15514_),
    .A3(_17454_),
    .ZN(_17455_));
 NAND3_X1 _44225_ (.A1(_17452_),
    .A2(_15409_),
    .A3(_17455_),
    .ZN(_17456_));
 AND2_X1 _44226_ (.A1(_17448_),
    .A2(_17456_),
    .ZN(_17457_));
 OAI21_X1 _44227_ (.A(_17442_),
    .B1(_17457_),
    .B2(_17404_),
    .ZN(_05318_));
 NAND2_X1 _44228_ (.A1(_17354_),
    .A2(\icache.lce.lce_cmd_inst.data_r [488]),
    .ZN(_17458_));
 BUF_X16 _44229_ (.A(_15483_),
    .Z(_17459_));
 NAND2_X1 _44230_ (.A1(_15671_),
    .A2(\icache.data_mems_7__data_mem.data_o [40]),
    .ZN(_17460_));
 NAND2_X1 _44231_ (.A1(_15725_),
    .A2(\icache.data_mems_6__data_mem.data_o [40]),
    .ZN(_17461_));
 AOI21_X2 _44232_ (.A(_17459_),
    .B1(_17460_),
    .B2(_17461_),
    .ZN(_17462_));
 NAND2_X1 _44233_ (.A1(_15719_),
    .A2(\icache.data_mems_5__data_mem.data_o [40]),
    .ZN(_17463_));
 NAND2_X1 _44234_ (.A1(_15475_),
    .A2(\icache.data_mems_4__data_mem.data_o [40]),
    .ZN(_17464_));
 AOI21_X1 _44235_ (.A(_15477_),
    .B1(_17463_),
    .B2(_17464_),
    .ZN(_17465_));
 OAI21_X1 _44236_ (.A(_16631_),
    .B1(_17462_),
    .B2(_17465_),
    .ZN(_17466_));
 NAND2_X1 _44237_ (.A1(_15719_),
    .A2(\icache.data_mems_3__data_mem.data_o [40]),
    .ZN(_17467_));
 NAND2_X1 _44238_ (.A1(_15967_),
    .A2(\icache.data_mems_2__data_mem.data_o [40]),
    .ZN(_17468_));
 NAND3_X1 _44239_ (.A1(_17467_),
    .A2(_15395_),
    .A3(_17468_),
    .ZN(_17469_));
 NAND2_X1 _44240_ (.A1(_16169_),
    .A2(\icache.data_mems_0__data_mem.data_o [40]),
    .ZN(_17470_));
 OAI211_X4 _44241_ (.A(_17470_),
    .B(_17459_),
    .C1(_15324_),
    .C2(_16168_),
    .ZN(_17471_));
 NAND3_X1 _44242_ (.A1(_17469_),
    .A2(_16372_),
    .A3(_17471_),
    .ZN(_17472_));
 AND2_X4 _44243_ (.A1(_17466_),
    .A2(_17472_),
    .ZN(_17473_));
 OAI21_X1 _44244_ (.A(_17458_),
    .B1(_17473_),
    .B2(_17404_),
    .ZN(_05319_));
 NAND2_X1 _44245_ (.A1(_17354_),
    .A2(\icache.lce.lce_cmd_inst.data_r [489]),
    .ZN(_17474_));
 NOR2_X2 _44246_ (.A1(_16186_),
    .A2(_15533_),
    .ZN(_17475_));
 AND2_X1 _44247_ (.A1(_15471_),
    .A2(\icache.data_mems_2__data_mem.data_o [41]),
    .ZN(_17476_));
 OAI21_X2 _44248_ (.A(_15432_),
    .B1(_17475_),
    .B2(_17476_),
    .ZN(_17477_));
 NAND2_X2 _44249_ (.A1(_15554_),
    .A2(_16192_),
    .ZN(_17478_));
 NAND2_X2 _44250_ (.A1(_16190_),
    .A2(_15714_),
    .ZN(_17479_));
 NAND3_X4 _44251_ (.A1(_17478_),
    .A2(_17479_),
    .A3(_15369_),
    .ZN(_17480_));
 AND3_X1 _44252_ (.A1(_17477_),
    .A2(_15699_),
    .A3(_17480_),
    .ZN(_17481_));
 NAND2_X1 _44253_ (.A1(_15398_),
    .A2(\icache.data_mems_5__data_mem.data_o [41]),
    .ZN(_17482_));
 NAND2_X1 _44254_ (.A1(_15955_),
    .A2(\icache.data_mems_4__data_mem.data_o [41]),
    .ZN(_17483_));
 NAND3_X1 _44255_ (.A1(_17482_),
    .A2(_17459_),
    .A3(_17483_),
    .ZN(_17484_));
 NAND2_X1 _44256_ (.A1(_16253_),
    .A2(\icache.data_mems_6__data_mem.data_o [41]),
    .ZN(_17485_));
 OAI211_X4 _44257_ (.A(_17485_),
    .B(_15678_),
    .C1(_15909_),
    .C2(_16181_),
    .ZN(_17486_));
 AOI21_X1 _44258_ (.A(_15579_),
    .B1(_17484_),
    .B2(_17486_),
    .ZN(_17487_));
 OR2_X2 _44259_ (.A1(_17481_),
    .A2(_17487_),
    .ZN(_17488_));
 OAI21_X1 _44260_ (.A(_17474_),
    .B1(_17488_),
    .B2(_17404_),
    .ZN(_05320_));
 NAND2_X1 _44261_ (.A1(_17354_),
    .A2(\icache.lce.lce_cmd_inst.data_r [507]),
    .ZN(_17489_));
 OR2_X1 _44262_ (.A1(_15317_),
    .A2(\icache.data_mems_5__data_mem.data_o [59]),
    .ZN(_17490_));
 NAND2_X1 _44263_ (.A1(_16569_),
    .A2(_15955_),
    .ZN(_17491_));
 NAND2_X1 _44264_ (.A1(_17490_),
    .A2(_17491_),
    .ZN(_17492_));
 NAND2_X1 _44265_ (.A1(_17492_),
    .A2(_16256_),
    .ZN(_17493_));
 OR2_X1 _44266_ (.A1(_15387_),
    .A2(\icache.data_mems_7__data_mem.data_o [59]),
    .ZN(_17494_));
 NAND2_X1 _44267_ (.A1(_16565_),
    .A2(_15391_),
    .ZN(_17495_));
 NAND2_X1 _44268_ (.A1(_17494_),
    .A2(_17495_),
    .ZN(_17496_));
 NAND2_X1 _44269_ (.A1(_17496_),
    .A2(_16262_),
    .ZN(_17497_));
 NAND2_X1 _44270_ (.A1(_17493_),
    .A2(_17497_),
    .ZN(_17498_));
 NAND2_X1 _44271_ (.A1(_17498_),
    .A2(_16266_),
    .ZN(_17499_));
 BUF_X16 _44272_ (.A(_15644_),
    .Z(_17500_));
 NOR2_X1 _44273_ (.A1(_16552_),
    .A2(_15505_),
    .ZN(_17501_));
 AND2_X1 _44274_ (.A1(_15700_),
    .A2(\icache.data_mems_0__data_mem.data_o [59]),
    .ZN(_17502_));
 NOR3_X2 _44275_ (.A1(_17501_),
    .A2(_17502_),
    .A3(_15779_),
    .ZN(_17503_));
 NAND2_X1 _44276_ (.A1(_15491_),
    .A2(_16558_),
    .ZN(_17504_));
 NAND2_X1 _44277_ (.A1(_16556_),
    .A2(_16067_),
    .ZN(_17505_));
 AOI21_X2 _44278_ (.A(_17016_),
    .B1(_17504_),
    .B2(_17505_),
    .ZN(_17506_));
 OAI21_X4 _44279_ (.A(_17500_),
    .B1(_17503_),
    .B2(_17506_),
    .ZN(_17507_));
 NAND2_X4 _44280_ (.A1(_17499_),
    .A2(_17507_),
    .ZN(_17508_));
 OAI21_X1 _44281_ (.A(_17489_),
    .B1(_17508_),
    .B2(_17404_),
    .ZN(_05341_));
 NAND2_X1 _44282_ (.A1(_17354_),
    .A2(\icache.lce.lce_cmd_inst.data_r [490]),
    .ZN(_17509_));
 NAND2_X1 _44283_ (.A1(_16155_),
    .A2(\icache.data_mems_3__data_mem.data_o [42]),
    .ZN(_17510_));
 BUF_X8 _44284_ (.A(_15320_),
    .Z(_17511_));
 OAI211_X1 _44285_ (.A(_17510_),
    .B(_17511_),
    .C1(_15721_),
    .C2(_16204_),
    .ZN(_17512_));
 NAND2_X1 _44286_ (.A1(_16343_),
    .A2(\icache.data_mems_1__data_mem.data_o [42]),
    .ZN(_17513_));
 NAND2_X1 _44287_ (.A1(_16015_),
    .A2(\icache.data_mems_0__data_mem.data_o [42]),
    .ZN(_17514_));
 NAND3_X1 _44288_ (.A1(_17513_),
    .A2(_17264_),
    .A3(_17514_),
    .ZN(_17515_));
 AND3_X1 _44289_ (.A1(_17512_),
    .A2(_15474_),
    .A3(_17515_),
    .ZN(_17516_));
 BUF_X16 _44290_ (.A(_15328_),
    .Z(_17517_));
 NOR2_X1 _44291_ (.A1(_16215_),
    .A2(_16867_),
    .ZN(_17518_));
 AND2_X1 _44292_ (.A1(_15916_),
    .A2(\icache.data_mems_4__data_mem.data_o [42]),
    .ZN(_17519_));
 OAI21_X2 _44293_ (.A(_16865_),
    .B1(_17518_),
    .B2(_17519_),
    .ZN(_17520_));
 OR2_X1 _44294_ (.A1(_16272_),
    .A2(\icache.data_mems_7__data_mem.data_o [42]),
    .ZN(_17521_));
 NAND2_X1 _44295_ (.A1(_16210_),
    .A2(_16805_),
    .ZN(_17522_));
 NAND3_X2 _44296_ (.A1(_17521_),
    .A2(_17522_),
    .A3(_16583_),
    .ZN(_17523_));
 AOI21_X2 _44297_ (.A(_17517_),
    .B1(_17520_),
    .B2(_17523_),
    .ZN(_17524_));
 NOR2_X4 _44298_ (.A1(_17516_),
    .A2(_17524_),
    .ZN(_17525_));
 OAI21_X1 _44299_ (.A(_17509_),
    .B1(_17525_),
    .B2(_17404_),
    .ZN(_05322_));
 BUF_X16 _44300_ (.A(_16724_),
    .Z(_17526_));
 NAND2_X1 _44301_ (.A1(_17526_),
    .A2(\icache.lce.lce_cmd_inst.data_r [491]),
    .ZN(_17527_));
 NAND2_X1 _44302_ (.A1(_15569_),
    .A2(_16240_),
    .ZN(_17528_));
 NAND2_X1 _44303_ (.A1(_16238_),
    .A2(_15573_),
    .ZN(_17529_));
 NAND2_X2 _44304_ (.A1(_17528_),
    .A2(_17529_),
    .ZN(_17530_));
 NAND2_X1 _44305_ (.A1(_17530_),
    .A2(_16256_),
    .ZN(_17531_));
 NAND2_X2 _44306_ (.A1(_15569_),
    .A2(_16245_),
    .ZN(_17532_));
 NAND2_X1 _44307_ (.A1(_16243_),
    .A2(_15564_),
    .ZN(_17533_));
 NAND2_X1 _44308_ (.A1(_17532_),
    .A2(_17533_),
    .ZN(_17534_));
 NAND2_X1 _44309_ (.A1(_17534_),
    .A2(_16262_),
    .ZN(_17535_));
 NAND2_X1 _44310_ (.A1(_17531_),
    .A2(_17535_),
    .ZN(_17536_));
 NAND2_X1 _44311_ (.A1(_17536_),
    .A2(_15580_),
    .ZN(_17537_));
 NAND2_X1 _44312_ (.A1(_16391_),
    .A2(\icache.data_mems_7__data_mem.data_o [43]),
    .ZN(_17538_));
 NAND2_X1 _44313_ (.A1(_15475_),
    .A2(\icache.data_mems_6__data_mem.data_o [43]),
    .ZN(_17539_));
 AND3_X1 _44314_ (.A1(_17538_),
    .A2(_16541_),
    .A3(_17539_),
    .ZN(_17540_));
 NAND2_X1 _44315_ (.A1(_15772_),
    .A2(_16233_),
    .ZN(_17541_));
 NAND2_X1 _44316_ (.A1(_16231_),
    .A2(_15955_),
    .ZN(_17542_));
 AOI21_X2 _44317_ (.A(_16544_),
    .B1(_17541_),
    .B2(_17542_),
    .ZN(_17543_));
 OAI21_X2 _44318_ (.A(_16013_),
    .B1(_17540_),
    .B2(_17543_),
    .ZN(_17544_));
 NAND2_X4 _44319_ (.A1(_17537_),
    .A2(_17544_),
    .ZN(_17545_));
 OAI21_X1 _44320_ (.A(_17527_),
    .B1(_17545_),
    .B2(_17404_),
    .ZN(_05323_));
 NAND2_X1 _44321_ (.A1(_17526_),
    .A2(\icache.lce.lce_cmd_inst.data_r [492]),
    .ZN(_17546_));
 NOR2_X1 _44322_ (.A1(_16259_),
    .A2(_15359_),
    .ZN(_17547_));
 AND2_X1 _44323_ (.A1(_16319_),
    .A2(\icache.data_mems_6__data_mem.data_o [44]),
    .ZN(_17548_));
 OAI21_X2 _44324_ (.A(_16209_),
    .B1(_17547_),
    .B2(_17548_),
    .ZN(_17549_));
 NOR2_X1 _44325_ (.A1(_16252_),
    .A2(_15334_),
    .ZN(_17550_));
 AND2_X1 _44326_ (.A1(_15322_),
    .A2(\icache.data_mems_4__data_mem.data_o [44]),
    .ZN(_17551_));
 OAI21_X2 _44327_ (.A(_15553_),
    .B1(_17550_),
    .B2(_17551_),
    .ZN(_17552_));
 AOI21_X2 _44328_ (.A(_17300_),
    .B1(_17549_),
    .B2(_17552_),
    .ZN(_17553_));
 BUF_X16 _44329_ (.A(_15331_),
    .Z(_17554_));
 NOR2_X1 _44330_ (.A1(_16274_),
    .A2(_15533_),
    .ZN(_17555_));
 AND2_X1 _44331_ (.A1(_15784_),
    .A2(\icache.data_mems_2__data_mem.data_o [44]),
    .ZN(_17556_));
 OAI21_X2 _44332_ (.A(_17554_),
    .B1(_17555_),
    .B2(_17556_),
    .ZN(_17557_));
 NOR2_X2 _44333_ (.A1(_16269_),
    .A2(_15518_),
    .ZN(_17558_));
 AND2_X1 _44334_ (.A1(_16061_),
    .A2(\icache.data_mems_0__data_mem.data_o [44]),
    .ZN(_17559_));
 OAI21_X2 _44335_ (.A(_15650_),
    .B1(_17558_),
    .B2(_17559_),
    .ZN(_17560_));
 AOI21_X2 _44336_ (.A(_16714_),
    .B1(_17557_),
    .B2(_17560_),
    .ZN(_17561_));
 NOR2_X4 _44337_ (.A1(_17553_),
    .A2(_17561_),
    .ZN(_17562_));
 OAI21_X1 _44338_ (.A(_17546_),
    .B1(_17562_),
    .B2(_17404_),
    .ZN(_05324_));
 NAND2_X1 _44339_ (.A1(_17526_),
    .A2(\icache.lce.lce_cmd_inst.data_r [394]),
    .ZN(_17563_));
 NOR2_X2 _44340_ (.A1(_16854_),
    .A2(_15318_),
    .ZN(_17564_));
 AND2_X1 _44341_ (.A1(_15541_),
    .A2(\icache.data_mems_3__data_mem.data_o [10]),
    .ZN(_17565_));
 OAI21_X2 _44342_ (.A(_16099_),
    .B1(_17564_),
    .B2(_17565_),
    .ZN(_17566_));
 BUF_X16 _44343_ (.A(_15734_),
    .Z(_17567_));
 NAND2_X1 _44344_ (.A1(_16391_),
    .A2(_16860_),
    .ZN(_17568_));
 NAND2_X1 _44345_ (.A1(_16858_),
    .A2(_16394_),
    .ZN(_17569_));
 NAND3_X2 _44346_ (.A1(_17568_),
    .A2(_17569_),
    .A3(_15446_),
    .ZN(_17570_));
 NAND3_X2 _44347_ (.A1(_17566_),
    .A2(_17567_),
    .A3(_17570_),
    .ZN(_17571_));
 NOR2_X1 _44348_ (.A1(_16872_),
    .A2(_15443_),
    .ZN(_17572_));
 AND2_X1 _44349_ (.A1(_15438_),
    .A2(\icache.data_mems_7__data_mem.data_o [10]),
    .ZN(_17573_));
 OAI21_X2 _44350_ (.A(_15450_),
    .B1(_17572_),
    .B2(_17573_),
    .ZN(_17574_));
 OR2_X1 _44351_ (.A1(_15776_),
    .A2(\icache.data_mems_4__data_mem.data_o [10]),
    .ZN(_17575_));
 NAND2_X1 _44352_ (.A1(_16866_),
    .A2(_16169_),
    .ZN(_17576_));
 NAND3_X2 _44353_ (.A1(_17575_),
    .A2(_17576_),
    .A3(_15994_),
    .ZN(_17577_));
 NAND3_X2 _44354_ (.A1(_17574_),
    .A2(_16823_),
    .A3(_17577_),
    .ZN(_17578_));
 NAND2_X4 _44355_ (.A1(_17571_),
    .A2(_17578_),
    .ZN(_17579_));
 BUF_X4 _44356_ (.A(_16785_),
    .Z(_17580_));
 OAI21_X1 _44357_ (.A(_17563_),
    .B1(_17579_),
    .B2(_17580_),
    .ZN(_05215_));
 NAND2_X1 _44358_ (.A1(_17526_),
    .A2(\icache.lce.lce_cmd_inst.data_r [395]),
    .ZN(_17581_));
 BUF_X8 _44359_ (.A(_15597_),
    .Z(_17582_));
 OR2_X2 _44360_ (.A1(_16015_),
    .A2(\icache.data_mems_4__data_mem.data_o [11]),
    .ZN(_17583_));
 NAND2_X2 _44361_ (.A1(_16878_),
    .A2(_16018_),
    .ZN(_17584_));
 AOI21_X2 _44362_ (.A(_15379_),
    .B1(_17583_),
    .B2(_17584_),
    .ZN(_17585_));
 INV_X1 _44363_ (.A(\icache.data_mems_6__data_mem.data_o [11]),
    .ZN(_17586_));
 NAND2_X2 _44364_ (.A1(_15747_),
    .A2(_17586_),
    .ZN(_17587_));
 NAND2_X2 _44365_ (.A1(_16883_),
    .A2(_15752_),
    .ZN(_17588_));
 AOI21_X2 _44366_ (.A(_16005_),
    .B1(_17587_),
    .B2(_17588_),
    .ZN(_17589_));
 OAI21_X2 _44367_ (.A(_17582_),
    .B1(_17585_),
    .B2(_17589_),
    .ZN(_17590_));
 NAND2_X1 _44368_ (.A1(_15671_),
    .A2(\icache.data_mems_0__data_mem.data_o [11]),
    .ZN(_17591_));
 NAND2_X1 _44369_ (.A1(_15967_),
    .A2(\icache.data_mems_1__data_mem.data_o [11]),
    .ZN(_17592_));
 AND3_X1 _44370_ (.A1(_17591_),
    .A2(_16418_),
    .A3(_17592_),
    .ZN(_17593_));
 NAND2_X1 _44371_ (.A1(_15537_),
    .A2(_16891_),
    .ZN(_17594_));
 NAND2_X1 _44372_ (.A1(_16889_),
    .A2(_15810_),
    .ZN(_17595_));
 AOI21_X2 _44373_ (.A(_17016_),
    .B1(_17594_),
    .B2(_17595_),
    .ZN(_17596_));
 OAI21_X2 _44374_ (.A(_17500_),
    .B1(_17593_),
    .B2(_17596_),
    .ZN(_17597_));
 NAND2_X4 _44375_ (.A1(_17590_),
    .A2(_17597_),
    .ZN(_17598_));
 OAI21_X1 _44376_ (.A(_17581_),
    .B1(_17598_),
    .B2(_17580_),
    .ZN(_05216_));
 NAND2_X1 _44377_ (.A1(_17526_),
    .A2(\icache.lce.lce_cmd_inst.data_r [396]),
    .ZN(_17599_));
 NOR2_X1 _44378_ (.A1(_16901_),
    .A2(_15478_),
    .ZN(_17600_));
 AND2_X1 _44379_ (.A1(_15876_),
    .A2(\icache.data_mems_7__data_mem.data_o [12]),
    .ZN(_17601_));
 OR3_X1 _44380_ (.A1(_17600_),
    .A2(_17601_),
    .A3(_16226_),
    .ZN(_17602_));
 NAND2_X1 _44381_ (.A1(_15756_),
    .A2(\icache.data_mems_4__data_mem.data_o [12]),
    .ZN(_17603_));
 NAND2_X1 _44382_ (.A1(_15443_),
    .A2(\icache.data_mems_5__data_mem.data_o [12]),
    .ZN(_17604_));
 NAND3_X1 _44383_ (.A1(_17603_),
    .A2(_15932_),
    .A3(_17604_),
    .ZN(_17605_));
 NAND3_X1 _44384_ (.A1(_17602_),
    .A2(_16360_),
    .A3(_17605_),
    .ZN(_17606_));
 NAND2_X1 _44385_ (.A1(_16155_),
    .A2(_16909_),
    .ZN(_17607_));
 NAND2_X1 _44386_ (.A1(_16907_),
    .A2(_15338_),
    .ZN(_17608_));
 AND3_X1 _44387_ (.A1(_17607_),
    .A2(_17608_),
    .A3(_16634_),
    .ZN(_17609_));
 NAND2_X1 _44388_ (.A1(_15671_),
    .A2(\icache.data_mems_2__data_mem.data_o [12]),
    .ZN(_17610_));
 NAND2_X1 _44389_ (.A1(_15725_),
    .A2(\icache.data_mems_3__data_mem.data_o [12]),
    .ZN(_17611_));
 AOI21_X1 _44390_ (.A(_15727_),
    .B1(_17610_),
    .B2(_17611_),
    .ZN(_17612_));
 OAI21_X1 _44391_ (.A(_16640_),
    .B1(_17609_),
    .B2(_17612_),
    .ZN(_17613_));
 AND2_X4 _44392_ (.A1(_17606_),
    .A2(_17613_),
    .ZN(_17614_));
 OAI21_X1 _44393_ (.A(_17599_),
    .B1(_17614_),
    .B2(_17580_),
    .ZN(_05217_));
 NAND2_X1 _44394_ (.A1(_17526_),
    .A2(\icache.lce.lce_cmd_inst.data_r [397]),
    .ZN(_17615_));
 OR2_X1 _44395_ (.A1(_15714_),
    .A2(\icache.data_mems_6__data_mem.data_o [13]),
    .ZN(_17616_));
 NAND2_X1 _44396_ (.A1(_16924_),
    .A2(_16408_),
    .ZN(_17617_));
 NAND2_X1 _44397_ (.A1(_17616_),
    .A2(_17617_),
    .ZN(_17618_));
 NAND2_X1 _44398_ (.A1(_17618_),
    .A2(_16341_),
    .ZN(_17619_));
 NAND2_X1 _44399_ (.A1(_15398_),
    .A2(_16930_),
    .ZN(_17620_));
 NAND2_X1 _44400_ (.A1(_16928_),
    .A2(_15402_),
    .ZN(_17621_));
 NAND2_X1 _44401_ (.A1(_17620_),
    .A2(_17621_),
    .ZN(_17622_));
 NAND2_X1 _44402_ (.A1(_17622_),
    .A2(_16347_),
    .ZN(_17623_));
 NAND2_X1 _44403_ (.A1(_17619_),
    .A2(_17623_),
    .ZN(_17624_));
 NAND2_X1 _44404_ (.A1(_17624_),
    .A2(_16266_),
    .ZN(_17625_));
 NAND2_X1 _44405_ (.A1(_15836_),
    .A2(_16920_),
    .ZN(_17626_));
 NAND2_X1 _44406_ (.A1(_16918_),
    .A2(_15541_),
    .ZN(_17627_));
 NAND2_X2 _44407_ (.A1(_17626_),
    .A2(_17627_),
    .ZN(_17628_));
 NAND2_X1 _44408_ (.A1(_17628_),
    .A2(_15587_),
    .ZN(_17629_));
 NAND2_X1 _44409_ (.A1(_16343_),
    .A2(\icache.data_mems_2__data_mem.data_o [13]),
    .ZN(_17630_));
 NAND2_X1 _44410_ (.A1(_16083_),
    .A2(\icache.data_mems_3__data_mem.data_o [13]),
    .ZN(_17631_));
 NAND3_X1 _44411_ (.A1(_17630_),
    .A2(_15395_),
    .A3(_17631_),
    .ZN(_17632_));
 NAND2_X1 _44412_ (.A1(_17629_),
    .A2(_17632_),
    .ZN(_17633_));
 BUF_X16 _44413_ (.A(_16314_),
    .Z(_17634_));
 NAND2_X1 _44414_ (.A1(_17633_),
    .A2(_17634_),
    .ZN(_17635_));
 NAND2_X4 _44415_ (.A1(_17625_),
    .A2(_17635_),
    .ZN(_17636_));
 OAI21_X1 _44416_ (.A(_17615_),
    .B1(_17636_),
    .B2(_17580_),
    .ZN(_05218_));
 NAND2_X1 _44417_ (.A1(_17526_),
    .A2(\icache.lce.lce_cmd_inst.data_r [398]),
    .ZN(_17637_));
 NOR2_X1 _44418_ (.A1(_16950_),
    .A2(_15541_),
    .ZN(_17638_));
 AND2_X1 _44419_ (.A1(_15334_),
    .A2(\icache.data_mems_5__data_mem.data_o [14]),
    .ZN(_17639_));
 NOR2_X1 _44420_ (.A1(_17638_),
    .A2(_17639_),
    .ZN(_17640_));
 NOR2_X1 _44421_ (.A1(_17640_),
    .A2(_15545_),
    .ZN(_17641_));
 NAND2_X1 _44422_ (.A1(_15719_),
    .A2(\icache.data_mems_6__data_mem.data_o [14]),
    .ZN(_17642_));
 NAND2_X1 _44423_ (.A1(_15475_),
    .A2(\icache.data_mems_7__data_mem.data_o [14]),
    .ZN(_17643_));
 AOI21_X1 _44424_ (.A(_16056_),
    .B1(_17642_),
    .B2(_17643_),
    .ZN(_17644_));
 OAI21_X1 _44425_ (.A(_16631_),
    .B1(_17641_),
    .B2(_17644_),
    .ZN(_17645_));
 NAND2_X1 _44426_ (.A1(_16391_),
    .A2(\icache.data_mems_2__data_mem.data_o [14]),
    .ZN(_17646_));
 OAI211_X2 _44427_ (.A(_17646_),
    .B(_15425_),
    .C1(_15721_),
    .C2(_16940_),
    .ZN(_17647_));
 NAND2_X1 _44428_ (.A1(_16222_),
    .A2(\icache.data_mems_0__data_mem.data_o [14]),
    .ZN(_17648_));
 NAND2_X1 _44429_ (.A1(_15725_),
    .A2(\icache.data_mems_1__data_mem.data_o [14]),
    .ZN(_17649_));
 NAND3_X2 _44430_ (.A1(_17648_),
    .A2(_15406_),
    .A3(_17649_),
    .ZN(_17650_));
 NAND3_X1 _44431_ (.A1(_17647_),
    .A2(_16372_),
    .A3(_17650_),
    .ZN(_17651_));
 AND2_X4 _44432_ (.A1(_17645_),
    .A2(_17651_),
    .ZN(_17652_));
 OAI21_X1 _44433_ (.A(_17637_),
    .B1(_17652_),
    .B2(_17580_),
    .ZN(_05219_));
 NAND2_X1 _44434_ (.A1(_17526_),
    .A2(\icache.lce.lce_cmd_inst.data_r [399]),
    .ZN(_17653_));
 OR2_X1 _44435_ (.A1(_15967_),
    .A2(\icache.data_mems_0__data_mem.data_o [15]),
    .ZN(_17654_));
 NAND2_X1 _44436_ (.A1(_16961_),
    .A2(_15728_),
    .ZN(_17655_));
 AOI21_X2 _44437_ (.A(_15379_),
    .B1(_17654_),
    .B2(_17655_),
    .ZN(_17656_));
 OR2_X1 _44438_ (.A1(_15573_),
    .A2(\icache.data_mems_2__data_mem.data_o [15]),
    .ZN(_17657_));
 NAND2_X2 _44439_ (.A1(_16957_),
    .A2(_15752_),
    .ZN(_17658_));
 AOI21_X2 _44440_ (.A(_16005_),
    .B1(_17657_),
    .B2(_17658_),
    .ZN(_17659_));
 OAI21_X2 _44441_ (.A(_15735_),
    .B1(_17656_),
    .B2(_17659_),
    .ZN(_17660_));
 OR2_X1 _44442_ (.A1(_15967_),
    .A2(\icache.data_mems_4__data_mem.data_o [15]),
    .ZN(_17661_));
 NAND2_X1 _44443_ (.A1(_16966_),
    .A2(_15728_),
    .ZN(_17662_));
 NAND3_X2 _44444_ (.A1(_17661_),
    .A2(_17662_),
    .A3(_15761_),
    .ZN(_17663_));
 NAND2_X2 _44445_ (.A1(_15747_),
    .A2(_16972_),
    .ZN(_17664_));
 NAND2_X2 _44446_ (.A1(_16970_),
    .A2(_15752_),
    .ZN(_17665_));
 NAND3_X2 _44447_ (.A1(_17664_),
    .A2(_17665_),
    .A3(_15708_),
    .ZN(_17666_));
 NAND3_X2 _44448_ (.A1(_17663_),
    .A2(_17666_),
    .A3(_15656_),
    .ZN(_17667_));
 NAND2_X4 _44449_ (.A1(_17660_),
    .A2(_17667_),
    .ZN(_17668_));
 OAI21_X1 _44450_ (.A(_17653_),
    .B1(_17668_),
    .B2(_17580_),
    .ZN(_05220_));
 NAND2_X1 _44451_ (.A1(_17526_),
    .A2(\icache.lce.lce_cmd_inst.data_r [400]),
    .ZN(_17669_));
 NOR2_X1 _44452_ (.A1(_16992_),
    .A2(_15505_),
    .ZN(_17670_));
 AND2_X1 _44453_ (.A1(_15471_),
    .A2(\icache.data_mems_3__data_mem.data_o [16]),
    .ZN(_17671_));
 OR3_X1 _44454_ (.A1(_17670_),
    .A2(_17671_),
    .A3(_16226_),
    .ZN(_17672_));
 OR2_X1 _44455_ (.A1(_15317_),
    .A2(\icache.data_mems_0__data_mem.data_o [16]),
    .ZN(_17673_));
 NAND2_X1 _44456_ (.A1(_16987_),
    .A2(_15402_),
    .ZN(_17674_));
 NAND2_X1 _44457_ (.A1(_17673_),
    .A2(_17674_),
    .ZN(_17675_));
 NAND2_X1 _44458_ (.A1(_17675_),
    .A2(_16347_),
    .ZN(_17676_));
 NAND2_X1 _44459_ (.A1(_17672_),
    .A2(_17676_),
    .ZN(_17677_));
 NAND2_X1 _44460_ (.A1(_17677_),
    .A2(_15580_),
    .ZN(_17678_));
 NAND2_X1 _44461_ (.A1(_16155_),
    .A2(\icache.data_mems_4__data_mem.data_o [16]),
    .ZN(_17679_));
 NAND2_X1 _44462_ (.A1(_15606_),
    .A2(\icache.data_mems_5__data_mem.data_o [16]),
    .ZN(_17680_));
 AND3_X1 _44463_ (.A1(_17679_),
    .A2(_16418_),
    .A3(_17680_),
    .ZN(_17681_));
 NAND2_X1 _44464_ (.A1(_15491_),
    .A2(_16983_),
    .ZN(_17682_));
 NAND2_X2 _44465_ (.A1(_16981_),
    .A2(_16067_),
    .ZN(_17683_));
 AOI21_X2 _44466_ (.A(_17016_),
    .B1(_17682_),
    .B2(_17683_),
    .ZN(_17684_));
 OAI21_X2 _44467_ (.A(_16013_),
    .B1(_17681_),
    .B2(_17684_),
    .ZN(_17685_));
 NAND2_X4 _44468_ (.A1(_17678_),
    .A2(_17685_),
    .ZN(_17686_));
 OAI21_X1 _44469_ (.A(_17669_),
    .B1(_17686_),
    .B2(_17580_),
    .ZN(_05223_));
 NAND2_X1 _44470_ (.A1(_17526_),
    .A2(\icache.lce.lce_cmd_inst.data_r [401]),
    .ZN(_17687_));
 NOR2_X4 _44471_ (.A1(_17000_),
    .A2(_15810_),
    .ZN(_17688_));
 AND2_X1 _44472_ (.A1(_15550_),
    .A2(\icache.data_mems_3__data_mem.data_o [17]),
    .ZN(_17689_));
 OR3_X1 _44473_ (.A1(_17688_),
    .A2(_17689_),
    .A3(_16226_),
    .ZN(_17690_));
 NAND2_X1 _44474_ (.A1(_15569_),
    .A2(_17006_),
    .ZN(_17691_));
 NAND2_X1 _44475_ (.A1(_17004_),
    .A2(_15564_),
    .ZN(_17692_));
 NAND2_X1 _44476_ (.A1(_17691_),
    .A2(_17692_),
    .ZN(_17693_));
 NAND2_X1 _44477_ (.A1(_17693_),
    .A2(_16347_),
    .ZN(_17694_));
 NAND2_X2 _44478_ (.A1(_17690_),
    .A2(_17694_),
    .ZN(_17695_));
 NAND2_X2 _44479_ (.A1(_17695_),
    .A2(_15580_),
    .ZN(_17696_));
 NOR2_X2 _44480_ (.A1(_17018_),
    .A2(_15436_),
    .ZN(_17697_));
 AND2_X1 _44481_ (.A1(_15916_),
    .A2(\icache.data_mems_7__data_mem.data_o [17]),
    .ZN(_17698_));
 NOR3_X2 _44482_ (.A1(_17697_),
    .A2(_17698_),
    .A3(_15932_),
    .ZN(_17699_));
 OR2_X1 _44483_ (.A1(_16272_),
    .A2(\icache.data_mems_4__data_mem.data_o [17]),
    .ZN(_17700_));
 NAND2_X1 _44484_ (.A1(_17012_),
    .A2(_16805_),
    .ZN(_17701_));
 AOI21_X2 _44485_ (.A(_16544_),
    .B1(_17700_),
    .B2(_17701_),
    .ZN(_17702_));
 OAI21_X2 _44486_ (.A(_16013_),
    .B1(_17699_),
    .B2(_17702_),
    .ZN(_17703_));
 NAND2_X4 _44487_ (.A1(_17696_),
    .A2(_17703_),
    .ZN(_17704_));
 OAI21_X1 _44488_ (.A(_17687_),
    .B1(_17704_),
    .B2(_17580_),
    .ZN(_05224_));
 BUF_X4 _44489_ (.A(_16724_),
    .Z(_17705_));
 NAND2_X1 _44490_ (.A1(_17705_),
    .A2(\icache.lce.lce_cmd_inst.data_r [402]),
    .ZN(_17706_));
 OR2_X1 _44491_ (.A1(_16083_),
    .A2(\icache.data_mems_2__data_mem.data_o [18]),
    .ZN(_17707_));
 NAND2_X2 _44492_ (.A1(_17033_),
    .A2(_15986_),
    .ZN(_17708_));
 AOI21_X2 _44493_ (.A(_15343_),
    .B1(_17707_),
    .B2(_17708_),
    .ZN(_17709_));
 BUF_X16 _44494_ (.A(_15394_),
    .Z(_17710_));
 NAND2_X1 _44495_ (.A1(_15747_),
    .A2(_17039_),
    .ZN(_17711_));
 NAND2_X2 _44496_ (.A1(_17037_),
    .A2(_15752_),
    .ZN(_17712_));
 AOI21_X2 _44497_ (.A(_17710_),
    .B1(_17711_),
    .B2(_17712_),
    .ZN(_17713_));
 OAI21_X2 _44498_ (.A(_15735_),
    .B1(_17709_),
    .B2(_17713_),
    .ZN(_17714_));
 NAND2_X1 _44499_ (.A1(_15671_),
    .A2(\icache.data_mems_6__data_mem.data_o [18]),
    .ZN(_17715_));
 NAND2_X1 _44500_ (.A1(_15725_),
    .A2(\icache.data_mems_7__data_mem.data_o [18]),
    .ZN(_17716_));
 AND3_X1 _44501_ (.A1(_17715_),
    .A2(_16541_),
    .A3(_17716_),
    .ZN(_17717_));
 NAND2_X1 _44502_ (.A1(_15537_),
    .A2(_17029_),
    .ZN(_17718_));
 NAND2_X1 _44503_ (.A1(_17027_),
    .A2(_15810_),
    .ZN(_17719_));
 AOI21_X2 _44504_ (.A(_16544_),
    .B1(_17718_),
    .B2(_17719_),
    .ZN(_17720_));
 OAI21_X2 _44505_ (.A(_16013_),
    .B1(_17717_),
    .B2(_17720_),
    .ZN(_17721_));
 NAND2_X4 _44506_ (.A1(_17714_),
    .A2(_17721_),
    .ZN(_17722_));
 OAI21_X1 _44507_ (.A(_17706_),
    .B1(_17722_),
    .B2(_17580_),
    .ZN(_05225_));
 NAND2_X1 _44508_ (.A1(_17705_),
    .A2(\icache.lce.lce_cmd_inst.data_r [403]),
    .ZN(_17723_));
 NOR2_X1 _44509_ (.A1(_17049_),
    .A2(_15460_),
    .ZN(_17724_));
 AND2_X1 _44510_ (.A1(_15308_),
    .A2(\icache.data_mems_3__data_mem.data_o [19]),
    .ZN(_17725_));
 OR3_X1 _44511_ (.A1(_17724_),
    .A2(_17725_),
    .A3(_16226_),
    .ZN(_17726_));
 NAND2_X1 _44512_ (.A1(_16391_),
    .A2(\icache.data_mems_0__data_mem.data_o [19]),
    .ZN(_17727_));
 NAND2_X1 _44513_ (.A1(_16394_),
    .A2(\icache.data_mems_1__data_mem.data_o [19]),
    .ZN(_17728_));
 NAND3_X1 _44514_ (.A1(_17727_),
    .A2(_15610_),
    .A3(_17728_),
    .ZN(_17729_));
 NAND2_X2 _44515_ (.A1(_17726_),
    .A2(_17729_),
    .ZN(_17730_));
 BUF_X16 _44516_ (.A(_15579_),
    .Z(_17731_));
 NAND2_X1 _44517_ (.A1(_17730_),
    .A2(_17731_),
    .ZN(_17732_));
 NAND2_X1 _44518_ (.A1(_15674_),
    .A2(_17060_),
    .ZN(_17733_));
 NAND2_X1 _44519_ (.A1(_17058_),
    .A2(_15986_),
    .ZN(_17734_));
 AOI21_X2 _44520_ (.A(_16014_),
    .B1(_17733_),
    .B2(_17734_),
    .ZN(_17735_));
 NAND2_X1 _44521_ (.A1(_16580_),
    .A2(_17055_),
    .ZN(_17736_));
 NAND2_X1 _44522_ (.A1(_17053_),
    .A2(_16805_),
    .ZN(_17737_));
 AOI21_X2 _44523_ (.A(_17016_),
    .B1(_17736_),
    .B2(_17737_),
    .ZN(_17738_));
 OAI21_X2 _44524_ (.A(_16013_),
    .B1(_17735_),
    .B2(_17738_),
    .ZN(_17739_));
 NAND2_X4 _44525_ (.A1(_17732_),
    .A2(_17739_),
    .ZN(_17740_));
 OAI21_X1 _44526_ (.A(_17723_),
    .B1(_17740_),
    .B2(_17580_),
    .ZN(_05226_));
 NAND2_X1 _44527_ (.A1(_17705_),
    .A2(\icache.lce.lce_cmd_inst.data_r [404]),
    .ZN(_17741_));
 NOR2_X1 _44528_ (.A1(_17071_),
    .A2(_15460_),
    .ZN(_17742_));
 AND2_X1 _44529_ (.A1(_15488_),
    .A2(\icache.data_mems_1__data_mem.data_o [20]),
    .ZN(_17743_));
 NOR2_X1 _44530_ (.A1(_17742_),
    .A2(_17743_),
    .ZN(_17744_));
 NOR2_X1 _44531_ (.A1(_17744_),
    .A2(_15545_),
    .ZN(_17745_));
 NAND2_X1 _44532_ (.A1(_15836_),
    .A2(\icache.data_mems_2__data_mem.data_o [20]),
    .ZN(_17746_));
 NAND2_X1 _44533_ (.A1(_15511_),
    .A2(\icache.data_mems_3__data_mem.data_o [20]),
    .ZN(_17747_));
 AOI21_X1 _44534_ (.A(_16056_),
    .B1(_17746_),
    .B2(_17747_),
    .ZN(_17748_));
 OAI21_X1 _44535_ (.A(_16438_),
    .B1(_17745_),
    .B2(_17748_),
    .ZN(_17749_));
 NOR2_X1 _44536_ (.A1(_17075_),
    .A2(_15460_),
    .ZN(_17750_));
 AND2_X1 _44537_ (.A1(_15784_),
    .A2(\icache.data_mems_5__data_mem.data_o [20]),
    .ZN(_17751_));
 OR3_X1 _44538_ (.A1(_17750_),
    .A2(_17751_),
    .A3(_15311_),
    .ZN(_17752_));
 NAND2_X1 _44539_ (.A1(_15335_),
    .A2(\icache.data_mems_7__data_mem.data_o [20]),
    .ZN(_17753_));
 OAI211_X2 _44540_ (.A(_17753_),
    .B(_17511_),
    .C1(_15324_),
    .C2(_17081_),
    .ZN(_17754_));
 NAND3_X1 _44541_ (.A1(_17752_),
    .A2(_15409_),
    .A3(_17754_),
    .ZN(_17755_));
 AND2_X4 _44542_ (.A1(_17749_),
    .A2(_17755_),
    .ZN(_17756_));
 BUF_X4 _44543_ (.A(_16785_),
    .Z(_17757_));
 OAI21_X1 _44544_ (.A(_17741_),
    .B1(_17756_),
    .B2(_17757_),
    .ZN(_05227_));
 NAND2_X1 _44545_ (.A1(_17705_),
    .A2(\icache.lce.lce_cmd_inst.data_r [405]),
    .ZN(_17758_));
 NOR2_X1 _44546_ (.A1(_15523_),
    .A2(\icache.data_mems_1__data_mem.data_o [21]),
    .ZN(_17759_));
 AOI211_X1 _44547_ (.A(_16229_),
    .B(_17759_),
    .C1(_15679_),
    .C2(_17103_),
    .ZN(_17760_));
 NAND2_X1 _44548_ (.A1(_15612_),
    .A2(\icache.data_mems_2__data_mem.data_o [21]),
    .ZN(_17761_));
 NAND2_X1 _44549_ (.A1(_15346_),
    .A2(\icache.data_mems_3__data_mem.data_o [21]),
    .ZN(_17762_));
 AOI21_X1 _44550_ (.A(_16634_),
    .B1(_17761_),
    .B2(_17762_),
    .ZN(_17763_));
 OAI21_X1 _44551_ (.A(_16438_),
    .B1(_17760_),
    .B2(_17763_),
    .ZN(_17764_));
 NOR2_X1 _44552_ (.A1(_17093_),
    .A2(_15317_),
    .ZN(_17765_));
 AND2_X1 _44553_ (.A1(_15322_),
    .A2(\icache.data_mems_7__data_mem.data_o [21]),
    .ZN(_17766_));
 OR3_X2 _44554_ (.A1(_17765_),
    .A2(_17766_),
    .A3(_15483_),
    .ZN(_17767_));
 NAND2_X1 _44555_ (.A1(_15372_),
    .A2(\icache.data_mems_4__data_mem.data_o [21]),
    .ZN(_17768_));
 OAI211_X2 _44556_ (.A(_17768_),
    .B(_16307_),
    .C1(_15756_),
    .C2(_17088_),
    .ZN(_17769_));
 NAND3_X1 _44557_ (.A1(_17767_),
    .A2(_17415_),
    .A3(_17769_),
    .ZN(_17770_));
 AND2_X4 _44558_ (.A1(_17764_),
    .A2(_17770_),
    .ZN(_17771_));
 OAI21_X1 _44559_ (.A(_17758_),
    .B1(_17771_),
    .B2(_17757_),
    .ZN(_05228_));
 NAND2_X1 _44560_ (.A1(_17705_),
    .A2(\icache.lce.lce_cmd_inst.data_r [406]),
    .ZN(_17772_));
 OR2_X1 _44561_ (.A1(_15533_),
    .A2(\icache.data_mems_4__data_mem.data_o [22]),
    .ZN(_17773_));
 NAND2_X1 _44562_ (.A1(_17120_),
    .A2(_15573_),
    .ZN(_17774_));
 NAND2_X1 _44563_ (.A1(_17773_),
    .A2(_17774_),
    .ZN(_17775_));
 NAND2_X1 _44564_ (.A1(_17775_),
    .A2(_16256_),
    .ZN(_17776_));
 OR2_X1 _44565_ (.A1(_15486_),
    .A2(\icache.data_mems_6__data_mem.data_o [22]),
    .ZN(_17777_));
 NAND2_X1 _44566_ (.A1(_17116_),
    .A2(_15564_),
    .ZN(_17778_));
 NAND2_X1 _44567_ (.A1(_17777_),
    .A2(_17778_),
    .ZN(_17779_));
 NAND2_X1 _44568_ (.A1(_17779_),
    .A2(_16262_),
    .ZN(_17780_));
 NAND2_X2 _44569_ (.A1(_17776_),
    .A2(_17780_),
    .ZN(_17781_));
 NAND2_X1 _44570_ (.A1(_17781_),
    .A2(_16266_),
    .ZN(_17782_));
 NAND2_X1 _44571_ (.A1(_16391_),
    .A2(\icache.data_mems_0__data_mem.data_o [22]),
    .ZN(_17783_));
 NAND2_X1 _44572_ (.A1(_16394_),
    .A2(\icache.data_mems_1__data_mem.data_o [22]),
    .ZN(_17784_));
 NAND3_X1 _44573_ (.A1(_17783_),
    .A2(_15610_),
    .A3(_17784_),
    .ZN(_17785_));
 NAND2_X1 _44574_ (.A1(_16222_),
    .A2(\icache.data_mems_2__data_mem.data_o [22]),
    .ZN(_17786_));
 NAND2_X1 _44575_ (.A1(_15725_),
    .A2(\icache.data_mems_3__data_mem.data_o [22]),
    .ZN(_17787_));
 NAND3_X1 _44576_ (.A1(_17786_),
    .A2(_15395_),
    .A3(_17787_),
    .ZN(_17788_));
 NAND2_X2 _44577_ (.A1(_17785_),
    .A2(_17788_),
    .ZN(_17789_));
 NAND2_X1 _44578_ (.A1(_17789_),
    .A2(_17634_),
    .ZN(_17790_));
 NAND2_X4 _44579_ (.A1(_17782_),
    .A2(_17790_),
    .ZN(_17791_));
 OAI21_X1 _44580_ (.A(_17772_),
    .B1(_17791_),
    .B2(_17757_),
    .ZN(_05229_));
 NAND2_X1 _44581_ (.A1(_17705_),
    .A2(\icache.lce.lce_cmd_inst.data_r [407]),
    .ZN(_17792_));
 NAND2_X1 _44582_ (.A1(_15537_),
    .A2(_17132_),
    .ZN(_17793_));
 NAND2_X2 _44583_ (.A1(_17130_),
    .A2(_15810_),
    .ZN(_17794_));
 AND3_X1 _44584_ (.A1(_17793_),
    .A2(_17794_),
    .A3(_15445_),
    .ZN(_17795_));
 NAND2_X2 _44585_ (.A1(_15671_),
    .A2(\icache.data_mems_6__data_mem.data_o [23]),
    .ZN(_17796_));
 NAND2_X2 _44586_ (.A1(_15725_),
    .A2(\icache.data_mems_7__data_mem.data_o [23]),
    .ZN(_17797_));
 AOI21_X4 _44587_ (.A(_15727_),
    .B1(_17796_),
    .B2(_17797_),
    .ZN(_17798_));
 NOR2_X2 _44588_ (.A1(_17795_),
    .A2(_17798_),
    .ZN(_17799_));
 NOR2_X1 _44589_ (.A1(_17799_),
    .A2(_15354_),
    .ZN(_17800_));
 NOR2_X2 _44590_ (.A1(_17139_),
    .A2(_16867_),
    .ZN(_17801_));
 AND2_X1 _44591_ (.A1(_15454_),
    .A2(\icache.data_mems_1__data_mem.data_o [23]),
    .ZN(_17802_));
 OAI21_X2 _44592_ (.A(_16865_),
    .B1(_17801_),
    .B2(_17802_),
    .ZN(_17803_));
 NAND2_X1 _44593_ (.A1(_15747_),
    .A2(_17144_),
    .ZN(_17804_));
 NAND2_X2 _44594_ (.A1(_17142_),
    .A2(_15461_),
    .ZN(_17805_));
 NAND3_X2 _44595_ (.A1(_17804_),
    .A2(_17805_),
    .A3(_16583_),
    .ZN(_17806_));
 AOI21_X2 _44596_ (.A(_16714_),
    .B1(_17803_),
    .B2(_17806_),
    .ZN(_17807_));
 NOR2_X4 _44597_ (.A1(_17800_),
    .A2(_17807_),
    .ZN(_17808_));
 OAI21_X1 _44598_ (.A(_17792_),
    .B1(_17808_),
    .B2(_17757_),
    .ZN(_05230_));
 NAND2_X1 _44599_ (.A1(_17705_),
    .A2(\icache.lce.lce_cmd_inst.data_r [408]),
    .ZN(_17809_));
 NOR2_X2 _44600_ (.A1(_17163_),
    .A2(_16001_),
    .ZN(_17810_));
 AND2_X1 _44601_ (.A1(_16253_),
    .A2(\icache.data_mems_7__data_mem.data_o [24]),
    .ZN(_17811_));
 OAI21_X2 _44602_ (.A(_15708_),
    .B1(_17810_),
    .B2(_17811_),
    .ZN(_17812_));
 NOR2_X1 _44603_ (.A1(_17167_),
    .A2(_15436_),
    .ZN(_17813_));
 AND2_X1 _44604_ (.A1(_16272_),
    .A2(\icache.data_mems_5__data_mem.data_o [24]),
    .ZN(_17814_));
 OAI21_X2 _44605_ (.A(_15712_),
    .B1(_17813_),
    .B2(_17814_),
    .ZN(_17815_));
 AOI21_X2 _44606_ (.A(_17300_),
    .B1(_17812_),
    .B2(_17815_),
    .ZN(_17816_));
 BUF_X16 _44607_ (.A(_15367_),
    .Z(_17817_));
 NAND2_X1 _44608_ (.A1(_15674_),
    .A2(_17158_),
    .ZN(_17818_));
 NAND2_X2 _44609_ (.A1(_17156_),
    .A2(_15986_),
    .ZN(_17819_));
 NAND3_X2 _44610_ (.A1(_17818_),
    .A2(_17819_),
    .A3(_15988_),
    .ZN(_17820_));
 NAND2_X2 _44611_ (.A1(_15747_),
    .A2(_17153_),
    .ZN(_17821_));
 NAND2_X1 _44612_ (.A1(_17151_),
    .A2(_15461_),
    .ZN(_17822_));
 NAND3_X2 _44613_ (.A1(_17821_),
    .A2(_17822_),
    .A3(_16217_),
    .ZN(_17823_));
 AOI21_X2 _44614_ (.A(_17817_),
    .B1(_17820_),
    .B2(_17823_),
    .ZN(_17824_));
 NOR2_X4 _44615_ (.A1(_17816_),
    .A2(_17824_),
    .ZN(_17825_));
 OAI21_X1 _44616_ (.A(_17809_),
    .B1(_17825_),
    .B2(_17757_),
    .ZN(_05231_));
 NAND2_X1 _44617_ (.A1(_17705_),
    .A2(\icache.lce.lce_cmd_inst.data_r [409]),
    .ZN(_17826_));
 BUF_X16 _44618_ (.A(_15734_),
    .Z(_17827_));
 NOR2_X1 _44619_ (.A1(_17191_),
    .A2(_16867_),
    .ZN(_17828_));
 AND2_X1 _44620_ (.A1(_15606_),
    .A2(\icache.data_mems_3__data_mem.data_o [25]),
    .ZN(_17829_));
 NOR3_X2 _44621_ (.A1(_17828_),
    .A2(_17829_),
    .A3(_15932_),
    .ZN(_17830_));
 OR2_X1 _44622_ (.A1(_16272_),
    .A2(\icache.data_mems_0__data_mem.data_o [25]),
    .ZN(_17831_));
 NAND2_X1 _44623_ (.A1(_17186_),
    .A2(_16805_),
    .ZN(_17832_));
 AOI21_X2 _44624_ (.A(_16544_),
    .B1(_17831_),
    .B2(_17832_),
    .ZN(_17833_));
 OAI21_X2 _44625_ (.A(_17827_),
    .B1(_17830_),
    .B2(_17833_),
    .ZN(_17834_));
 NOR2_X1 _44626_ (.A1(_17174_),
    .A2(_16867_),
    .ZN(_17835_));
 AND2_X1 _44627_ (.A1(_15606_),
    .A2(\icache.data_mems_7__data_mem.data_o [25]),
    .ZN(_17836_));
 NOR3_X2 _44628_ (.A1(_17835_),
    .A2(_17836_),
    .A3(_15932_),
    .ZN(_17837_));
 NAND2_X1 _44629_ (.A1(_16580_),
    .A2(_17180_),
    .ZN(_17838_));
 BUF_X16 _44630_ (.A(_15486_),
    .Z(_17839_));
 NAND2_X2 _44631_ (.A1(_17178_),
    .A2(_17839_),
    .ZN(_17840_));
 AOI21_X2 _44632_ (.A(_16544_),
    .B1(_17838_),
    .B2(_17840_),
    .ZN(_17841_));
 OAI21_X2 _44633_ (.A(_16013_),
    .B1(_17837_),
    .B2(_17841_),
    .ZN(_17842_));
 NAND2_X4 _44634_ (.A1(_17834_),
    .A2(_17842_),
    .ZN(_17843_));
 OAI21_X1 _44635_ (.A(_17826_),
    .B1(_17843_),
    .B2(_17757_),
    .ZN(_05232_));
 NAND2_X1 _44636_ (.A1(_17705_),
    .A2(\icache.lce.lce_cmd_inst.data_r [410]),
    .ZN(_17844_));
 INV_X1 _44637_ (.A(\icache.data_mems_4__data_mem.data_o [26]),
    .ZN(_17845_));
 NAND2_X1 _44638_ (.A1(_15491_),
    .A2(_17845_),
    .ZN(_17846_));
 NAND2_X1 _44639_ (.A1(_17201_),
    .A2(_15985_),
    .ZN(_17847_));
 AND3_X1 _44640_ (.A1(_17846_),
    .A2(_17847_),
    .A3(_15463_),
    .ZN(_17848_));
 NAND2_X1 _44641_ (.A1(_15736_),
    .A2(\icache.data_mems_6__data_mem.data_o [26]),
    .ZN(_17849_));
 NAND2_X1 _44642_ (.A1(_15606_),
    .A2(\icache.data_mems_7__data_mem.data_o [26]),
    .ZN(_17850_));
 AOI21_X2 _44643_ (.A(_16634_),
    .B1(_17849_),
    .B2(_17850_),
    .ZN(_17851_));
 OR3_X2 _44644_ (.A1(_17848_),
    .A2(_17851_),
    .A3(_15699_),
    .ZN(_17852_));
 NOR2_X2 _44645_ (.A1(_17205_),
    .A2(_15452_),
    .ZN(_17853_));
 AND2_X1 _44646_ (.A1(_15738_),
    .A2(\icache.data_mems_3__data_mem.data_o [26]),
    .ZN(_17854_));
 OAI21_X2 _44647_ (.A(_16621_),
    .B1(_17853_),
    .B2(_17854_),
    .ZN(_17855_));
 NAND2_X1 _44648_ (.A1(_15627_),
    .A2(_17211_),
    .ZN(_17856_));
 NAND2_X1 _44649_ (.A1(_17209_),
    .A2(_16112_),
    .ZN(_17857_));
 NAND3_X2 _44650_ (.A1(_17856_),
    .A2(_17857_),
    .A3(_15901_),
    .ZN(_17858_));
 NAND3_X2 _44651_ (.A1(_17855_),
    .A2(_16390_),
    .A3(_17858_),
    .ZN(_17859_));
 NAND2_X4 _44652_ (.A1(_17852_),
    .A2(_17859_),
    .ZN(_17860_));
 OAI21_X1 _44653_ (.A(_17844_),
    .B1(_17860_),
    .B2(_17757_),
    .ZN(_05234_));
 NAND2_X1 _44654_ (.A1(_17705_),
    .A2(\icache.lce.lce_cmd_inst.data_r [411]),
    .ZN(_17861_));
 NOR2_X1 _44655_ (.A1(_17224_),
    .A2(_16867_),
    .ZN(_17862_));
 AND2_X1 _44656_ (.A1(_15438_),
    .A2(\icache.data_mems_5__data_mem.data_o [27]),
    .ZN(_17863_));
 OAI21_X2 _44657_ (.A(_16865_),
    .B1(_17862_),
    .B2(_17863_),
    .ZN(_17864_));
 OR2_X1 _44658_ (.A1(_15776_),
    .A2(\icache.data_mems_6__data_mem.data_o [27]),
    .ZN(_17865_));
 NAND2_X2 _44659_ (.A1(_17219_),
    .A2(_16169_),
    .ZN(_17866_));
 NAND3_X2 _44660_ (.A1(_17865_),
    .A2(_17866_),
    .A3(_16583_),
    .ZN(_17867_));
 AOI21_X2 _44661_ (.A(_17300_),
    .B1(_17864_),
    .B2(_17867_),
    .ZN(_17868_));
 NOR2_X1 _44662_ (.A1(_17234_),
    .A2(_15452_),
    .ZN(_17869_));
 AND2_X1 _44663_ (.A1(_15738_),
    .A2(\icache.data_mems_3__data_mem.data_o [27]),
    .ZN(_17870_));
 OAI21_X2 _44664_ (.A(_17554_),
    .B1(_17869_),
    .B2(_17870_),
    .ZN(_17871_));
 OR2_X1 _44665_ (.A1(_15457_),
    .A2(\icache.data_mems_0__data_mem.data_o [27]),
    .ZN(_17872_));
 NAND2_X1 _44666_ (.A1(_17229_),
    .A2(_16112_),
    .ZN(_17873_));
 NAND3_X2 _44667_ (.A1(_17872_),
    .A2(_17873_),
    .A3(_16217_),
    .ZN(_17874_));
 AOI21_X2 _44668_ (.A(_17817_),
    .B1(_17871_),
    .B2(_17874_),
    .ZN(_17875_));
 NOR2_X4 _44669_ (.A1(_17868_),
    .A2(_17875_),
    .ZN(_17876_));
 OAI21_X1 _44670_ (.A(_17861_),
    .B1(_17876_),
    .B2(_17757_),
    .ZN(_05235_));
 BUF_X16 _44671_ (.A(_16724_),
    .Z(_17877_));
 NAND2_X1 _44672_ (.A1(_17877_),
    .A2(\icache.lce.lce_cmd_inst.data_r [412]),
    .ZN(_17878_));
 OR2_X1 _44673_ (.A1(_15714_),
    .A2(\icache.data_mems_4__data_mem.data_o [28]),
    .ZN(_17879_));
 NAND2_X1 _44674_ (.A1(_17254_),
    .A2(_16408_),
    .ZN(_17880_));
 NAND2_X1 _44675_ (.A1(_17879_),
    .A2(_17880_),
    .ZN(_17881_));
 NAND2_X1 _44676_ (.A1(_17881_),
    .A2(_15770_),
    .ZN(_17882_));
 OR2_X1 _44677_ (.A1(_15317_),
    .A2(\icache.data_mems_6__data_mem.data_o [28]),
    .ZN(_17883_));
 NAND2_X1 _44678_ (.A1(_17250_),
    .A2(_15402_),
    .ZN(_17884_));
 NAND2_X1 _44679_ (.A1(_17883_),
    .A2(_17884_),
    .ZN(_17885_));
 NAND2_X1 _44680_ (.A1(_17885_),
    .A2(_15804_),
    .ZN(_17886_));
 NAND3_X1 _44681_ (.A1(_17882_),
    .A2(_17886_),
    .A3(_15409_),
    .ZN(_17887_));
 NAND2_X1 _44682_ (.A1(_15836_),
    .A2(_17246_),
    .ZN(_17888_));
 NAND2_X1 _44683_ (.A1(_17244_),
    .A2(_15541_),
    .ZN(_17889_));
 NAND2_X1 _44684_ (.A1(_17888_),
    .A2(_17889_),
    .ZN(_17890_));
 NAND2_X1 _44685_ (.A1(_17890_),
    .A2(_17273_),
    .ZN(_17891_));
 NAND2_X1 _44686_ (.A1(_16343_),
    .A2(\icache.data_mems_0__data_mem.data_o [28]),
    .ZN(_17892_));
 NAND2_X1 _44687_ (.A1(_16083_),
    .A2(\icache.data_mems_1__data_mem.data_o [28]),
    .ZN(_17893_));
 NAND3_X1 _44688_ (.A1(_17892_),
    .A2(_15673_),
    .A3(_17893_),
    .ZN(_17894_));
 NAND3_X1 _44689_ (.A1(_17891_),
    .A2(_16372_),
    .A3(_17894_),
    .ZN(_17895_));
 AND2_X4 _44690_ (.A1(_17887_),
    .A2(_17895_),
    .ZN(_17896_));
 OAI21_X1 _44691_ (.A(_17878_),
    .B1(_17896_),
    .B2(_17757_),
    .ZN(_05236_));
 NAND2_X1 _44692_ (.A1(_17877_),
    .A2(\icache.lce.lce_cmd_inst.data_r [391]),
    .ZN(_17897_));
 NOR2_X1 _44693_ (.A1(_16793_),
    .A2(_15460_),
    .ZN(_17898_));
 AND2_X1 _44694_ (.A1(_15308_),
    .A2(\icache.data_mems_7__data_mem.data_o [7]),
    .ZN(_17899_));
 OR3_X1 _44695_ (.A1(_17898_),
    .A2(_17899_),
    .A3(_15405_),
    .ZN(_17900_));
 OR2_X1 _44696_ (.A1(_15334_),
    .A2(\icache.data_mems_4__data_mem.data_o [7]),
    .ZN(_17901_));
 NAND2_X1 _44697_ (.A1(_16788_),
    .A2(_15338_),
    .ZN(_17902_));
 NAND2_X1 _44698_ (.A1(_17901_),
    .A2(_17902_),
    .ZN(_17903_));
 NAND2_X1 _44699_ (.A1(_17903_),
    .A2(_15932_),
    .ZN(_17904_));
 AND3_X1 _44700_ (.A1(_17900_),
    .A2(_16033_),
    .A3(_17904_),
    .ZN(_17905_));
 NAND2_X1 _44701_ (.A1(_15674_),
    .A2(_16799_),
    .ZN(_17906_));
 NAND2_X2 _44702_ (.A1(_16797_),
    .A2(_15986_),
    .ZN(_17907_));
 NAND3_X2 _44703_ (.A1(_17906_),
    .A2(_17907_),
    .A3(_15988_),
    .ZN(_17908_));
 NAND2_X1 _44704_ (.A1(_16580_),
    .A2(_16804_),
    .ZN(_17909_));
 NAND2_X1 _44705_ (.A1(_16802_),
    .A2(_17839_),
    .ZN(_17910_));
 NAND3_X2 _44706_ (.A1(_17909_),
    .A2(_17910_),
    .A3(_16217_),
    .ZN(_17911_));
 AOI21_X2 _44707_ (.A(_17817_),
    .B1(_17908_),
    .B2(_17911_),
    .ZN(_17912_));
 NOR2_X4 _44708_ (.A1(_17905_),
    .A2(_17912_),
    .ZN(_17913_));
 OAI21_X1 _44709_ (.A(_17897_),
    .B1(_17913_),
    .B2(_17757_),
    .ZN(_05212_));
 NAND2_X1 _44710_ (.A1(_17877_),
    .A2(\icache.lce.lce_cmd_inst.data_r [392]),
    .ZN(_17914_));
 NOR2_X1 _44711_ (.A1(_16825_),
    .A2(_15541_),
    .ZN(_17915_));
 AND2_X1 _44712_ (.A1(_15317_),
    .A2(\icache.data_mems_7__data_mem.data_o [8]),
    .ZN(_17916_));
 NOR2_X2 _44713_ (.A1(_17915_),
    .A2(_17916_),
    .ZN(_17917_));
 NOR2_X1 _44714_ (.A1(_17917_),
    .A2(_16512_),
    .ZN(_17918_));
 NAND2_X1 _44715_ (.A1(_15719_),
    .A2(\icache.data_mems_4__data_mem.data_o [8]),
    .ZN(_17919_));
 NAND2_X1 _44716_ (.A1(_15967_),
    .A2(\icache.data_mems_5__data_mem.data_o [8]),
    .ZN(_17920_));
 AOI21_X1 _44717_ (.A(_15477_),
    .B1(_17919_),
    .B2(_17920_),
    .ZN(_17921_));
 OAI21_X1 _44718_ (.A(_16631_),
    .B1(_17918_),
    .B2(_17921_),
    .ZN(_17922_));
 NAND2_X1 _44719_ (.A1(_16155_),
    .A2(_16816_),
    .ZN(_17923_));
 NAND2_X1 _44720_ (.A1(_16814_),
    .A2(_15338_),
    .ZN(_17924_));
 AND3_X1 _44721_ (.A1(_17923_),
    .A2(_17924_),
    .A3(_16643_),
    .ZN(_17925_));
 NAND2_X1 _44722_ (.A1(_16222_),
    .A2(\icache.data_mems_0__data_mem.data_o [8]),
    .ZN(_17926_));
 NAND2_X1 _44723_ (.A1(_15725_),
    .A2(\icache.data_mems_1__data_mem.data_o [8]),
    .ZN(_17927_));
 AOI21_X2 _44724_ (.A(_16324_),
    .B1(_17926_),
    .B2(_17927_),
    .ZN(_17928_));
 OAI21_X1 _44725_ (.A(_16640_),
    .B1(_17925_),
    .B2(_17928_),
    .ZN(_17929_));
 AND2_X4 _44726_ (.A1(_17922_),
    .A2(_17929_),
    .ZN(_17930_));
 BUF_X16 _44727_ (.A(_16785_),
    .Z(_17931_));
 OAI21_X1 _44728_ (.A(_17914_),
    .B1(_17930_),
    .B2(_17931_),
    .ZN(_05213_));
 NAND2_X1 _44729_ (.A1(_17877_),
    .A2(\icache.lce.lce_cmd_inst.data_r [393]),
    .ZN(_17932_));
 OR2_X1 _44730_ (.A1(_15967_),
    .A2(\icache.data_mems_4__data_mem.data_o [9]),
    .ZN(_17933_));
 NAND2_X1 _44731_ (.A1(_16835_),
    .A2(_15728_),
    .ZN(_17934_));
 AOI21_X1 _44732_ (.A(_15379_),
    .B1(_17933_),
    .B2(_17934_),
    .ZN(_17935_));
 OR2_X1 _44733_ (.A1(_15573_),
    .A2(\icache.data_mems_6__data_mem.data_o [9]),
    .ZN(_17936_));
 NAND2_X1 _44734_ (.A1(_16831_),
    .A2(_15752_),
    .ZN(_17937_));
 AOI21_X2 _44735_ (.A(_16005_),
    .B1(_17936_),
    .B2(_17937_),
    .ZN(_17938_));
 OAI21_X2 _44736_ (.A(_17582_),
    .B1(_17935_),
    .B2(_17938_),
    .ZN(_17939_));
 NAND2_X1 _44737_ (.A1(_15674_),
    .A2(_16847_),
    .ZN(_17940_));
 NAND2_X1 _44738_ (.A1(_16845_),
    .A2(_15986_),
    .ZN(_17941_));
 AOI21_X2 _44739_ (.A(_16014_),
    .B1(_17940_),
    .B2(_17941_),
    .ZN(_17942_));
 NAND2_X1 _44740_ (.A1(_16580_),
    .A2(_16842_),
    .ZN(_17943_));
 NAND2_X1 _44741_ (.A1(_16840_),
    .A2(_17839_),
    .ZN(_17944_));
 AOI21_X2 _44742_ (.A(_17016_),
    .B1(_17943_),
    .B2(_17944_),
    .ZN(_17945_));
 OAI21_X2 _44743_ (.A(_17500_),
    .B1(_17942_),
    .B2(_17945_),
    .ZN(_17946_));
 NAND2_X4 _44744_ (.A1(_17939_),
    .A2(_17946_),
    .ZN(_17947_));
 OAI21_X1 _44745_ (.A(_17932_),
    .B1(_17947_),
    .B2(_17931_),
    .ZN(_05214_));
 NAND2_X1 _44746_ (.A1(_17877_),
    .A2(\icache.lce.lce_cmd_inst.data_r [314]),
    .ZN(_17948_));
 NAND2_X1 _44747_ (.A1(_16536_),
    .A2(_15770_),
    .ZN(_17949_));
 NAND2_X1 _44748_ (.A1(_16532_),
    .A2(_15514_),
    .ZN(_17950_));
 AOI21_X1 _44749_ (.A(_15686_),
    .B1(_17949_),
    .B2(_17950_),
    .ZN(_17951_));
 AND3_X1 _44750_ (.A1(_16545_),
    .A2(_16546_),
    .A3(_16229_),
    .ZN(_17952_));
 AOI21_X2 _44751_ (.A(_15664_),
    .B1(_16540_),
    .B2(_16542_),
    .ZN(_17953_));
 NOR3_X1 _44752_ (.A1(_17952_),
    .A2(_17953_),
    .A3(_15597_),
    .ZN(_17954_));
 OR2_X4 _44753_ (.A1(_17951_),
    .A2(_17954_),
    .ZN(_17955_));
 OAI21_X1 _44754_ (.A(_17948_),
    .B1(_17955_),
    .B2(_17931_),
    .ZN(_05127_));
 NAND2_X1 _44755_ (.A1(_17877_),
    .A2(\icache.lce.lce_cmd_inst.data_r [315]),
    .ZN(_17956_));
 OR3_X2 _44756_ (.A1(_16566_),
    .A2(_16567_),
    .A3(_15394_),
    .ZN(_17957_));
 OR3_X2 _44757_ (.A1(_16570_),
    .A2(_16571_),
    .A3(_15405_),
    .ZN(_17958_));
 NAND2_X4 _44758_ (.A1(_17957_),
    .A2(_17958_),
    .ZN(_17959_));
 BUF_X16 _44759_ (.A(_16265_),
    .Z(_17960_));
 NAND2_X1 _44760_ (.A1(_17959_),
    .A2(_17960_),
    .ZN(_17961_));
 NAND2_X1 _44761_ (.A1(_16554_),
    .A2(_15567_),
    .ZN(_17962_));
 NAND2_X1 _44762_ (.A1(_16560_),
    .A2(_15576_),
    .ZN(_17963_));
 NAND2_X4 _44763_ (.A1(_17962_),
    .A2(_17963_),
    .ZN(_17964_));
 NAND2_X1 _44764_ (.A1(_17964_),
    .A2(_17567_),
    .ZN(_17965_));
 NAND2_X4 _44765_ (.A1(_17961_),
    .A2(_17965_),
    .ZN(_17966_));
 OAI21_X1 _44766_ (.A(_17956_),
    .B1(_17966_),
    .B2(_17931_),
    .ZN(_05128_));
 NAND2_X1 _44767_ (.A1(_17877_),
    .A2(\icache.lce.lce_cmd_inst.data_r [316]),
    .ZN(_17967_));
 AOI21_X4 _44768_ (.A(_15576_),
    .B1(_16586_),
    .B2(_16587_),
    .ZN(_17968_));
 AOI21_X4 _44769_ (.A(_16544_),
    .B1(_16590_),
    .B2(_16591_),
    .ZN(_17969_));
 OAI21_X2 _44770_ (.A(_17827_),
    .B1(_17968_),
    .B2(_17969_),
    .ZN(_17970_));
 BUF_X16 _44771_ (.A(_16012_),
    .Z(_17971_));
 AOI21_X4 _44772_ (.A(_15576_),
    .B1(_16576_),
    .B2(_16577_),
    .ZN(_17972_));
 AOI21_X4 _44773_ (.A(_16544_),
    .B1(_16581_),
    .B2(_16582_),
    .ZN(_17973_));
 OAI21_X2 _44774_ (.A(_17971_),
    .B1(_17972_),
    .B2(_17973_),
    .ZN(_17974_));
 NAND2_X4 _44775_ (.A1(_17970_),
    .A2(_17974_),
    .ZN(_17975_));
 OAI21_X1 _44776_ (.A(_17967_),
    .B1(_17975_),
    .B2(_17931_),
    .ZN(_05129_));
 NAND2_X1 _44777_ (.A1(_17877_),
    .A2(\icache.lce.lce_cmd_inst.data_r [317]),
    .ZN(_17976_));
 OR3_X1 _44778_ (.A1(_16597_),
    .A2(_16598_),
    .A3(_16226_),
    .ZN(_17977_));
 NAND2_X1 _44779_ (.A1(_16602_),
    .A2(_16347_),
    .ZN(_17978_));
 NAND2_X1 _44780_ (.A1(_17977_),
    .A2(_17978_),
    .ZN(_17979_));
 NAND2_X2 _44781_ (.A1(_17979_),
    .A2(_17960_),
    .ZN(_17980_));
 BUF_X16 _44782_ (.A(_15405_),
    .Z(_17981_));
 NOR3_X1 _44783_ (.A1(_16605_),
    .A2(_16606_),
    .A3(_17981_),
    .ZN(_17982_));
 AOI21_X2 _44784_ (.A(_16544_),
    .B1(_16608_),
    .B2(_16609_),
    .ZN(_17983_));
 OAI21_X2 _44785_ (.A(_17500_),
    .B1(_17982_),
    .B2(_17983_),
    .ZN(_17984_));
 NAND2_X4 _44786_ (.A1(_17980_),
    .A2(_17984_),
    .ZN(_17985_));
 OAI21_X1 _44787_ (.A(_17976_),
    .B1(_17985_),
    .B2(_17931_),
    .ZN(_05130_));
 NAND2_X1 _44788_ (.A1(_17877_),
    .A2(\icache.lce.lce_cmd_inst.data_r [318]),
    .ZN(_17986_));
 NOR3_X2 _44789_ (.A1(_16622_),
    .A2(_16623_),
    .A3(_17273_),
    .ZN(_17987_));
 BUF_X16 _44790_ (.A(_15405_),
    .Z(_17988_));
 AOI21_X2 _44791_ (.A(_17988_),
    .B1(_16625_),
    .B2(_16626_),
    .ZN(_17989_));
 BUF_X16 _44792_ (.A(_15833_),
    .Z(_17990_));
 NOR3_X2 _44793_ (.A1(_17987_),
    .A2(_17989_),
    .A3(_17990_),
    .ZN(_17991_));
 OAI21_X2 _44794_ (.A(_15450_),
    .B1(_16614_),
    .B2(_16615_),
    .ZN(_17992_));
 NAND3_X2 _44795_ (.A1(_16617_),
    .A2(_16618_),
    .A3(_15994_),
    .ZN(_17993_));
 AOI21_X2 _44796_ (.A(_17817_),
    .B1(_17992_),
    .B2(_17993_),
    .ZN(_17994_));
 NOR2_X4 _44797_ (.A1(_17991_),
    .A2(_17994_),
    .ZN(_17995_));
 OAI21_X1 _44798_ (.A(_17986_),
    .B1(_17995_),
    .B2(_17931_),
    .ZN(_05131_));
 NAND2_X1 _44799_ (.A1(_17877_),
    .A2(\icache.lce.lce_cmd_inst.data_r [319]),
    .ZN(_17996_));
 AND3_X1 _44800_ (.A1(_16632_),
    .A2(_16633_),
    .A3(_15378_),
    .ZN(_17997_));
 AOI21_X1 _44801_ (.A(_15331_),
    .B1(_16636_),
    .B2(_16637_),
    .ZN(_17998_));
 OR3_X2 _44802_ (.A1(_17997_),
    .A2(_15734_),
    .A3(_17998_),
    .ZN(_17999_));
 AND3_X1 _44803_ (.A1(_16645_),
    .A2(_16541_),
    .A3(_16646_),
    .ZN(_18000_));
 AOI21_X2 _44804_ (.A(_16544_),
    .B1(_16641_),
    .B2(_16642_),
    .ZN(_18001_));
 OAI21_X2 _44805_ (.A(_17500_),
    .B1(_18000_),
    .B2(_18001_),
    .ZN(_18002_));
 NAND2_X4 _44806_ (.A1(_17999_),
    .A2(_18002_),
    .ZN(_18003_));
 OAI21_X1 _44807_ (.A(_17996_),
    .B1(_18003_),
    .B2(_17931_),
    .ZN(_05132_));
 BUF_X8 _44808_ (.A(_16724_),
    .Z(_18004_));
 NAND2_X1 _44809_ (.A1(_18004_),
    .A2(\icache.lce.lce_cmd_inst.data_r [320]),
    .ZN(_18005_));
 NOR2_X1 _44810_ (.A1(_15554_),
    .A2(\icache.data_mems_4__data_mem.data_o [0]),
    .ZN(_18006_));
 AOI211_X2 _44811_ (.A(_16226_),
    .B(_18006_),
    .C1(_15756_),
    .C2(_16662_),
    .ZN(_18007_));
 AOI21_X2 _44812_ (.A(_15812_),
    .B1(_16658_),
    .B2(_16659_),
    .ZN(_18008_));
 OR3_X2 _44813_ (.A1(_18007_),
    .A2(_18008_),
    .A3(_15699_),
    .ZN(_18009_));
 AOI21_X1 _44814_ (.A(_15544_),
    .B1(_16651_),
    .B2(_16652_),
    .ZN(_18010_));
 AOI21_X1 _44815_ (.A(_17068_),
    .B1(_16654_),
    .B2(_16655_),
    .ZN(_18011_));
 OAI21_X2 _44816_ (.A(_17500_),
    .B1(_18010_),
    .B2(_18011_),
    .ZN(_18012_));
 NAND2_X4 _44817_ (.A1(_18009_),
    .A2(_18012_),
    .ZN(_18013_));
 OAI21_X1 _44818_ (.A(_18005_),
    .B1(_18013_),
    .B2(_17931_),
    .ZN(_05134_));
 NAND2_X1 _44819_ (.A1(_18004_),
    .A2(\icache.lce.lce_cmd_inst.data_r [321]),
    .ZN(_18014_));
 OR3_X1 _44820_ (.A1(_16675_),
    .A2(_16676_),
    .A3(_16321_),
    .ZN(_18015_));
 OR3_X2 _44821_ (.A1(_16679_),
    .A2(_16680_),
    .A3(_17068_),
    .ZN(_18016_));
 AOI21_X1 _44822_ (.A(_16049_),
    .B1(_18015_),
    .B2(_18016_),
    .ZN(_18017_));
 OAI21_X1 _44823_ (.A(_16327_),
    .B1(_16668_),
    .B2(_16669_),
    .ZN(_18018_));
 INV_X1 _44824_ (.A(\icache.data_mems_6__data_mem.data_o [1]),
    .ZN(_18019_));
 NAND2_X1 _44825_ (.A1(_18019_),
    .A2(_15495_),
    .ZN(_18020_));
 OAI211_X4 _44826_ (.A(_18020_),
    .B(_15609_),
    .C1(_15725_),
    .C2(\icache.data_mems_7__data_mem.data_o [1]),
    .ZN(_18021_));
 AND3_X1 _44827_ (.A1(_18018_),
    .A2(_18021_),
    .A3(_15819_),
    .ZN(_18022_));
 OR2_X4 _44828_ (.A1(_18017_),
    .A2(_18022_),
    .ZN(_18023_));
 OAI21_X1 _44829_ (.A(_18014_),
    .B1(_18023_),
    .B2(_17931_),
    .ZN(_05135_));
 NAND2_X1 _44830_ (.A1(_18004_),
    .A2(\icache.lce.lce_cmd_inst.data_r [322]),
    .ZN(_18024_));
 NOR3_X2 _44831_ (.A1(_16694_),
    .A2(_16695_),
    .A3(_17273_),
    .ZN(_18025_));
 AOI21_X2 _44832_ (.A(_17988_),
    .B1(_16697_),
    .B2(_16699_),
    .ZN(_18026_));
 OAI21_X1 _44833_ (.A(_17582_),
    .B1(_18025_),
    .B2(_18026_),
    .ZN(_18027_));
 OAI21_X2 _44834_ (.A(_17308_),
    .B1(_16686_),
    .B2(_16687_),
    .ZN(_18028_));
 NAND2_X1 _44835_ (.A1(_16690_),
    .A2(_17839_),
    .ZN(_18029_));
 OAI211_X4 _44836_ (.A(_18029_),
    .B(_15779_),
    .C1(_15324_),
    .C2(\icache.data_mems_1__data_mem.data_o [2]),
    .ZN(_18030_));
 NAND3_X1 _44837_ (.A1(_18028_),
    .A2(_18030_),
    .A3(_15996_),
    .ZN(_18031_));
 NAND2_X2 _44838_ (.A1(_18027_),
    .A2(_18031_),
    .ZN(_18032_));
 BUF_X4 _44839_ (.A(_16785_),
    .Z(_18033_));
 OAI21_X1 _44840_ (.A(_18024_),
    .B1(_18032_),
    .B2(_18033_),
    .ZN(_05136_));
 NAND2_X1 _44841_ (.A1(_18004_),
    .A2(\icache.lce.lce_cmd_inst.data_r [323]),
    .ZN(_18034_));
 OR3_X2 _44842_ (.A1(_16705_),
    .A2(_16706_),
    .A3(_16053_),
    .ZN(_18035_));
 NAND2_X1 _44843_ (.A1(_16711_),
    .A2(_15406_),
    .ZN(_18036_));
 AND3_X1 _44844_ (.A1(_18035_),
    .A2(_16033_),
    .A3(_18036_),
    .ZN(_18037_));
 OAI21_X1 _44845_ (.A(_15484_),
    .B1(_16715_),
    .B2(_16716_),
    .ZN(_18038_));
 OAI21_X2 _44846_ (.A(_15497_),
    .B1(_16719_),
    .B2(_16720_),
    .ZN(_18039_));
 AOI21_X1 _44847_ (.A(_17817_),
    .B1(_18038_),
    .B2(_18039_),
    .ZN(_18040_));
 NOR2_X2 _44848_ (.A1(_18037_),
    .A2(_18040_),
    .ZN(_18041_));
 OAI21_X1 _44849_ (.A(_18034_),
    .B1(_18041_),
    .B2(_18033_),
    .ZN(_05137_));
 NAND2_X1 _44850_ (.A1(_18004_),
    .A2(\icache.lce.lce_cmd_inst.data_r [324]),
    .ZN(_18042_));
 NOR3_X1 _44851_ (.A1(_16728_),
    .A2(_16729_),
    .A3(_15619_),
    .ZN(_18043_));
 AOI21_X2 _44852_ (.A(_16005_),
    .B1(_16731_),
    .B2(_16733_),
    .ZN(_18044_));
 OAI21_X1 _44853_ (.A(_17582_),
    .B1(_18043_),
    .B2(_18044_),
    .ZN(_18045_));
 AOI21_X2 _44854_ (.A(_16014_),
    .B1(_16736_),
    .B2(_16738_),
    .ZN(_18046_));
 AOI21_X1 _44855_ (.A(_17016_),
    .B1(_16741_),
    .B2(_16743_),
    .ZN(_18047_));
 OAI21_X1 _44856_ (.A(_17500_),
    .B1(_18046_),
    .B2(_18047_),
    .ZN(_18048_));
 NAND2_X2 _44857_ (.A1(_18045_),
    .A2(_18048_),
    .ZN(_18049_));
 OAI21_X1 _44858_ (.A(_18042_),
    .B1(_18049_),
    .B2(_18033_),
    .ZN(_05138_));
 NAND2_X1 _44859_ (.A1(_18004_),
    .A2(\icache.lce.lce_cmd_inst.data_r [325]),
    .ZN(_18050_));
 OR3_X2 _44860_ (.A1(_16748_),
    .A2(_16749_),
    .A3(_16053_),
    .ZN(_18051_));
 NAND2_X1 _44861_ (.A1(_16755_),
    .A2(_15406_),
    .ZN(_18052_));
 AOI21_X2 _44862_ (.A(_15686_),
    .B1(_18051_),
    .B2(_18052_),
    .ZN(_18053_));
 OAI21_X1 _44863_ (.A(_15484_),
    .B1(_16758_),
    .B2(_16759_),
    .ZN(_18054_));
 NAND3_X1 _44864_ (.A1(_16761_),
    .A2(_16763_),
    .A3(_15378_),
    .ZN(_18055_));
 AND3_X1 _44865_ (.A1(_18054_),
    .A2(_15430_),
    .A3(_18055_),
    .ZN(_18056_));
 OR2_X4 _44866_ (.A1(_18053_),
    .A2(_18056_),
    .ZN(_18057_));
 OAI21_X1 _44867_ (.A(_18050_),
    .B1(_18057_),
    .B2(_18033_),
    .ZN(_05139_));
 NAND2_X1 _44868_ (.A1(_18004_),
    .A2(\icache.lce.lce_cmd_inst.data_r [326]),
    .ZN(_18058_));
 OAI21_X4 _44869_ (.A(_15708_),
    .B1(_16768_),
    .B2(_16769_),
    .ZN(_18059_));
 OAI21_X4 _44870_ (.A(_15712_),
    .B1(_16771_),
    .B2(_16772_),
    .ZN(_18060_));
 AOI21_X4 _44871_ (.A(_17300_),
    .B1(_18059_),
    .B2(_18060_),
    .ZN(_18061_));
 OAI21_X2 _44872_ (.A(_17554_),
    .B1(_16776_),
    .B2(_16777_),
    .ZN(_18062_));
 NAND3_X2 _44873_ (.A1(_16779_),
    .A2(_16781_),
    .A3(_16217_),
    .ZN(_18063_));
 AOI21_X2 _44874_ (.A(_17817_),
    .B1(_18062_),
    .B2(_18063_),
    .ZN(_18064_));
 NOR2_X4 _44875_ (.A1(_18061_),
    .A2(_18064_),
    .ZN(_18065_));
 OAI21_X1 _44876_ (.A(_18058_),
    .B1(_18065_),
    .B2(_18033_),
    .ZN(_05140_));
 NAND2_X1 _44877_ (.A1(_18004_),
    .A2(\icache.lce.lce_cmd_inst.data_r [327]),
    .ZN(_18066_));
 NOR3_X2 _44878_ (.A1(_16789_),
    .A2(_16790_),
    .A3(_16227_),
    .ZN(_18067_));
 AOI21_X1 _44879_ (.A(_17710_),
    .B1(_16792_),
    .B2(_16794_),
    .ZN(_18068_));
 OAI21_X1 _44880_ (.A(_17582_),
    .B1(_18067_),
    .B2(_18068_),
    .ZN(_18069_));
 AOI21_X2 _44881_ (.A(_16014_),
    .B1(_16798_),
    .B2(_16800_),
    .ZN(_18070_));
 AOI21_X2 _44882_ (.A(_17016_),
    .B1(_16803_),
    .B2(_16806_),
    .ZN(_18071_));
 OAI21_X1 _44883_ (.A(_17500_),
    .B1(_18070_),
    .B2(_18071_),
    .ZN(_18072_));
 NAND2_X2 _44884_ (.A1(_18069_),
    .A2(_18072_),
    .ZN(_18073_));
 OAI21_X1 _44885_ (.A(_18066_),
    .B1(_18073_),
    .B2(_18033_),
    .ZN(_05141_));
 NAND2_X1 _44886_ (.A1(_18004_),
    .A2(\icache.lce.lce_cmd_inst.data_r [328]),
    .ZN(_18074_));
 NOR3_X2 _44887_ (.A1(_16820_),
    .A2(_16821_),
    .A3(_16512_),
    .ZN(_18075_));
 AOI21_X2 _44888_ (.A(_17710_),
    .B1(_16824_),
    .B2(_16826_),
    .ZN(_18076_));
 OAI21_X1 _44889_ (.A(_17582_),
    .B1(_18075_),
    .B2(_18076_),
    .ZN(_18077_));
 OAI21_X1 _44890_ (.A(_16621_),
    .B1(_16811_),
    .B2(_16812_),
    .ZN(_18078_));
 NAND3_X4 _44891_ (.A1(_16815_),
    .A2(_16817_),
    .A3(_15901_),
    .ZN(_18079_));
 NAND3_X1 _44892_ (.A1(_18078_),
    .A2(_16390_),
    .A3(_18079_),
    .ZN(_18080_));
 NAND2_X2 _44893_ (.A1(_18077_),
    .A2(_18080_),
    .ZN(_18081_));
 OAI21_X1 _44894_ (.A(_18074_),
    .B1(_18081_),
    .B2(_18033_),
    .ZN(_05142_));
 NAND2_X1 _44895_ (.A1(_18004_),
    .A2(\icache.lce.lce_cmd_inst.data_r [329]),
    .ZN(_18082_));
 AOI21_X2 _44896_ (.A(_17710_),
    .B1(_16841_),
    .B2(_16843_),
    .ZN(_18083_));
 AOI21_X2 _44897_ (.A(_17988_),
    .B1(_16846_),
    .B2(_16848_),
    .ZN(_18084_));
 BUF_X16 _44898_ (.A(_15408_),
    .Z(_18085_));
 NOR3_X2 _44899_ (.A1(_18083_),
    .A2(_18084_),
    .A3(_18085_),
    .ZN(_18086_));
 OAI21_X4 _44900_ (.A(_15450_),
    .B1(_16836_),
    .B2(_16837_),
    .ZN(_18087_));
 OAI21_X2 _44901_ (.A(_15650_),
    .B1(_16832_),
    .B2(_16833_),
    .ZN(_18088_));
 AOI21_X2 _44902_ (.A(_17517_),
    .B1(_18087_),
    .B2(_18088_),
    .ZN(_18089_));
 NOR2_X4 _44903_ (.A1(_18086_),
    .A2(_18089_),
    .ZN(_18090_));
 OAI21_X1 _44904_ (.A(_18082_),
    .B1(_18090_),
    .B2(_18033_),
    .ZN(_05143_));
 BUF_X4 _44905_ (.A(_16724_),
    .Z(_18091_));
 NAND2_X1 _44906_ (.A1(_18091_),
    .A2(\icache.lce.lce_cmd_inst.data_r [330]),
    .ZN(_18092_));
 NAND2_X1 _44907_ (.A1(_16856_),
    .A2(_16256_),
    .ZN(_18093_));
 NAND2_X1 _44908_ (.A1(_16862_),
    .A2(_16262_),
    .ZN(_18094_));
 NAND2_X1 _44909_ (.A1(_18093_),
    .A2(_18094_),
    .ZN(_18095_));
 NAND2_X2 _44910_ (.A1(_18095_),
    .A2(_17731_),
    .ZN(_18096_));
 NOR3_X2 _44911_ (.A1(_16868_),
    .A2(_16869_),
    .A3(_17981_),
    .ZN(_18097_));
 AOI21_X1 _44912_ (.A(_15740_),
    .B1(_16871_),
    .B2(_16873_),
    .ZN(_18098_));
 OAI21_X1 _44913_ (.A(_17971_),
    .B1(_18097_),
    .B2(_18098_),
    .ZN(_18099_));
 NAND2_X4 _44914_ (.A1(_18096_),
    .A2(_18099_),
    .ZN(_18100_));
 OAI21_X1 _44915_ (.A(_18092_),
    .B1(_18100_),
    .B2(_18033_),
    .ZN(_05145_));
 NAND2_X1 _44916_ (.A1(_18091_),
    .A2(\icache.lce.lce_cmd_inst.data_r [331]),
    .ZN(_18101_));
 NOR3_X1 _44917_ (.A1(_16886_),
    .A2(_16887_),
    .A3(_16195_),
    .ZN(_18102_));
 AOI21_X1 _44918_ (.A(_15938_),
    .B1(_16890_),
    .B2(_16892_),
    .ZN(_18103_));
 OAI21_X1 _44919_ (.A(_17827_),
    .B1(_18102_),
    .B2(_18103_),
    .ZN(_18104_));
 OAI21_X2 _44920_ (.A(_15450_),
    .B1(_16879_),
    .B2(_16880_),
    .ZN(_18105_));
 NAND2_X1 _44921_ (.A1(_17586_),
    .A2(_17839_),
    .ZN(_18106_));
 OAI211_X4 _44922_ (.A(_18106_),
    .B(_17981_),
    .C1(_15324_),
    .C2(\icache.data_mems_7__data_mem.data_o [11]),
    .ZN(_18107_));
 NAND3_X2 _44923_ (.A1(_18105_),
    .A2(_18107_),
    .A3(_15656_),
    .ZN(_18108_));
 NAND2_X2 _44924_ (.A1(_18104_),
    .A2(_18108_),
    .ZN(_18109_));
 OAI21_X1 _44925_ (.A(_18101_),
    .B1(_18109_),
    .B2(_18033_),
    .ZN(_05146_));
 NAND2_X1 _44926_ (.A1(_18091_),
    .A2(\icache.lce.lce_cmd_inst.data_r [332]),
    .ZN(_18110_));
 NOR3_X2 _44927_ (.A1(_16904_),
    .A2(_16905_),
    .A3(_17273_),
    .ZN(_18111_));
 AOI21_X2 _44928_ (.A(_17988_),
    .B1(_16908_),
    .B2(_16910_),
    .ZN(_18112_));
 NOR3_X1 _44929_ (.A1(_18111_),
    .A2(_18112_),
    .A3(_18085_),
    .ZN(_18113_));
 OAI21_X1 _44930_ (.A(_15450_),
    .B1(_16897_),
    .B2(_16898_),
    .ZN(_18114_));
 NAND2_X1 _44931_ (.A1(_16901_),
    .A2(_17839_),
    .ZN(_18115_));
 BUF_X16 _44932_ (.A(_15511_),
    .Z(_18116_));
 OAI211_X4 _44933_ (.A(_18115_),
    .B(_15932_),
    .C1(_18116_),
    .C2(\icache.data_mems_7__data_mem.data_o [12]),
    .ZN(_18117_));
 AOI21_X1 _44934_ (.A(_17517_),
    .B1(_18114_),
    .B2(_18117_),
    .ZN(_18118_));
 NOR2_X2 _44935_ (.A1(_18113_),
    .A2(_18118_),
    .ZN(_18119_));
 BUF_X8 _44936_ (.A(_16785_),
    .Z(_18120_));
 OAI21_X1 _44937_ (.A(_18110_),
    .B1(_18119_),
    .B2(_18120_),
    .ZN(_05147_));
 NAND2_X1 _44938_ (.A1(_18091_),
    .A2(\icache.lce.lce_cmd_inst.data_r [333]),
    .ZN(_18121_));
 NOR3_X1 _44939_ (.A1(_16915_),
    .A2(_16916_),
    .A3(_15619_),
    .ZN(_18122_));
 AOI21_X2 _44940_ (.A(_16005_),
    .B1(_16919_),
    .B2(_16921_),
    .ZN(_18123_));
 OAI21_X1 _44941_ (.A(_17827_),
    .B1(_18122_),
    .B2(_18123_),
    .ZN(_18124_));
 OAI21_X2 _44942_ (.A(_16386_),
    .B1(_16925_),
    .B2(_16926_),
    .ZN(_18125_));
 NAND3_X2 _44943_ (.A1(_16929_),
    .A2(_16931_),
    .A3(_16396_),
    .ZN(_18126_));
 NAND3_X1 _44944_ (.A1(_18125_),
    .A2(_16823_),
    .A3(_18126_),
    .ZN(_18127_));
 NAND2_X2 _44945_ (.A1(_18124_),
    .A2(_18127_),
    .ZN(_18128_));
 OAI21_X1 _44946_ (.A(_18121_),
    .B1(_18128_),
    .B2(_18120_),
    .ZN(_05148_));
 NAND2_X1 _44947_ (.A1(_18091_),
    .A2(\icache.lce.lce_cmd_inst.data_r [334]),
    .ZN(_18129_));
 NOR3_X2 _44948_ (.A1(_16946_),
    .A2(_16947_),
    .A3(_15938_),
    .ZN(_18130_));
 AOI21_X4 _44949_ (.A(_17264_),
    .B1(_16949_),
    .B2(_16951_),
    .ZN(_18131_));
 BUF_X16 _44950_ (.A(_15833_),
    .Z(_18132_));
 NOR3_X1 _44951_ (.A1(_18130_),
    .A2(_18131_),
    .A3(_18132_),
    .ZN(_18133_));
 OAI21_X2 _44952_ (.A(_17554_),
    .B1(_16937_),
    .B2(_16938_),
    .ZN(_18134_));
 OAI21_X2 _44953_ (.A(_15650_),
    .B1(_16941_),
    .B2(_16942_),
    .ZN(_18135_));
 AOI21_X1 _44954_ (.A(_17817_),
    .B1(_18134_),
    .B2(_18135_),
    .ZN(_18136_));
 NOR2_X2 _44955_ (.A1(_18133_),
    .A2(_18136_),
    .ZN(_18137_));
 OAI21_X1 _44956_ (.A(_18129_),
    .B1(_18137_),
    .B2(_18120_),
    .ZN(_05149_));
 NAND2_X1 _44957_ (.A1(_18091_),
    .A2(\icache.lce.lce_cmd_inst.data_r [335]),
    .ZN(_18138_));
 OR3_X1 _44958_ (.A1(_16958_),
    .A2(_16959_),
    .A3(_16321_),
    .ZN(_18139_));
 OR3_X2 _44959_ (.A1(_16962_),
    .A2(_16963_),
    .A3(_17068_),
    .ZN(_18140_));
 AOI21_X1 _44960_ (.A(_16049_),
    .B1(_18139_),
    .B2(_18140_),
    .ZN(_18141_));
 OAI21_X1 _44961_ (.A(_16327_),
    .B1(_16967_),
    .B2(_16968_),
    .ZN(_18142_));
 NAND3_X1 _44962_ (.A1(_16971_),
    .A2(_16973_),
    .A3(_15342_),
    .ZN(_18143_));
 AND3_X1 _44963_ (.A1(_18142_),
    .A2(_15522_),
    .A3(_18143_),
    .ZN(_18144_));
 OR2_X2 _44964_ (.A1(_18141_),
    .A2(_18144_),
    .ZN(_18145_));
 OAI21_X1 _44965_ (.A(_18138_),
    .B1(_18145_),
    .B2(_18120_),
    .ZN(_05150_));
 NAND2_X1 _44966_ (.A1(_18091_),
    .A2(\icache.lce.lce_cmd_inst.data_r [336]),
    .ZN(_18146_));
 NOR3_X2 _44967_ (.A1(_16978_),
    .A2(_16979_),
    .A3(_16512_),
    .ZN(_18147_));
 AOI21_X2 _44968_ (.A(_17710_),
    .B1(_16982_),
    .B2(_16984_),
    .ZN(_18148_));
 OAI21_X1 _44969_ (.A(_17582_),
    .B1(_18147_),
    .B2(_18148_),
    .ZN(_18149_));
 NOR3_X2 _44970_ (.A1(_16988_),
    .A2(_16989_),
    .A3(_17981_),
    .ZN(_18150_));
 AOI21_X2 _44971_ (.A(_15740_),
    .B1(_16991_),
    .B2(_16993_),
    .ZN(_18151_));
 OAI21_X1 _44972_ (.A(_17500_),
    .B1(_18150_),
    .B2(_18151_),
    .ZN(_18152_));
 NAND2_X2 _44973_ (.A1(_18149_),
    .A2(_18152_),
    .ZN(_18153_));
 OAI21_X1 _44974_ (.A(_18146_),
    .B1(_18153_),
    .B2(_18120_),
    .ZN(_05151_));
 NAND2_X1 _44975_ (.A1(_18091_),
    .A2(\icache.lce.lce_cmd_inst.data_r [337]),
    .ZN(_18154_));
 NAND2_X2 _44976_ (.A1(_17002_),
    .A2(_16021_),
    .ZN(_18155_));
 NAND2_X2 _44977_ (.A1(_17008_),
    .A2(_15804_),
    .ZN(_18156_));
 AND3_X2 _44978_ (.A1(_18155_),
    .A2(_18156_),
    .A3(_16562_),
    .ZN(_18157_));
 OAI21_X1 _44979_ (.A(_16327_),
    .B1(_17013_),
    .B2(_17014_),
    .ZN(_18158_));
 NAND3_X1 _44980_ (.A1(_17017_),
    .A2(_17019_),
    .A3(_15342_),
    .ZN(_18159_));
 AOI21_X2 _44981_ (.A(_17517_),
    .B1(_18158_),
    .B2(_18159_),
    .ZN(_18160_));
 NOR2_X4 _44982_ (.A1(_18157_),
    .A2(_18160_),
    .ZN(_18161_));
 OAI21_X1 _44983_ (.A(_18154_),
    .B1(_18161_),
    .B2(_18120_),
    .ZN(_05152_));
 NAND2_X1 _44984_ (.A1(_18091_),
    .A2(\icache.lce.lce_cmd_inst.data_r [338]),
    .ZN(_18162_));
 NOR3_X2 _44985_ (.A1(_17024_),
    .A2(_17025_),
    .A3(_15619_),
    .ZN(_18163_));
 BUF_X16 _44986_ (.A(_15609_),
    .Z(_18164_));
 AOI21_X4 _44987_ (.A(_18164_),
    .B1(_17028_),
    .B2(_17030_),
    .ZN(_18165_));
 OAI21_X1 _44988_ (.A(_17582_),
    .B1(_18163_),
    .B2(_18165_),
    .ZN(_18166_));
 OAI21_X2 _44989_ (.A(_16386_),
    .B1(_17034_),
    .B2(_17035_),
    .ZN(_18167_));
 NAND3_X2 _44990_ (.A1(_17038_),
    .A2(_17040_),
    .A3(_16396_),
    .ZN(_18168_));
 NAND3_X1 _44991_ (.A1(_18167_),
    .A2(_16390_),
    .A3(_18168_),
    .ZN(_18169_));
 NAND2_X2 _44992_ (.A1(_18166_),
    .A2(_18169_),
    .ZN(_18170_));
 OAI21_X1 _44993_ (.A(_18162_),
    .B1(_18170_),
    .B2(_18120_),
    .ZN(_05153_));
 NAND2_X1 _44994_ (.A1(_18091_),
    .A2(\icache.lce.lce_cmd_inst.data_r [339]),
    .ZN(_18171_));
 NOR3_X1 _44995_ (.A1(_17045_),
    .A2(_17046_),
    .A3(_16512_),
    .ZN(_18172_));
 AOI21_X2 _44996_ (.A(_17710_),
    .B1(_17048_),
    .B2(_17050_),
    .ZN(_18173_));
 OAI21_X1 _44997_ (.A(_17827_),
    .B1(_18172_),
    .B2(_18173_),
    .ZN(_18174_));
 AOI21_X1 _44998_ (.A(_16014_),
    .B1(_17054_),
    .B2(_17056_),
    .ZN(_18175_));
 AOI21_X1 _44999_ (.A(_17016_),
    .B1(_17059_),
    .B2(_17061_),
    .ZN(_18176_));
 OAI21_X1 _45000_ (.A(_17971_),
    .B1(_18175_),
    .B2(_18176_),
    .ZN(_18177_));
 NAND2_X2 _45001_ (.A1(_18174_),
    .A2(_18177_),
    .ZN(_18178_));
 OAI21_X1 _45002_ (.A(_18171_),
    .B1(_18178_),
    .B2(_18120_),
    .ZN(_05154_));
 BUF_X4 _45003_ (.A(_16724_),
    .Z(_18179_));
 NAND2_X1 _45004_ (.A1(_18179_),
    .A2(\icache.lce.lce_cmd_inst.data_r [340]),
    .ZN(_18180_));
 NAND2_X1 _45005_ (.A1(_17077_),
    .A2(_15545_),
    .ZN(_18181_));
 NAND2_X1 _45006_ (.A1(_17083_),
    .A2(_17988_),
    .ZN(_18182_));
 AND3_X1 _45007_ (.A1(_18181_),
    .A2(_18182_),
    .A3(_15940_),
    .ZN(_18183_));
 OAI21_X1 _45008_ (.A(_15660_),
    .B1(_17066_),
    .B2(_17067_),
    .ZN(_18184_));
 OR2_X1 _45009_ (.A1(_15488_),
    .A2(\icache.data_mems_1__data_mem.data_o [20]),
    .ZN(_18185_));
 OAI211_X2 _45010_ (.A(_18185_),
    .B(_16229_),
    .C1(_15671_),
    .C2(\icache.data_mems_0__data_mem.data_o [20]),
    .ZN(_18186_));
 AOI21_X2 _45011_ (.A(_17817_),
    .B1(_18184_),
    .B2(_18186_),
    .ZN(_18187_));
 NOR2_X4 _45012_ (.A1(_18183_),
    .A2(_18187_),
    .ZN(_18188_));
 OAI21_X1 _45013_ (.A(_18180_),
    .B1(_18188_),
    .B2(_18120_),
    .ZN(_05156_));
 NAND2_X1 _45014_ (.A1(_18179_),
    .A2(\icache.lce.lce_cmd_inst.data_r [341]),
    .ZN(_18189_));
 OR3_X2 _45015_ (.A1(_17089_),
    .A2(_17090_),
    .A3(_16226_),
    .ZN(_18190_));
 NAND2_X1 _45016_ (.A1(_17095_),
    .A2(_16347_),
    .ZN(_18191_));
 NAND2_X4 _45017_ (.A1(_18190_),
    .A2(_18191_),
    .ZN(_18192_));
 NAND2_X1 _45018_ (.A1(_18192_),
    .A2(_17960_),
    .ZN(_18193_));
 OAI21_X2 _45019_ (.A(_16386_),
    .B1(_17099_),
    .B2(_17100_),
    .ZN(_18194_));
 NAND3_X1 _45020_ (.A1(_17102_),
    .A2(_17104_),
    .A3(_16396_),
    .ZN(_18195_));
 NAND3_X1 _45021_ (.A1(_18194_),
    .A2(_16390_),
    .A3(_18195_),
    .ZN(_18196_));
 NAND2_X2 _45022_ (.A1(_18193_),
    .A2(_18196_),
    .ZN(_18197_));
 OAI21_X1 _45023_ (.A(_18189_),
    .B1(_18197_),
    .B2(_18120_),
    .ZN(_05157_));
 NAND2_X1 _45024_ (.A1(_18179_),
    .A2(\icache.lce.lce_cmd_inst.data_r [342]),
    .ZN(_18198_));
 OAI21_X1 _45025_ (.A(_16099_),
    .B1(_17112_),
    .B2(_17113_),
    .ZN(_18199_));
 OAI21_X2 _45026_ (.A(_15370_),
    .B1(_17109_),
    .B2(_17110_),
    .ZN(_18200_));
 AOI21_X2 _45027_ (.A(_16956_),
    .B1(_18199_),
    .B2(_18200_),
    .ZN(_18201_));
 OAI21_X2 _45028_ (.A(_15860_),
    .B1(_17121_),
    .B2(_17122_),
    .ZN(_18202_));
 OAI21_X2 _45029_ (.A(_15650_),
    .B1(_17117_),
    .B2(_17118_),
    .ZN(_18203_));
 AOI21_X2 _45030_ (.A(_17517_),
    .B1(_18202_),
    .B2(_18203_),
    .ZN(_18204_));
 NOR2_X4 _45031_ (.A1(_18201_),
    .A2(_18204_),
    .ZN(_18205_));
 BUF_X8 _45032_ (.A(_16785_),
    .Z(_18206_));
 OAI21_X1 _45033_ (.A(_18198_),
    .B1(_18205_),
    .B2(_18206_),
    .ZN(_05158_));
 NAND2_X1 _45034_ (.A1(_18179_),
    .A2(\icache.lce.lce_cmd_inst.data_r [343]),
    .ZN(_18207_));
 OR3_X4 _45035_ (.A1(_17127_),
    .A2(_17128_),
    .A3(_15394_),
    .ZN(_18208_));
 BUF_X16 _45036_ (.A(_15497_),
    .Z(_18209_));
 NAND2_X1 _45037_ (.A1(_17134_),
    .A2(_18209_),
    .ZN(_18210_));
 NAND2_X4 _45038_ (.A1(_18208_),
    .A2(_18210_),
    .ZN(_18211_));
 NAND2_X1 _45039_ (.A1(_18211_),
    .A2(_17960_),
    .ZN(_18212_));
 AOI21_X2 _45040_ (.A(_15576_),
    .B1(_17138_),
    .B2(_17140_),
    .ZN(_18213_));
 AOI21_X2 _45041_ (.A(_15740_),
    .B1(_17143_),
    .B2(_17145_),
    .ZN(_18214_));
 OAI21_X2 _45042_ (.A(_17500_),
    .B1(_18213_),
    .B2(_18214_),
    .ZN(_18215_));
 NAND2_X4 _45043_ (.A1(_18212_),
    .A2(_18215_),
    .ZN(_18216_));
 OAI21_X1 _45044_ (.A(_18207_),
    .B1(_18216_),
    .B2(_18206_),
    .ZN(_05159_));
 NAND2_X1 _45045_ (.A1(_18179_),
    .A2(\icache.lce.lce_cmd_inst.data_r [344]),
    .ZN(_18217_));
 AOI21_X2 _45046_ (.A(_15379_),
    .B1(_17162_),
    .B2(_17164_),
    .ZN(_18218_));
 AOI21_X2 _45047_ (.A(_18164_),
    .B1(_17166_),
    .B2(_17168_),
    .ZN(_18219_));
 OAI21_X2 _45048_ (.A(_17582_),
    .B1(_18218_),
    .B2(_18219_),
    .ZN(_18220_));
 NAND3_X2 _45049_ (.A1(_17152_),
    .A2(_17154_),
    .A3(_15754_),
    .ZN(_18221_));
 NAND3_X2 _45050_ (.A1(_17157_),
    .A2(_17159_),
    .A3(_15761_),
    .ZN(_18222_));
 NAND3_X2 _45051_ (.A1(_18221_),
    .A2(_18222_),
    .A3(_15996_),
    .ZN(_18223_));
 NAND2_X4 _45052_ (.A1(_18220_),
    .A2(_18223_),
    .ZN(_18224_));
 OAI21_X1 _45053_ (.A(_18217_),
    .B1(_18224_),
    .B2(_18206_),
    .ZN(_05160_));
 NAND2_X1 _45054_ (.A1(_18179_),
    .A2(\icache.lce.lce_cmd_inst.data_r [345]),
    .ZN(_18225_));
 NAND2_X1 _45055_ (.A1(_17176_),
    .A2(_17228_),
    .ZN(_18226_));
 NAND2_X1 _45056_ (.A1(_17182_),
    .A2(_18209_),
    .ZN(_18227_));
 NAND2_X2 _45057_ (.A1(_18226_),
    .A2(_18227_),
    .ZN(_18228_));
 NAND2_X1 _45058_ (.A1(_18228_),
    .A2(_17960_),
    .ZN(_18229_));
 OAI21_X2 _45059_ (.A(_16621_),
    .B1(_17187_),
    .B2(_17188_),
    .ZN(_18230_));
 NAND3_X2 _45060_ (.A1(_17190_),
    .A2(_17192_),
    .A3(_15901_),
    .ZN(_18231_));
 NAND3_X2 _45061_ (.A1(_18230_),
    .A2(_16390_),
    .A3(_18231_),
    .ZN(_18232_));
 NAND2_X4 _45062_ (.A1(_18229_),
    .A2(_18232_),
    .ZN(_18233_));
 OAI21_X1 _45063_ (.A(_18225_),
    .B1(_18233_),
    .B2(_18206_),
    .ZN(_05161_));
 NAND2_X1 _45064_ (.A1(_18179_),
    .A2(\icache.lce.lce_cmd_inst.data_r [346]),
    .ZN(_18234_));
 NAND2_X1 _45065_ (.A1(_17207_),
    .A2(_17228_),
    .ZN(_18235_));
 NAND2_X1 _45066_ (.A1(_17213_),
    .A2(_18209_),
    .ZN(_18236_));
 NAND2_X2 _45067_ (.A1(_18235_),
    .A2(_18236_),
    .ZN(_18237_));
 NAND2_X1 _45068_ (.A1(_18237_),
    .A2(_17731_),
    .ZN(_18238_));
 OAI21_X4 _45069_ (.A(_16386_),
    .B1(_17197_),
    .B2(_17198_),
    .ZN(_18239_));
 NAND2_X1 _45070_ (.A1(_15721_),
    .A2(_17201_),
    .ZN(_18240_));
 OAI211_X2 _45071_ (.A(_18240_),
    .B(_15567_),
    .C1(_15721_),
    .C2(\icache.data_mems_4__data_mem.data_o [26]),
    .ZN(_18241_));
 NAND3_X2 _45072_ (.A1(_18239_),
    .A2(_16823_),
    .A3(_18241_),
    .ZN(_18242_));
 NAND2_X4 _45073_ (.A1(_18238_),
    .A2(_18242_),
    .ZN(_18243_));
 OAI21_X1 _45074_ (.A(_18234_),
    .B1(_18243_),
    .B2(_18206_),
    .ZN(_05162_));
 NAND2_X1 _45075_ (.A1(_18179_),
    .A2(\icache.lce.lce_cmd_inst.data_r [347]),
    .ZN(_18244_));
 NOR3_X2 _45076_ (.A1(_17220_),
    .A2(_17221_),
    .A3(_15619_),
    .ZN(_18245_));
 AOI21_X2 _45077_ (.A(_18164_),
    .B1(_17223_),
    .B2(_17225_),
    .ZN(_18246_));
 OAI21_X2 _45078_ (.A(_17582_),
    .B1(_18245_),
    .B2(_18246_),
    .ZN(_18247_));
 OAI21_X2 _45079_ (.A(_16621_),
    .B1(_17230_),
    .B2(_17231_),
    .ZN(_18248_));
 NAND3_X2 _45080_ (.A1(_17233_),
    .A2(_17235_),
    .A3(_15901_),
    .ZN(_18249_));
 NAND3_X2 _45081_ (.A1(_18248_),
    .A2(_16390_),
    .A3(_18249_),
    .ZN(_18250_));
 NAND2_X4 _45082_ (.A1(_18247_),
    .A2(_18250_),
    .ZN(_18251_));
 OAI21_X1 _45083_ (.A(_18244_),
    .B1(_18251_),
    .B2(_18206_),
    .ZN(_05163_));
 NAND2_X1 _45084_ (.A1(_18179_),
    .A2(\icache.lce.lce_cmd_inst.data_r [348]),
    .ZN(_18252_));
 OAI21_X2 _45085_ (.A(_15708_),
    .B1(_17241_),
    .B2(_17242_),
    .ZN(_18253_));
 NAND3_X2 _45086_ (.A1(_17245_),
    .A2(_17247_),
    .A3(_15446_),
    .ZN(_18254_));
 AOI21_X2 _45087_ (.A(_16956_),
    .B1(_18253_),
    .B2(_18254_),
    .ZN(_18255_));
 OAI21_X2 _45088_ (.A(_17554_),
    .B1(_17255_),
    .B2(_17256_),
    .ZN(_18256_));
 OAI21_X1 _45089_ (.A(_15650_),
    .B1(_17251_),
    .B2(_17252_),
    .ZN(_18257_));
 AOI21_X2 _45090_ (.A(_17517_),
    .B1(_18256_),
    .B2(_18257_),
    .ZN(_18258_));
 NOR2_X4 _45091_ (.A1(_18255_),
    .A2(_18258_),
    .ZN(_18259_));
 OAI21_X1 _45092_ (.A(_18252_),
    .B1(_18259_),
    .B2(_18206_),
    .ZN(_05164_));
 NAND2_X1 _45093_ (.A1(_18179_),
    .A2(\icache.lce.lce_cmd_inst.data_r [349]),
    .ZN(_18260_));
 NOR2_X1 _45094_ (.A1(_17263_),
    .A2(_15545_),
    .ZN(_18261_));
 AOI21_X2 _45095_ (.A(_16056_),
    .B1(_17266_),
    .B2(_17267_),
    .ZN(_18262_));
 OAI21_X1 _45096_ (.A(_16631_),
    .B1(_18261_),
    .B2(_18262_),
    .ZN(_18263_));
 NAND2_X1 _45097_ (.A1(_17272_),
    .A2(_15343_),
    .ZN(_18264_));
 NAND2_X1 _45098_ (.A1(_17277_),
    .A2(_16230_),
    .ZN(_18265_));
 NAND3_X1 _45099_ (.A1(_18264_),
    .A2(_18265_),
    .A3(_15315_),
    .ZN(_18266_));
 AND2_X4 _45100_ (.A1(_18263_),
    .A2(_18266_),
    .ZN(_18267_));
 OAI21_X1 _45101_ (.A(_18260_),
    .B1(_18267_),
    .B2(_18206_),
    .ZN(_05165_));
 BUF_X16 _45102_ (.A(_15301_),
    .Z(_18268_));
 BUF_X8 _45103_ (.A(_18268_),
    .Z(_18269_));
 NAND2_X1 _45104_ (.A1(_18269_),
    .A2(\icache.lce.lce_cmd_inst.data_r [350]),
    .ZN(_18270_));
 NOR2_X4 _45105_ (.A1(_17284_),
    .A2(_16418_),
    .ZN(_18271_));
 AOI21_X4 _45106_ (.A(_15331_),
    .B1(_17286_),
    .B2(_17287_),
    .ZN(_18272_));
 OR3_X2 _45107_ (.A1(_18271_),
    .A2(_15597_),
    .A3(_18272_),
    .ZN(_18273_));
 OAI21_X2 _45108_ (.A(_16621_),
    .B1(_17294_),
    .B2(_17295_),
    .ZN(_18274_));
 OAI21_X2 _45109_ (.A(_15761_),
    .B1(_17291_),
    .B2(_17292_),
    .ZN(_18275_));
 NAND3_X2 _45110_ (.A1(_18274_),
    .A2(_18275_),
    .A3(_15656_),
    .ZN(_18276_));
 NAND2_X4 _45111_ (.A1(_18273_),
    .A2(_18276_),
    .ZN(_18277_));
 OAI21_X1 _45112_ (.A(_18270_),
    .B1(_18277_),
    .B2(_18206_),
    .ZN(_05167_));
 NAND2_X1 _45113_ (.A1(_18269_),
    .A2(\icache.lce.lce_cmd_inst.data_r [351]),
    .ZN(_18278_));
 OAI21_X2 _45114_ (.A(_16099_),
    .B1(_17309_),
    .B2(_17310_),
    .ZN(_18279_));
 NAND3_X2 _45115_ (.A1(_17313_),
    .A2(_17314_),
    .A3(_16578_),
    .ZN(_18280_));
 NAND3_X2 _45116_ (.A1(_18279_),
    .A2(_17567_),
    .A3(_18280_),
    .ZN(_18281_));
 OAI21_X2 _45117_ (.A(_15860_),
    .B1(_17301_),
    .B2(_17302_),
    .ZN(_18282_));
 NAND3_X2 _45118_ (.A1(_17304_),
    .A2(_17305_),
    .A3(_15994_),
    .ZN(_18283_));
 NAND3_X2 _45119_ (.A1(_18282_),
    .A2(_16823_),
    .A3(_18283_),
    .ZN(_18284_));
 NAND2_X4 _45120_ (.A1(_18281_),
    .A2(_18284_),
    .ZN(_18285_));
 OAI21_X1 _45121_ (.A(_18278_),
    .B1(_18285_),
    .B2(_18206_),
    .ZN(_05168_));
 NAND2_X1 _45122_ (.A1(_18269_),
    .A2(\icache.lce.lce_cmd_inst.data_r [352]),
    .ZN(_18286_));
 NOR2_X1 _45123_ (.A1(_17321_),
    .A2(_17264_),
    .ZN(_18287_));
 AOI21_X1 _45124_ (.A(_16643_),
    .B1(_17323_),
    .B2(_17324_),
    .ZN(_18288_));
 NOR3_X1 _45125_ (.A1(_18287_),
    .A2(_15724_),
    .A3(_18288_),
    .ZN(_18289_));
 NAND2_X1 _45126_ (.A1(_17333_),
    .A2(_16195_),
    .ZN(_18290_));
 NAND2_X1 _45127_ (.A1(_17329_),
    .A2(_16541_),
    .ZN(_18291_));
 AOI21_X1 _45128_ (.A(_15670_),
    .B1(_18290_),
    .B2(_18291_),
    .ZN(_18292_));
 OR2_X4 _45129_ (.A1(_18289_),
    .A2(_18292_),
    .ZN(_18293_));
 BUF_X16 _45130_ (.A(_15302_),
    .Z(_18294_));
 BUF_X16 _45131_ (.A(_18294_),
    .Z(_18295_));
 OAI21_X1 _45132_ (.A(_18286_),
    .B1(_18293_),
    .B2(_18295_),
    .ZN(_05169_));
 NAND2_X1 _45133_ (.A1(_18269_),
    .A2(\icache.lce.lce_cmd_inst.data_r [353]),
    .ZN(_18296_));
 OR3_X1 _45134_ (.A1(_17338_),
    .A2(_17339_),
    .A3(_15394_),
    .ZN(_18297_));
 NAND2_X1 _45135_ (.A1(_17343_),
    .A2(_18209_),
    .ZN(_18298_));
 NAND2_X2 _45136_ (.A1(_18297_),
    .A2(_18298_),
    .ZN(_18299_));
 NAND2_X1 _45137_ (.A1(_18299_),
    .A2(_17731_),
    .ZN(_18300_));
 OAI21_X2 _45138_ (.A(_16621_),
    .B1(_17346_),
    .B2(_17347_),
    .ZN(_18301_));
 NAND3_X2 _45139_ (.A1(_17349_),
    .A2(_17350_),
    .A3(_15901_),
    .ZN(_18302_));
 NAND3_X2 _45140_ (.A1(_18301_),
    .A2(_16823_),
    .A3(_18302_),
    .ZN(_18303_));
 NAND2_X4 _45141_ (.A1(_18300_),
    .A2(_18303_),
    .ZN(_18304_));
 OAI21_X1 _45142_ (.A(_18296_),
    .B1(_18304_),
    .B2(_18295_),
    .ZN(_05170_));
 NAND2_X1 _45143_ (.A1(_18269_),
    .A2(\icache.lce.lce_cmd_inst.data_r [354]),
    .ZN(_18305_));
 NOR2_X1 _45144_ (.A1(_15421_),
    .A2(\icache.data_mems_3__data_mem.data_o [34]),
    .ZN(_18306_));
 AOI211_X2 _45145_ (.A(_16229_),
    .B(_18306_),
    .C1(_16018_),
    .C2(_16042_),
    .ZN(_18307_));
 AOI21_X1 _45146_ (.A(_16307_),
    .B1(_17364_),
    .B2(_17365_),
    .ZN(_18308_));
 NOR3_X1 _45147_ (.A1(_18307_),
    .A2(_18308_),
    .A3(_16265_),
    .ZN(_18309_));
 NAND3_X1 _45148_ (.A1(_17358_),
    .A2(_17511_),
    .A3(_17359_),
    .ZN(_18310_));
 NAND2_X1 _45149_ (.A1(_16083_),
    .A2(\icache.data_mems_6__data_mem.data_o [34]),
    .ZN(_18311_));
 OAI211_X1 _45150_ (.A(_18311_),
    .B(_16307_),
    .C1(_15909_),
    .C2(_16036_),
    .ZN(_18312_));
 AOI21_X1 _45151_ (.A(_15579_),
    .B1(_18310_),
    .B2(_18312_),
    .ZN(_18313_));
 OR2_X4 _45152_ (.A1(_18309_),
    .A2(_18313_),
    .ZN(_18314_));
 OAI21_X1 _45153_ (.A(_18305_),
    .B1(_18314_),
    .B2(_18295_),
    .ZN(_05171_));
 NAND2_X1 _45154_ (.A1(_18269_),
    .A2(\icache.lce.lce_cmd_inst.data_r [355]),
    .ZN(_18315_));
 NAND2_X1 _45155_ (.A1(_17372_),
    .A2(_15770_),
    .ZN(_18316_));
 NAND2_X1 _45156_ (.A1(_17377_),
    .A2(_15514_),
    .ZN(_18317_));
 NAND3_X1 _45157_ (.A1(_18316_),
    .A2(_18317_),
    .A3(_15834_),
    .ZN(_18318_));
 AND3_X1 _45158_ (.A1(_17381_),
    .A2(_17382_),
    .A3(_16229_),
    .ZN(_18319_));
 AOI21_X2 _45159_ (.A(_15664_),
    .B1(_17384_),
    .B2(_17385_),
    .ZN(_18320_));
 OAI21_X1 _45160_ (.A(_17415_),
    .B1(_18319_),
    .B2(_18320_),
    .ZN(_18321_));
 AND2_X4 _45161_ (.A1(_18318_),
    .A2(_18321_),
    .ZN(_18322_));
 OAI21_X1 _45162_ (.A(_18315_),
    .B1(_18322_),
    .B2(_18295_),
    .ZN(_05172_));
 NAND2_X1 _45163_ (.A1(_18269_),
    .A2(\icache.lce.lce_cmd_inst.data_r [356]),
    .ZN(_18323_));
 BUF_X16 _45164_ (.A(_15597_),
    .Z(_18324_));
 NOR3_X2 _45165_ (.A1(_17396_),
    .A2(_17397_),
    .A3(_15619_),
    .ZN(_18325_));
 AOI21_X2 _45166_ (.A(_18164_),
    .B1(_17399_),
    .B2(_17400_),
    .ZN(_18326_));
 OAI21_X2 _45167_ (.A(_18324_),
    .B1(_18325_),
    .B2(_18326_),
    .ZN(_18327_));
 OAI21_X2 _45168_ (.A(_16621_),
    .B1(_17390_),
    .B2(_17391_),
    .ZN(_18328_));
 NAND2_X1 _45169_ (.A1(_16077_),
    .A2(_15479_),
    .ZN(_18329_));
 OAI211_X2 _45170_ (.A(_18329_),
    .B(_16578_),
    .C1(_18116_),
    .C2(\icache.data_mems_3__data_mem.data_o [36]),
    .ZN(_18330_));
 NAND3_X2 _45171_ (.A1(_18328_),
    .A2(_18330_),
    .A3(_15996_),
    .ZN(_18331_));
 NAND2_X4 _45172_ (.A1(_18327_),
    .A2(_18331_),
    .ZN(_18332_));
 OAI21_X1 _45173_ (.A(_18323_),
    .B1(_18332_),
    .B2(_18295_),
    .ZN(_05173_));
 NAND2_X1 _45174_ (.A1(_18269_),
    .A2(\icache.lce.lce_cmd_inst.data_r [357]),
    .ZN(_18333_));
 NAND2_X1 _45175_ (.A1(_17408_),
    .A2(_17228_),
    .ZN(_18334_));
 NAND2_X1 _45176_ (.A1(_17412_),
    .A2(_18209_),
    .ZN(_18335_));
 NAND2_X1 _45177_ (.A1(_18334_),
    .A2(_18335_),
    .ZN(_18336_));
 NAND2_X1 _45178_ (.A1(_18336_),
    .A2(_17731_),
    .ZN(_18337_));
 AND3_X1 _45179_ (.A1(_17419_),
    .A2(_16541_),
    .A3(_17420_),
    .ZN(_18338_));
 AOI21_X2 _45180_ (.A(_15740_),
    .B1(_17416_),
    .B2(_17417_),
    .ZN(_18339_));
 OAI21_X1 _45181_ (.A(_17971_),
    .B1(_18338_),
    .B2(_18339_),
    .ZN(_18340_));
 NAND2_X2 _45182_ (.A1(_18337_),
    .A2(_18340_),
    .ZN(_18341_));
 OAI21_X1 _45183_ (.A(_18333_),
    .B1(_18341_),
    .B2(_18295_),
    .ZN(_05174_));
 NAND2_X1 _45184_ (.A1(_18269_),
    .A2(\icache.lce.lce_cmd_inst.data_r [358]),
    .ZN(_18342_));
 NOR2_X1 _45185_ (.A1(_17427_),
    .A2(_15425_),
    .ZN(_18343_));
 AOI21_X1 _45186_ (.A(_16634_),
    .B1(_17429_),
    .B2(_17430_),
    .ZN(_18344_));
 OAI21_X1 _45187_ (.A(_16631_),
    .B1(_18343_),
    .B2(_18344_),
    .ZN(_18345_));
 NAND2_X1 _45188_ (.A1(_17435_),
    .A2(_17273_),
    .ZN(_18346_));
 NAND3_X1 _45189_ (.A1(_17437_),
    .A2(_15673_),
    .A3(_17438_),
    .ZN(_18347_));
 NAND3_X1 _45190_ (.A1(_18346_),
    .A2(_16372_),
    .A3(_18347_),
    .ZN(_18348_));
 AND2_X2 _45191_ (.A1(_18345_),
    .A2(_18348_),
    .ZN(_18349_));
 OAI21_X1 _45192_ (.A(_18342_),
    .B1(_18349_),
    .B2(_18295_),
    .ZN(_05175_));
 NAND2_X1 _45193_ (.A1(_18269_),
    .A2(\icache.lce.lce_cmd_inst.data_r [359]),
    .ZN(_18350_));
 BUF_X16 _45194_ (.A(_15314_),
    .Z(_18351_));
 NAND2_X1 _45195_ (.A1(_17451_),
    .A2(_15395_),
    .ZN(_18352_));
 NAND3_X2 _45196_ (.A1(_17453_),
    .A2(_16418_),
    .A3(_17454_),
    .ZN(_18353_));
 AOI21_X1 _45197_ (.A(_18351_),
    .B1(_18352_),
    .B2(_18353_),
    .ZN(_18354_));
 NAND3_X2 _45198_ (.A1(_17445_),
    .A2(_17459_),
    .A3(_17446_),
    .ZN(_18355_));
 NAND2_X1 _45199_ (.A1(_16083_),
    .A2(\icache.data_mems_0__data_mem.data_o [39]),
    .ZN(_18356_));
 OAI211_X4 _45200_ (.A(_18356_),
    .B(_15678_),
    .C1(_15909_),
    .C2(_16149_),
    .ZN(_18357_));
 AOI21_X1 _45201_ (.A(_15670_),
    .B1(_18355_),
    .B2(_18357_),
    .ZN(_18358_));
 OR2_X2 _45202_ (.A1(_18354_),
    .A2(_18358_),
    .ZN(_18359_));
 OAI21_X1 _45203_ (.A(_18350_),
    .B1(_18359_),
    .B2(_18295_),
    .ZN(_05176_));
 BUF_X4 _45204_ (.A(_18268_),
    .Z(_18360_));
 NAND2_X1 _45205_ (.A1(_18360_),
    .A2(\icache.lce.lce_cmd_inst.data_r [360]),
    .ZN(_18361_));
 NOR2_X1 _45206_ (.A1(_15537_),
    .A2(\icache.data_mems_0__data_mem.data_o [40]),
    .ZN(_18362_));
 AOI211_X2 _45207_ (.A(_15445_),
    .B(_18362_),
    .C1(_16035_),
    .C2(_16168_),
    .ZN(_18363_));
 AOI21_X1 _45208_ (.A(_15477_),
    .B1(_17467_),
    .B2(_17468_),
    .ZN(_18364_));
 OAI21_X1 _45209_ (.A(_16438_),
    .B1(_18363_),
    .B2(_18364_),
    .ZN(_18365_));
 BUF_X8 _45210_ (.A(_15408_),
    .Z(_18366_));
 AOI21_X1 _45211_ (.A(_17459_),
    .B1(_17463_),
    .B2(_17464_),
    .ZN(_18367_));
 AOI21_X1 _45212_ (.A(_16324_),
    .B1(_17460_),
    .B2(_17461_),
    .ZN(_18368_));
 OAI21_X1 _45213_ (.A(_18366_),
    .B1(_18367_),
    .B2(_18368_),
    .ZN(_18369_));
 AND2_X4 _45214_ (.A1(_18365_),
    .A2(_18369_),
    .ZN(_18370_));
 OAI21_X1 _45215_ (.A(_18361_),
    .B1(_18370_),
    .B2(_18295_),
    .ZN(_05178_));
 NAND2_X1 _45216_ (.A1(_18360_),
    .A2(\icache.lce.lce_cmd_inst.data_r [361]),
    .ZN(_18371_));
 NOR2_X1 _45217_ (.A1(_15751_),
    .A2(\icache.data_mems_7__data_mem.data_o [41]),
    .ZN(_18372_));
 AOI211_X2 _45218_ (.A(_15544_),
    .B(_18372_),
    .C1(_16112_),
    .C2(_16179_),
    .ZN(_18373_));
 AOI21_X2 _45219_ (.A(_15369_),
    .B1(_17482_),
    .B2(_17483_),
    .ZN(_18374_));
 OR3_X2 _45220_ (.A1(_18373_),
    .A2(_18374_),
    .A3(_15699_),
    .ZN(_18375_));
 BUF_X32 _45221_ (.A(_15644_),
    .Z(_18376_));
 NOR3_X2 _45222_ (.A1(_17475_),
    .A2(_17476_),
    .A3(_15311_),
    .ZN(_18377_));
 AOI21_X4 _45223_ (.A(_16053_),
    .B1(_17478_),
    .B2(_17479_),
    .ZN(_18378_));
 OAI21_X2 _45224_ (.A(_18376_),
    .B1(_18377_),
    .B2(_18378_),
    .ZN(_18379_));
 NAND2_X4 _45225_ (.A1(_18375_),
    .A2(_18379_),
    .ZN(_18380_));
 OAI21_X1 _45226_ (.A(_18371_),
    .B1(_18380_),
    .B2(_18295_),
    .ZN(_05179_));
 NAND2_X1 _45227_ (.A1(_18360_),
    .A2(\icache.lce.lce_cmd_inst.data_r [362]),
    .ZN(_18381_));
 AOI21_X1 _45228_ (.A(_15727_),
    .B1(_17513_),
    .B2(_17514_),
    .ZN(_18382_));
 NAND2_X1 _45229_ (.A1(_15573_),
    .A2(\icache.data_mems_2__data_mem.data_o [42]),
    .ZN(_18383_));
 AOI21_X1 _45230_ (.A(_16643_),
    .B1(_17510_),
    .B2(_18383_),
    .ZN(_18384_));
 OR3_X1 _45231_ (.A1(_18382_),
    .A2(_18384_),
    .A3(_15655_),
    .ZN(_18385_));
 NOR3_X2 _45232_ (.A1(_17518_),
    .A2(_17519_),
    .A3(_17981_),
    .ZN(_18386_));
 AOI21_X2 _45233_ (.A(_15740_),
    .B1(_17521_),
    .B2(_17522_),
    .ZN(_18387_));
 OAI21_X2 _45234_ (.A(_17971_),
    .B1(_18386_),
    .B2(_18387_),
    .ZN(_18388_));
 NAND2_X4 _45235_ (.A1(_18385_),
    .A2(_18388_),
    .ZN(_18389_));
 BUF_X4 _45236_ (.A(_18294_),
    .Z(_18390_));
 OAI21_X1 _45237_ (.A(_18381_),
    .B1(_18389_),
    .B2(_18390_),
    .ZN(_05180_));
 NAND2_X1 _45238_ (.A1(_18360_),
    .A2(\icache.lce.lce_cmd_inst.data_r [363]),
    .ZN(_18391_));
 NAND2_X1 _45239_ (.A1(_17534_),
    .A2(_16578_),
    .ZN(_18392_));
 NAND2_X1 _45240_ (.A1(_17530_),
    .A2(_15594_),
    .ZN(_18393_));
 NAND3_X1 _45241_ (.A1(_18392_),
    .A2(_18393_),
    .A3(_15834_),
    .ZN(_18394_));
 AND3_X1 _45242_ (.A1(_17541_),
    .A2(_17542_),
    .A3(_16643_),
    .ZN(_18395_));
 AOI21_X1 _45243_ (.A(_16324_),
    .B1(_17538_),
    .B2(_17539_),
    .ZN(_18396_));
 OAI21_X1 _45244_ (.A(_18366_),
    .B1(_18395_),
    .B2(_18396_),
    .ZN(_18397_));
 AND2_X4 _45245_ (.A1(_18394_),
    .A2(_18397_),
    .ZN(_18398_));
 OAI21_X1 _45246_ (.A(_18391_),
    .B1(_18398_),
    .B2(_18390_),
    .ZN(_05181_));
 NAND2_X1 _45247_ (.A1(_18360_),
    .A2(\icache.lce.lce_cmd_inst.data_r [364]),
    .ZN(_18399_));
 OR3_X1 _45248_ (.A1(_17547_),
    .A2(_17548_),
    .A3(_16321_),
    .ZN(_18400_));
 OR3_X1 _45249_ (.A1(_17550_),
    .A2(_17551_),
    .A3(_17068_),
    .ZN(_18401_));
 AOI21_X1 _45250_ (.A(_18351_),
    .B1(_18400_),
    .B2(_18401_),
    .ZN(_18402_));
 OAI21_X2 _45251_ (.A(_16327_),
    .B1(_17558_),
    .B2(_17559_),
    .ZN(_18403_));
 OAI21_X1 _45252_ (.A(_15445_),
    .B1(_17555_),
    .B2(_17556_),
    .ZN(_18404_));
 AND3_X1 _45253_ (.A1(_18403_),
    .A2(_18404_),
    .A3(_15328_),
    .ZN(_18405_));
 OR2_X2 _45254_ (.A1(_18402_),
    .A2(_18405_),
    .ZN(_18406_));
 OAI21_X1 _45255_ (.A(_18399_),
    .B1(_18406_),
    .B2(_18390_),
    .ZN(_05182_));
 NAND2_X1 _45256_ (.A1(_18360_),
    .A2(\icache.lce.lce_cmd_inst.data_r [365]),
    .ZN(_18407_));
 OR3_X1 _45257_ (.A1(_15506_),
    .A2(_15507_),
    .A3(_16053_),
    .ZN(_18408_));
 NAND2_X1 _45258_ (.A1(_15513_),
    .A2(_15932_),
    .ZN(_18409_));
 AND3_X1 _45259_ (.A1(_18408_),
    .A2(_15474_),
    .A3(_18409_),
    .ZN(_18410_));
 OAI21_X1 _45260_ (.A(_17554_),
    .B1(_15519_),
    .B2(_15520_),
    .ZN(_18411_));
 NAND3_X2 _45261_ (.A1(_15525_),
    .A2(_15527_),
    .A3(_16217_),
    .ZN(_18412_));
 AOI21_X1 _45262_ (.A(_17517_),
    .B1(_18411_),
    .B2(_18412_),
    .ZN(_18413_));
 NOR2_X2 _45263_ (.A1(_18410_),
    .A2(_18413_),
    .ZN(_18414_));
 OAI21_X1 _45264_ (.A(_18407_),
    .B1(_18414_),
    .B2(_18390_),
    .ZN(_05183_));
 NAND2_X1 _45265_ (.A1(_18360_),
    .A2(\icache.lce.lce_cmd_inst.data_r [366]),
    .ZN(_18415_));
 OAI21_X2 _45266_ (.A(_15432_),
    .B1(_15555_),
    .B2(_15557_),
    .ZN(_18416_));
 OAI21_X2 _45267_ (.A(_16634_),
    .B1(_15549_),
    .B2(_15551_),
    .ZN(_18417_));
 AND3_X1 _45268_ (.A1(_18416_),
    .A2(_18417_),
    .A3(_15522_),
    .ZN(_18418_));
 BUF_X16 _45269_ (.A(_15502_),
    .Z(_18419_));
 OR3_X1 _45270_ (.A1(_15534_),
    .A2(_15535_),
    .A3(_17068_),
    .ZN(_18420_));
 NAND2_X1 _45271_ (.A1(_15543_),
    .A2(_17988_),
    .ZN(_18421_));
 AOI21_X1 _45272_ (.A(_18419_),
    .B1(_18420_),
    .B2(_18421_),
    .ZN(_18422_));
 OR2_X2 _45273_ (.A1(_18418_),
    .A2(_18422_),
    .ZN(_18423_));
 OAI21_X1 _45274_ (.A(_18415_),
    .B1(_18423_),
    .B2(_18390_),
    .ZN(_05184_));
 NAND2_X1 _45275_ (.A1(_18360_),
    .A2(\icache.lce.lce_cmd_inst.data_r [367]),
    .ZN(_18424_));
 NAND2_X1 _45276_ (.A1(_15566_),
    .A2(_15587_),
    .ZN(_18425_));
 NAND2_X1 _45277_ (.A1(_15575_),
    .A2(_15594_),
    .ZN(_18426_));
 NAND2_X1 _45278_ (.A1(_18425_),
    .A2(_18426_),
    .ZN(_18427_));
 NAND2_X1 _45279_ (.A1(_18427_),
    .A2(_17731_),
    .ZN(_18428_));
 NAND2_X1 _45280_ (.A1(_15585_),
    .A2(_15567_),
    .ZN(_18429_));
 NAND2_X1 _45281_ (.A1(_15593_),
    .A2(_15576_),
    .ZN(_18430_));
 NAND2_X1 _45282_ (.A1(_18429_),
    .A2(_18430_),
    .ZN(_18431_));
 NAND2_X1 _45283_ (.A1(_18431_),
    .A2(_15598_),
    .ZN(_18432_));
 NAND2_X2 _45284_ (.A1(_18428_),
    .A2(_18432_),
    .ZN(_18433_));
 OAI21_X1 _45285_ (.A(_18424_),
    .B1(_18433_),
    .B2(_18390_),
    .ZN(_05185_));
 NAND2_X1 _45286_ (.A1(_18360_),
    .A2(\icache.lce.lce_cmd_inst.data_r [368]),
    .ZN(_18434_));
 NAND2_X1 _45287_ (.A1(_15608_),
    .A2(_16341_),
    .ZN(_18435_));
 NAND2_X1 _45288_ (.A1(_15618_),
    .A2(_15587_),
    .ZN(_18436_));
 NAND2_X2 _45289_ (.A1(_18435_),
    .A2(_18436_),
    .ZN(_18437_));
 NAND2_X1 _45290_ (.A1(_18437_),
    .A2(_17731_),
    .ZN(_18438_));
 OAI21_X2 _45291_ (.A(_16386_),
    .B1(_15624_),
    .B2(_15625_),
    .ZN(_18439_));
 NAND3_X4 _45292_ (.A1(_15629_),
    .A2(_15631_),
    .A3(_16396_),
    .ZN(_18440_));
 NAND3_X4 _45293_ (.A1(_18439_),
    .A2(_16823_),
    .A3(_18440_),
    .ZN(_18441_));
 NAND2_X2 _45294_ (.A1(_18438_),
    .A2(_18441_),
    .ZN(_18442_));
 OAI21_X1 _45295_ (.A(_18434_),
    .B1(_18442_),
    .B2(_18390_),
    .ZN(_05186_));
 NAND2_X1 _45296_ (.A1(_18360_),
    .A2(\icache.lce.lce_cmd_inst.data_r [369]),
    .ZN(_18443_));
 OAI21_X2 _45297_ (.A(_15712_),
    .B1(_15637_),
    .B2(_15638_),
    .ZN(_18444_));
 OAI21_X2 _45298_ (.A(_15332_),
    .B1(_15641_),
    .B2(_15642_),
    .ZN(_18445_));
 NAND3_X2 _45299_ (.A1(_18444_),
    .A2(_17567_),
    .A3(_18445_),
    .ZN(_18446_));
 OAI21_X2 _45300_ (.A(_17308_),
    .B1(_15647_),
    .B2(_15648_),
    .ZN(_18447_));
 OAI21_X2 _45301_ (.A(_15594_),
    .B1(_15652_),
    .B2(_15653_),
    .ZN(_18448_));
 NAND3_X2 _45302_ (.A1(_18447_),
    .A2(_16823_),
    .A3(_18448_),
    .ZN(_18449_));
 NAND2_X4 _45303_ (.A1(_18446_),
    .A2(_18449_),
    .ZN(_18450_));
 OAI21_X1 _45304_ (.A(_18443_),
    .B1(_18450_),
    .B2(_18390_),
    .ZN(_05187_));
 BUF_X4 _45305_ (.A(_18268_),
    .Z(_18451_));
 NAND2_X1 _45306_ (.A1(_18451_),
    .A2(\icache.lce.lce_cmd_inst.data_r [370]),
    .ZN(_18452_));
 OAI21_X2 _45307_ (.A(_16099_),
    .B1(_15661_),
    .B2(_15662_),
    .ZN(_18453_));
 OAI21_X2 _45308_ (.A(_15370_),
    .B1(_15666_),
    .B2(_15667_),
    .ZN(_18454_));
 NAND3_X2 _45309_ (.A1(_18453_),
    .A2(_18454_),
    .A3(_16143_),
    .ZN(_18455_));
 NAND2_X1 _45310_ (.A1(_15675_),
    .A2(_15909_),
    .ZN(_18456_));
 OAI211_X2 _45311_ (.A(_18456_),
    .B(_15395_),
    .C1(_18116_),
    .C2(\icache.data_mems_1__data_mem.data_o [50]),
    .ZN(_18457_));
 NAND2_X1 _45312_ (.A1(_15680_),
    .A2(_17839_),
    .ZN(_18458_));
 OAI211_X4 _45313_ (.A(_18458_),
    .B(_17981_),
    .C1(_15324_),
    .C2(\icache.data_mems_3__data_mem.data_o [50]),
    .ZN(_18459_));
 BUF_X16 _45314_ (.A(_15644_),
    .Z(_18460_));
 NAND3_X2 _45315_ (.A1(_18457_),
    .A2(_18459_),
    .A3(_18460_),
    .ZN(_18461_));
 NAND2_X4 _45316_ (.A1(_18455_),
    .A2(_18461_),
    .ZN(_18462_));
 OAI21_X1 _45317_ (.A(_18452_),
    .B1(_18462_),
    .B2(_18390_),
    .ZN(_05189_));
 NAND2_X1 _45318_ (.A1(_18451_),
    .A2(\icache.lce.lce_cmd_inst.data_r [371]),
    .ZN(_18463_));
 OAI21_X1 _45319_ (.A(_15712_),
    .B1(_15696_),
    .B2(_15697_),
    .ZN(_18464_));
 NAND3_X4 _45320_ (.A1(_15701_),
    .A2(_15703_),
    .A3(_15911_),
    .ZN(_18465_));
 NAND3_X1 _45321_ (.A1(_18464_),
    .A2(_17567_),
    .A3(_18465_),
    .ZN(_18466_));
 OR2_X1 _45322_ (.A1(_15375_),
    .A2(\icache.data_mems_7__data_mem.data_o [51]),
    .ZN(_18467_));
 OAI211_X4 _45323_ (.A(_18467_),
    .B(_18164_),
    .C1(_15721_),
    .C2(\icache.data_mems_6__data_mem.data_o [51]),
    .ZN(_18468_));
 OAI21_X2 _45324_ (.A(_15594_),
    .B1(_15688_),
    .B2(_15689_),
    .ZN(_18469_));
 BUF_X16 _45325_ (.A(_15655_),
    .Z(_18470_));
 NAND3_X2 _45326_ (.A1(_18468_),
    .A2(_18469_),
    .A3(_18470_),
    .ZN(_18471_));
 NAND2_X4 _45327_ (.A1(_18466_),
    .A2(_18471_),
    .ZN(_18472_));
 OAI21_X1 _45328_ (.A(_18463_),
    .B1(_18472_),
    .B2(_18390_),
    .ZN(_05190_));
 NAND2_X1 _45329_ (.A1(_18451_),
    .A2(\icache.lce.lce_cmd_inst.data_r [372]),
    .ZN(_18473_));
 OR3_X1 _45330_ (.A1(_15709_),
    .A2(_15710_),
    .A3(_16321_),
    .ZN(_18474_));
 OR3_X1 _45331_ (.A1(_15715_),
    .A2(_15716_),
    .A3(_17068_),
    .ZN(_18475_));
 AND3_X1 _45332_ (.A1(_18474_),
    .A2(_18475_),
    .A3(_15940_),
    .ZN(_18476_));
 NAND2_X1 _45333_ (.A1(_16427_),
    .A2(_15478_),
    .ZN(_18477_));
 OAI211_X4 _45334_ (.A(_18477_),
    .B(_16229_),
    .C1(_16394_),
    .C2(\icache.data_mems_1__data_mem.data_o [52]),
    .ZN(_18478_));
 NAND2_X1 _45335_ (.A1(_15722_),
    .A2(_15495_),
    .ZN(_18479_));
 OAI211_X2 _45336_ (.A(_18479_),
    .B(_15609_),
    .C1(_15725_),
    .C2(\icache.data_mems_3__data_mem.data_o [52]),
    .ZN(_18480_));
 AOI21_X2 _45337_ (.A(_17817_),
    .B1(_18478_),
    .B2(_18480_),
    .ZN(_18481_));
 NOR2_X4 _45338_ (.A1(_18476_),
    .A2(_18481_),
    .ZN(_18482_));
 BUF_X8 _45339_ (.A(_18294_),
    .Z(_18483_));
 OAI21_X1 _45340_ (.A(_18473_),
    .B1(_18482_),
    .B2(_18483_),
    .ZN(_05191_));
 NAND2_X1 _45341_ (.A1(_18451_),
    .A2(\icache.lce.lce_cmd_inst.data_r [373]),
    .ZN(_18484_));
 AOI21_X4 _45342_ (.A(_17710_),
    .B1(_15749_),
    .B2(_15753_),
    .ZN(_18485_));
 AOI21_X2 _45343_ (.A(_17988_),
    .B1(_15758_),
    .B2(_15760_),
    .ZN(_18486_));
 NOR3_X2 _45344_ (.A1(_18485_),
    .A2(_18486_),
    .A3(_18132_),
    .ZN(_18487_));
 OAI21_X2 _45345_ (.A(_15860_),
    .B1(_15737_),
    .B2(_15739_),
    .ZN(_18488_));
 NAND3_X2 _45346_ (.A1(_15742_),
    .A2(_15744_),
    .A3(_15994_),
    .ZN(_18489_));
 AOI21_X2 _45347_ (.A(_17817_),
    .B1(_18488_),
    .B2(_18489_),
    .ZN(_18490_));
 NOR2_X4 _45348_ (.A1(_18487_),
    .A2(_18490_),
    .ZN(_18491_));
 OAI21_X1 _45349_ (.A(_18484_),
    .B1(_18491_),
    .B2(_18483_),
    .ZN(_05192_));
 NAND2_X1 _45350_ (.A1(_18451_),
    .A2(\icache.lce.lce_cmd_inst.data_r [374]),
    .ZN(_18492_));
 NAND2_X1 _45351_ (.A1(_15769_),
    .A2(_15395_),
    .ZN(_18493_));
 NAND2_X1 _45352_ (.A1(_15778_),
    .A2(_17981_),
    .ZN(_18494_));
 AOI21_X1 _45353_ (.A(_18351_),
    .B1(_18493_),
    .B2(_18494_),
    .ZN(_18495_));
 OAI21_X1 _45354_ (.A(_15812_),
    .B1(_15788_),
    .B2(_15789_),
    .ZN(_18496_));
 OAI21_X1 _45355_ (.A(_15445_),
    .B1(_15783_),
    .B2(_15785_),
    .ZN(_18497_));
 AND3_X1 _45356_ (.A1(_18496_),
    .A2(_18497_),
    .A3(_15328_),
    .ZN(_18498_));
 OR2_X2 _45357_ (.A1(_18495_),
    .A2(_18498_),
    .ZN(_18499_));
 OAI21_X1 _45358_ (.A(_18492_),
    .B1(_18499_),
    .B2(_18483_),
    .ZN(_05193_));
 NAND2_X1 _45359_ (.A1(_18451_),
    .A2(\icache.lce.lce_cmd_inst.data_r [375]),
    .ZN(_18500_));
 NAND2_X1 _45360_ (.A1(_15797_),
    .A2(_16341_),
    .ZN(_18501_));
 NAND2_X1 _45361_ (.A1(_15803_),
    .A2(_15587_),
    .ZN(_18502_));
 NAND2_X1 _45362_ (.A1(_18501_),
    .A2(_18502_),
    .ZN(_18503_));
 NAND2_X1 _45363_ (.A1(_18503_),
    .A2(_17731_),
    .ZN(_18504_));
 AOI21_X2 _45364_ (.A(_16014_),
    .B1(_15808_),
    .B2(_15811_),
    .ZN(_18505_));
 AOI21_X2 _45365_ (.A(_16227_),
    .B1(_15815_),
    .B2(_15817_),
    .ZN(_18506_));
 OAI21_X2 _45366_ (.A(_17971_),
    .B1(_18505_),
    .B2(_18506_),
    .ZN(_18507_));
 NAND2_X2 _45367_ (.A1(_18504_),
    .A2(_18507_),
    .ZN(_18508_));
 OAI21_X1 _45368_ (.A(_18500_),
    .B1(_18508_),
    .B2(_18483_),
    .ZN(_05194_));
 NAND2_X1 _45369_ (.A1(_18451_),
    .A2(\icache.lce.lce_cmd_inst.data_r [376]),
    .ZN(_18509_));
 NAND2_X1 _45370_ (.A1(_15831_),
    .A2(_17228_),
    .ZN(_18510_));
 NAND2_X1 _45371_ (.A1(_15826_),
    .A2(_18209_),
    .ZN(_18511_));
 NAND2_X1 _45372_ (.A1(_18510_),
    .A2(_18511_),
    .ZN(_18512_));
 NAND2_X1 _45373_ (.A1(_18512_),
    .A2(_17731_),
    .ZN(_18513_));
 NAND2_X1 _45374_ (.A1(_15847_),
    .A2(_15587_),
    .ZN(_18514_));
 NAND2_X1 _45375_ (.A1(_15841_),
    .A2(_15594_),
    .ZN(_18515_));
 NAND2_X1 _45376_ (.A1(_18514_),
    .A2(_18515_),
    .ZN(_18516_));
 NAND2_X1 _45377_ (.A1(_18516_),
    .A2(_15598_),
    .ZN(_18517_));
 NAND2_X2 _45378_ (.A1(_18513_),
    .A2(_18517_),
    .ZN(_18518_));
 OAI21_X1 _45379_ (.A(_18509_),
    .B1(_18518_),
    .B2(_18483_),
    .ZN(_05195_));
 NAND2_X1 _45380_ (.A1(_18451_),
    .A2(\icache.lce.lce_cmd_inst.data_r [377]),
    .ZN(_18519_));
 NOR3_X2 _45381_ (.A1(_15854_),
    .A2(_15855_),
    .A3(_16195_),
    .ZN(_18520_));
 AOI21_X2 _45382_ (.A(_15938_),
    .B1(_15857_),
    .B2(_15859_),
    .ZN(_18521_));
 OAI21_X2 _45383_ (.A(_18324_),
    .B1(_18520_),
    .B2(_18521_),
    .ZN(_18522_));
 OAI21_X2 _45384_ (.A(_15860_),
    .B1(_15868_),
    .B2(_15869_),
    .ZN(_18523_));
 OAI21_X2 _45385_ (.A(_15650_),
    .B1(_15864_),
    .B2(_15865_),
    .ZN(_18524_));
 NAND3_X2 _45386_ (.A1(_18523_),
    .A2(_18524_),
    .A3(_18460_),
    .ZN(_18525_));
 NAND2_X4 _45387_ (.A1(_18522_),
    .A2(_18525_),
    .ZN(_18526_));
 OAI21_X1 _45388_ (.A(_18519_),
    .B1(_18526_),
    .B2(_18483_),
    .ZN(_05196_));
 NAND2_X1 _45389_ (.A1(_18451_),
    .A2(\icache.lce.lce_cmd_inst.data_r [378]),
    .ZN(_18527_));
 NAND2_X1 _45390_ (.A1(_15895_),
    .A2(_15610_),
    .ZN(_18528_));
 NAND2_X1 _45391_ (.A1(_15889_),
    .A2(_15619_),
    .ZN(_18529_));
 AND3_X1 _45392_ (.A1(_18528_),
    .A2(_18529_),
    .A3(_15940_),
    .ZN(_18530_));
 BUF_X16 _45393_ (.A(_15367_),
    .Z(_18531_));
 OAI21_X4 _45394_ (.A(_16865_),
    .B1(_15875_),
    .B2(_15877_),
    .ZN(_18532_));
 OAI21_X4 _45395_ (.A(_15379_),
    .B1(_15880_),
    .B2(_15881_),
    .ZN(_18533_));
 AOI21_X4 _45396_ (.A(_18531_),
    .B1(_18532_),
    .B2(_18533_),
    .ZN(_18534_));
 NOR2_X4 _45397_ (.A1(_18530_),
    .A2(_18534_),
    .ZN(_18535_));
 OAI21_X1 _45398_ (.A(_18527_),
    .B1(_18535_),
    .B2(_18483_),
    .ZN(_05197_));
 NAND2_X1 _45399_ (.A1(_18451_),
    .A2(\icache.lce.lce_cmd_inst.data_r [379]),
    .ZN(_18536_));
 NAND2_X1 _45400_ (.A1(_17496_),
    .A2(_16021_),
    .ZN(_18537_));
 NAND2_X1 _45401_ (.A1(_17492_),
    .A2(_15804_),
    .ZN(_18538_));
 AOI21_X1 _45402_ (.A(_18351_),
    .B1(_18537_),
    .B2(_18538_),
    .ZN(_18539_));
 OAI21_X2 _45403_ (.A(_15812_),
    .B1(_17501_),
    .B2(_17502_),
    .ZN(_18540_));
 NAND3_X1 _45404_ (.A1(_17504_),
    .A2(_17505_),
    .A3(_15342_),
    .ZN(_18541_));
 AND3_X1 _45405_ (.A1(_18540_),
    .A2(_15430_),
    .A3(_18541_),
    .ZN(_18542_));
 OR2_X4 _45406_ (.A1(_18539_),
    .A2(_18542_),
    .ZN(_18543_));
 OAI21_X1 _45407_ (.A(_18536_),
    .B1(_18543_),
    .B2(_18483_),
    .ZN(_05198_));
 BUF_X8 _45408_ (.A(_18268_),
    .Z(_18544_));
 NAND2_X1 _45409_ (.A1(_18544_),
    .A2(\icache.lce.lce_cmd_inst.data_r [380]),
    .ZN(_18545_));
 OAI21_X1 _45410_ (.A(_15708_),
    .B1(_15470_),
    .B2(_15472_),
    .ZN(_18546_));
 NAND2_X1 _45411_ (.A1(_16589_),
    .A2(_15986_),
    .ZN(_18547_));
 OAI211_X2 _45412_ (.A(_18547_),
    .B(_15610_),
    .C1(_18116_),
    .C2(\icache.data_mems_3__data_mem.data_o [60]),
    .ZN(_18548_));
 AOI21_X2 _45413_ (.A(_16956_),
    .B1(_18546_),
    .B2(_18548_),
    .ZN(_18549_));
 OAI21_X2 _45414_ (.A(_17554_),
    .B1(_15487_),
    .B2(_15489_),
    .ZN(_18550_));
 NAND3_X1 _45415_ (.A1(_15493_),
    .A2(_15496_),
    .A3(_15464_),
    .ZN(_18551_));
 AOI21_X2 _45416_ (.A(_17517_),
    .B1(_18550_),
    .B2(_18551_),
    .ZN(_18552_));
 NOR2_X4 _45417_ (.A1(_18549_),
    .A2(_18552_),
    .ZN(_18553_));
 OAI21_X1 _45418_ (.A(_18545_),
    .B1(_18553_),
    .B2(_18483_),
    .ZN(_05200_));
 NAND2_X1 _45419_ (.A1(_18544_),
    .A2(\icache.lce.lce_cmd_inst.data_r [381]),
    .ZN(_18554_));
 NOR3_X2 _45420_ (.A1(_15437_),
    .A2(_15439_),
    .A3(_17273_),
    .ZN(_18555_));
 AOI21_X2 _45421_ (.A(_17988_),
    .B1(_15441_),
    .B2(_15444_),
    .ZN(_18556_));
 NOR3_X2 _45422_ (.A1(_18555_),
    .A2(_18556_),
    .A3(_18132_),
    .ZN(_18557_));
 OAI21_X2 _45423_ (.A(_17308_),
    .B1(_15453_),
    .B2(_15455_),
    .ZN(_18558_));
 NAND3_X2 _45424_ (.A1(_15458_),
    .A2(_15462_),
    .A3(_17236_),
    .ZN(_18559_));
 AOI21_X2 _45425_ (.A(_18531_),
    .B1(_18558_),
    .B2(_18559_),
    .ZN(_18560_));
 NOR2_X4 _45426_ (.A1(_18557_),
    .A2(_18560_),
    .ZN(_18561_));
 OAI21_X1 _45427_ (.A(_18554_),
    .B1(_18561_),
    .B2(_18483_),
    .ZN(_05201_));
 NAND2_X1 _45428_ (.A1(_18544_),
    .A2(\icache.lce.lce_cmd_inst.data_r [382]),
    .ZN(_18562_));
 NAND2_X1 _45429_ (.A1(_15415_),
    .A2(_15567_),
    .ZN(_18563_));
 NAND2_X1 _45430_ (.A1(_15423_),
    .A2(_15576_),
    .ZN(_18564_));
 NAND2_X1 _45431_ (.A1(_18563_),
    .A2(_18564_),
    .ZN(_18565_));
 NAND2_X1 _45432_ (.A1(_18565_),
    .A2(_17731_),
    .ZN(_18566_));
 NAND2_X1 _45433_ (.A1(_15393_),
    .A2(_15587_),
    .ZN(_18567_));
 NAND2_X1 _45434_ (.A1(_15404_),
    .A2(_15594_),
    .ZN(_18568_));
 NAND2_X1 _45435_ (.A1(_18567_),
    .A2(_18568_),
    .ZN(_18569_));
 NAND2_X1 _45436_ (.A1(_18569_),
    .A2(_15598_),
    .ZN(_18570_));
 NAND2_X2 _45437_ (.A1(_18566_),
    .A2(_18570_),
    .ZN(_18571_));
 BUF_X16 _45438_ (.A(_18294_),
    .Z(_18572_));
 OAI21_X1 _45439_ (.A(_18562_),
    .B1(_18571_),
    .B2(_18572_),
    .ZN(_05202_));
 NAND2_X1 _45440_ (.A1(_18544_),
    .A2(\icache.lce.lce_cmd_inst.data_r [383]),
    .ZN(_18573_));
 OR3_X1 _45441_ (.A1(_15355_),
    .A2(_15356_),
    .A3(_15424_),
    .ZN(_18574_));
 OR3_X1 _45442_ (.A1(_15360_),
    .A2(_15363_),
    .A3(_17068_),
    .ZN(_18575_));
 AND3_X1 _45443_ (.A1(_18574_),
    .A2(_18575_),
    .A3(_15940_),
    .ZN(_18576_));
 OAI21_X2 _45444_ (.A(_17554_),
    .B1(_15373_),
    .B2(_15376_),
    .ZN(_18577_));
 OAI21_X2 _45445_ (.A(_15650_),
    .B1(_15381_),
    .B2(_15382_),
    .ZN(_18578_));
 AOI21_X1 _45446_ (.A(_18531_),
    .B1(_18577_),
    .B2(_18578_),
    .ZN(_18579_));
 NOR2_X2 _45447_ (.A1(_18576_),
    .A2(_18579_),
    .ZN(_18580_));
 OAI21_X1 _45448_ (.A(_18573_),
    .B1(_18580_),
    .B2(_18572_),
    .ZN(_05203_));
 NAND2_X1 _45449_ (.A1(_18544_),
    .A2(\icache.lce.lce_cmd_inst.data_r [384]),
    .ZN(_18581_));
 OAI21_X2 _45450_ (.A(_16396_),
    .B1(_15307_),
    .B2(_15309_),
    .ZN(_18582_));
 NAND2_X1 _45451_ (.A1(_15747_),
    .A2(_15325_),
    .ZN(_18583_));
 OAI211_X4 _45452_ (.A(_18583_),
    .B(_15610_),
    .C1(_15721_),
    .C2(\icache.data_mems_5__data_mem.data_o [0]),
    .ZN(_18584_));
 AOI21_X2 _45453_ (.A(_17300_),
    .B1(_18582_),
    .B2(_18584_),
    .ZN(_18585_));
 OAI21_X2 _45454_ (.A(_17554_),
    .B1(_15345_),
    .B2(_15347_),
    .ZN(_18586_));
 OAI21_X2 _45455_ (.A(_15650_),
    .B1(_15336_),
    .B2(_15339_),
    .ZN(_18587_));
 AOI21_X2 _45456_ (.A(_18531_),
    .B1(_18586_),
    .B2(_18587_),
    .ZN(_18588_));
 NOR2_X4 _45457_ (.A1(_18585_),
    .A2(_18588_),
    .ZN(_18589_));
 OAI21_X1 _45458_ (.A(_18581_),
    .B1(_18589_),
    .B2(_18572_),
    .ZN(_05204_));
 NAND2_X1 _45459_ (.A1(_18544_),
    .A2(\icache.lce.lce_cmd_inst.data_r [385]),
    .ZN(_18590_));
 OR2_X1 _45460_ (.A1(_15714_),
    .A2(\icache.data_mems_4__data_mem.data_o [1]),
    .ZN(_18591_));
 NAND2_X1 _45461_ (.A1(_16667_),
    .A2(_16408_),
    .ZN(_18592_));
 NAND2_X1 _45462_ (.A1(_18591_),
    .A2(_18592_),
    .ZN(_18593_));
 NAND2_X1 _45463_ (.A1(_18593_),
    .A2(_15770_),
    .ZN(_18594_));
 NAND2_X1 _45464_ (.A1(_15398_),
    .A2(_18019_),
    .ZN(_18595_));
 NAND2_X1 _45465_ (.A1(_16672_),
    .A2(_15402_),
    .ZN(_18596_));
 NAND2_X1 _45466_ (.A1(_18595_),
    .A2(_18596_),
    .ZN(_18597_));
 NAND2_X1 _45467_ (.A1(_18597_),
    .A2(_15514_),
    .ZN(_18598_));
 NAND3_X1 _45468_ (.A1(_18594_),
    .A2(_18598_),
    .A3(_15409_),
    .ZN(_18599_));
 OR2_X1 _45469_ (.A1(_15876_),
    .A2(\icache.data_mems_0__data_mem.data_o [1]),
    .ZN(_18600_));
 NAND2_X1 _45470_ (.A1(_16678_),
    .A2(_16067_),
    .ZN(_18601_));
 AND3_X1 _45471_ (.A1(_18600_),
    .A2(_18601_),
    .A3(_15463_),
    .ZN(_18602_));
 NAND2_X1 _45472_ (.A1(_16155_),
    .A2(\icache.data_mems_2__data_mem.data_o [1]),
    .ZN(_18603_));
 NAND2_X1 _45473_ (.A1(_15606_),
    .A2(\icache.data_mems_3__data_mem.data_o [1]),
    .ZN(_18604_));
 AOI21_X1 _45474_ (.A(_16634_),
    .B1(_18603_),
    .B2(_18604_),
    .ZN(_18605_));
 OAI21_X1 _45475_ (.A(_16640_),
    .B1(_18602_),
    .B2(_18605_),
    .ZN(_18606_));
 AND2_X2 _45476_ (.A1(_18599_),
    .A2(_18606_),
    .ZN(_18607_));
 OAI21_X1 _45477_ (.A(_18590_),
    .B1(_18607_),
    .B2(_18572_),
    .ZN(_05205_));
 NAND2_X1 _45478_ (.A1(_18544_),
    .A2(\icache.lce.lce_cmd_inst.data_r [386]),
    .ZN(_18608_));
 NOR2_X1 _45479_ (.A1(_16698_),
    .A2(_16867_),
    .ZN(_18609_));
 AND2_X1 _45480_ (.A1(_15438_),
    .A2(\icache.data_mems_5__data_mem.data_o [2]),
    .ZN(_18610_));
 OAI21_X2 _45481_ (.A(_16865_),
    .B1(_18609_),
    .B2(_18610_),
    .ZN(_18611_));
 OR2_X1 _45482_ (.A1(_15776_),
    .A2(\icache.data_mems_6__data_mem.data_o [2]),
    .ZN(_18612_));
 NAND2_X2 _45483_ (.A1(_16693_),
    .A2(_16169_),
    .ZN(_18613_));
 NAND3_X2 _45484_ (.A1(_18612_),
    .A2(_18613_),
    .A3(_17236_),
    .ZN(_18614_));
 AOI21_X2 _45485_ (.A(_17300_),
    .B1(_18611_),
    .B2(_18614_),
    .ZN(_18615_));
 NOR2_X1 _45486_ (.A1(_16690_),
    .A2(_15443_),
    .ZN(_18616_));
 AND2_X1 _45487_ (.A1(_15738_),
    .A2(\icache.data_mems_1__data_mem.data_o [2]),
    .ZN(_18617_));
 OAI21_X2 _45488_ (.A(_16865_),
    .B1(_18616_),
    .B2(_18617_),
    .ZN(_18618_));
 OR2_X1 _45489_ (.A1(_15457_),
    .A2(\icache.data_mems_2__data_mem.data_o [2]),
    .ZN(_18619_));
 NAND2_X1 _45490_ (.A1(_16685_),
    .A2(_16112_),
    .ZN(_18620_));
 NAND3_X2 _45491_ (.A1(_18619_),
    .A2(_18620_),
    .A3(_17236_),
    .ZN(_18621_));
 AOI21_X2 _45492_ (.A(_18531_),
    .B1(_18618_),
    .B2(_18621_),
    .ZN(_18622_));
 NOR2_X4 _45493_ (.A1(_18615_),
    .A2(_18622_),
    .ZN(_18623_));
 OAI21_X1 _45494_ (.A(_18608_),
    .B1(_18623_),
    .B2(_18572_),
    .ZN(_05206_));
 NAND2_X1 _45495_ (.A1(_18544_),
    .A2(\icache.lce.lce_cmd_inst.data_r [387]),
    .ZN(_18624_));
 NOR2_X2 _45496_ (.A1(_16709_),
    .A2(_15435_),
    .ZN(_18625_));
 AND2_X1 _45497_ (.A1(_15471_),
    .A2(\icache.data_mems_7__data_mem.data_o [3]),
    .ZN(_18626_));
 OAI21_X1 _45498_ (.A(_15432_),
    .B1(_18625_),
    .B2(_18626_),
    .ZN(_18627_));
 OR2_X1 _45499_ (.A1(_15362_),
    .A2(\icache.data_mems_4__data_mem.data_o [3]),
    .ZN(_18628_));
 NAND2_X1 _45500_ (.A1(_16704_),
    .A2(_15714_),
    .ZN(_18629_));
 NAND3_X2 _45501_ (.A1(_18628_),
    .A2(_18629_),
    .A3(_15369_),
    .ZN(_18630_));
 AND3_X1 _45502_ (.A1(_18627_),
    .A2(_15655_),
    .A3(_18630_),
    .ZN(_18631_));
 NAND2_X2 _45503_ (.A1(_15372_),
    .A2(\icache.data_mems_0__data_mem.data_o [3]),
    .ZN(_18632_));
 OAI211_X4 _45504_ (.A(_18632_),
    .B(_15673_),
    .C1(_15674_),
    .C2(_16718_),
    .ZN(_18633_));
 NAND2_X1 _45505_ (.A1(_15398_),
    .A2(\icache.data_mems_2__data_mem.data_o [3]),
    .ZN(_18634_));
 NAND2_X1 _45506_ (.A1(_15955_),
    .A2(\icache.data_mems_3__data_mem.data_o [3]),
    .ZN(_18635_));
 NAND3_X1 _45507_ (.A1(_18634_),
    .A2(_17511_),
    .A3(_18635_),
    .ZN(_18636_));
 AOI21_X1 _45508_ (.A(_18419_),
    .B1(_18633_),
    .B2(_18636_),
    .ZN(_18637_));
 OR2_X4 _45509_ (.A1(_18631_),
    .A2(_18637_),
    .ZN(_18638_));
 OAI21_X1 _45510_ (.A(_18624_),
    .B1(_18638_),
    .B2(_18572_),
    .ZN(_05207_));
 NAND2_X1 _45511_ (.A1(_18544_),
    .A2(\icache.lce.lce_cmd_inst.data_r [388]),
    .ZN(_18639_));
 NOR2_X1 _45512_ (.A1(_16732_),
    .A2(_15533_),
    .ZN(_18640_));
 AND2_X1 _45513_ (.A1(_15390_),
    .A2(\icache.data_mems_5__data_mem.data_o [4]),
    .ZN(_18641_));
 OR3_X1 _45514_ (.A1(_18640_),
    .A2(_18641_),
    .A3(_15424_),
    .ZN(_18642_));
 NAND2_X1 _45515_ (.A1(_15719_),
    .A2(\icache.data_mems_6__data_mem.data_o [4]),
    .ZN(_18643_));
 OAI211_X1 _45516_ (.A(_18643_),
    .B(_15321_),
    .C1(_16035_),
    .C2(_16727_),
    .ZN(_18644_));
 AND3_X1 _45517_ (.A1(_18642_),
    .A2(_16033_),
    .A3(_18644_),
    .ZN(_18645_));
 NOR2_X1 _45518_ (.A1(_16737_),
    .A2(_15452_),
    .ZN(_18646_));
 AND2_X1 _45519_ (.A1(_15438_),
    .A2(\icache.data_mems_3__data_mem.data_o [4]),
    .ZN(_18647_));
 OAI21_X2 _45520_ (.A(_17554_),
    .B1(_18646_),
    .B2(_18647_),
    .ZN(_18648_));
 NAND2_X1 _45521_ (.A1(_15756_),
    .A2(_16742_),
    .ZN(_18649_));
 NAND2_X1 _45522_ (.A1(_16740_),
    .A2(_16169_),
    .ZN(_18650_));
 NAND3_X2 _45523_ (.A1(_18649_),
    .A2(_18650_),
    .A3(_15464_),
    .ZN(_18651_));
 AOI21_X2 _45524_ (.A(_18531_),
    .B1(_18648_),
    .B2(_18651_),
    .ZN(_18652_));
 NOR2_X4 _45525_ (.A1(_18645_),
    .A2(_18652_),
    .ZN(_18653_));
 OAI21_X1 _45526_ (.A(_18639_),
    .B1(_18653_),
    .B2(_18572_),
    .ZN(_05208_));
 NAND2_X1 _45527_ (.A1(_18544_),
    .A2(\icache.lce.lce_cmd_inst.data_r [389]),
    .ZN(_18654_));
 NOR2_X1 _45528_ (.A1(_16762_),
    .A2(_15478_),
    .ZN(_18655_));
 AND2_X1 _45529_ (.A1(_15876_),
    .A2(\icache.data_mems_1__data_mem.data_o [5]),
    .ZN(_18656_));
 OR3_X1 _45530_ (.A1(_18655_),
    .A2(_18656_),
    .A3(_15394_),
    .ZN(_18657_));
 NAND2_X1 _45531_ (.A1(_15756_),
    .A2(\icache.data_mems_2__data_mem.data_o [5]),
    .ZN(_18658_));
 NAND2_X1 _45532_ (.A1(_15443_),
    .A2(\icache.data_mems_3__data_mem.data_o [5]),
    .ZN(_18659_));
 NAND3_X1 _45533_ (.A1(_18658_),
    .A2(_16230_),
    .A3(_18659_),
    .ZN(_18660_));
 NAND2_X1 _45534_ (.A1(_18657_),
    .A2(_18660_),
    .ZN(_18661_));
 BUF_X16 _45535_ (.A(_15579_),
    .Z(_18662_));
 NAND2_X1 _45536_ (.A1(_18661_),
    .A2(_18662_),
    .ZN(_18663_));
 NAND2_X1 _45537_ (.A1(_15719_),
    .A2(\icache.data_mems_4__data_mem.data_o [5]),
    .ZN(_18664_));
 NAND2_X1 _45538_ (.A1(_15475_),
    .A2(\icache.data_mems_5__data_mem.data_o [5]),
    .ZN(_18665_));
 AND3_X2 _45539_ (.A1(_18664_),
    .A2(_16418_),
    .A3(_18665_),
    .ZN(_18666_));
 NAND2_X1 _45540_ (.A1(_15772_),
    .A2(_16753_),
    .ZN(_18667_));
 NAND2_X1 _45541_ (.A1(_16751_),
    .A2(_15402_),
    .ZN(_18668_));
 AOI21_X1 _45542_ (.A(_16227_),
    .B1(_18667_),
    .B2(_18668_),
    .ZN(_18669_));
 OAI21_X1 _45543_ (.A(_17971_),
    .B1(_18666_),
    .B2(_18669_),
    .ZN(_18670_));
 NAND2_X2 _45544_ (.A1(_18663_),
    .A2(_18670_),
    .ZN(_18671_));
 OAI21_X1 _45545_ (.A(_18654_),
    .B1(_18671_),
    .B2(_18572_),
    .ZN(_05209_));
 BUF_X8 _45546_ (.A(_18268_),
    .Z(_18672_));
 NAND2_X1 _45547_ (.A1(_18672_),
    .A2(\icache.lce.lce_cmd_inst.data_r [390]),
    .ZN(_18673_));
 NOR2_X1 _45548_ (.A1(_16780_),
    .A2(_15505_),
    .ZN(_18674_));
 AND2_X1 _45549_ (.A1(_15784_),
    .A2(\icache.data_mems_3__data_mem.data_o [6]),
    .ZN(_18675_));
 NOR2_X2 _45550_ (.A1(_18674_),
    .A2(_18675_),
    .ZN(_18676_));
 NOR2_X1 _45551_ (.A1(_18676_),
    .A2(_16512_),
    .ZN(_18677_));
 NAND2_X1 _45552_ (.A1(_15537_),
    .A2(\icache.data_mems_0__data_mem.data_o [6]),
    .ZN(_18678_));
 NAND2_X1 _45553_ (.A1(_15810_),
    .A2(\icache.data_mems_1__data_mem.data_o [6]),
    .ZN(_18679_));
 AOI21_X2 _45554_ (.A(_15477_),
    .B1(_18678_),
    .B2(_18679_),
    .ZN(_18680_));
 OAI21_X1 _45555_ (.A(_16438_),
    .B1(_18677_),
    .B2(_18680_),
    .ZN(_18681_));
 NAND2_X1 _45556_ (.A1(_15836_),
    .A2(\icache.data_mems_6__data_mem.data_o [6]),
    .ZN(_18682_));
 NAND2_X1 _45557_ (.A1(_15541_),
    .A2(\icache.data_mems_7__data_mem.data_o [6]),
    .ZN(_18683_));
 AOI21_X1 _45558_ (.A(_15673_),
    .B1(_18682_),
    .B2(_18683_),
    .ZN(_18684_));
 NAND2_X1 _45559_ (.A1(_15736_),
    .A2(\icache.data_mems_4__data_mem.data_o [6]),
    .ZN(_18685_));
 NAND2_X1 _45560_ (.A1(_15375_),
    .A2(\icache.data_mems_5__data_mem.data_o [6]),
    .ZN(_18686_));
 AOI21_X1 _45561_ (.A(_16324_),
    .B1(_18685_),
    .B2(_18686_),
    .ZN(_18687_));
 OAI21_X1 _45562_ (.A(_18366_),
    .B1(_18684_),
    .B2(_18687_),
    .ZN(_18688_));
 AND2_X4 _45563_ (.A1(_18681_),
    .A2(_18688_),
    .ZN(_18689_));
 OAI21_X1 _45564_ (.A(_18673_),
    .B1(_18689_),
    .B2(_18572_),
    .ZN(_05211_));
 NAND2_X1 _45565_ (.A1(_18672_),
    .A2(\icache.lce.lce_cmd_inst.data_r [295]),
    .ZN(_18690_));
 OAI21_X2 _45566_ (.A(_15712_),
    .B1(_16136_),
    .B2(_16137_),
    .ZN(_18691_));
 OAI21_X1 _45567_ (.A(_15332_),
    .B1(_16140_),
    .B2(_16141_),
    .ZN(_18692_));
 NAND3_X1 _45568_ (.A1(_18691_),
    .A2(_15905_),
    .A3(_18692_),
    .ZN(_18693_));
 OAI21_X2 _45569_ (.A(_17308_),
    .B1(_16145_),
    .B2(_16146_),
    .ZN(_18694_));
 NAND3_X2 _45570_ (.A1(_16148_),
    .A2(_16150_),
    .A3(_17236_),
    .ZN(_18695_));
 NAND3_X1 _45571_ (.A1(_18694_),
    .A2(_16390_),
    .A3(_18695_),
    .ZN(_18696_));
 NAND2_X2 _45572_ (.A1(_18693_),
    .A2(_18696_),
    .ZN(_18697_));
 OAI21_X1 _45573_ (.A(_18690_),
    .B1(_18697_),
    .B2(_18572_),
    .ZN(_05105_));
 NAND2_X1 _45574_ (.A1(_18672_),
    .A2(\icache.lce.lce_cmd_inst.data_r [296]),
    .ZN(_18698_));
 NOR3_X2 _45575_ (.A1(_16163_),
    .A2(_16164_),
    .A3(_17273_),
    .ZN(_18699_));
 AOI21_X2 _45576_ (.A(_17988_),
    .B1(_16167_),
    .B2(_16170_),
    .ZN(_18700_));
 OAI21_X1 _45577_ (.A(_17827_),
    .B1(_18699_),
    .B2(_18700_),
    .ZN(_18701_));
 OAI21_X1 _45578_ (.A(_15860_),
    .B1(_16159_),
    .B2(_16160_),
    .ZN(_18702_));
 OAI21_X1 _45579_ (.A(_15650_),
    .B1(_16156_),
    .B2(_16157_),
    .ZN(_18703_));
 NAND3_X1 _45580_ (.A1(_18702_),
    .A2(_18703_),
    .A3(_18470_),
    .ZN(_18704_));
 NAND2_X2 _45581_ (.A1(_18701_),
    .A2(_18704_),
    .ZN(_18705_));
 BUF_X4 _45582_ (.A(_18294_),
    .Z(_18706_));
 OAI21_X1 _45583_ (.A(_18698_),
    .B1(_18705_),
    .B2(_18706_),
    .ZN(_05106_));
 NAND2_X1 _45584_ (.A1(_18672_),
    .A2(\icache.lce.lce_cmd_inst.data_r [297]),
    .ZN(_18707_));
 NAND2_X1 _45585_ (.A1(_16188_),
    .A2(_17228_),
    .ZN(_18708_));
 NAND2_X1 _45586_ (.A1(_16194_),
    .A2(_18209_),
    .ZN(_18709_));
 NAND2_X1 _45587_ (.A1(_18708_),
    .A2(_18709_),
    .ZN(_18710_));
 NAND2_X1 _45588_ (.A1(_18710_),
    .A2(_18662_),
    .ZN(_18711_));
 NOR3_X1 _45589_ (.A1(_16176_),
    .A2(_16177_),
    .A3(_17981_),
    .ZN(_18712_));
 AOI21_X2 _45590_ (.A(_15740_),
    .B1(_16180_),
    .B2(_16182_),
    .ZN(_18713_));
 OAI21_X1 _45591_ (.A(_17971_),
    .B1(_18712_),
    .B2(_18713_),
    .ZN(_18714_));
 NAND2_X2 _45592_ (.A1(_18711_),
    .A2(_18714_),
    .ZN(_18715_));
 OAI21_X1 _45593_ (.A(_18707_),
    .B1(_18715_),
    .B2(_18706_),
    .ZN(_05107_));
 NAND2_X1 _45594_ (.A1(_18672_),
    .A2(\icache.lce.lce_cmd_inst.data_r [298]),
    .ZN(_18716_));
 OAI21_X2 _45595_ (.A(_16099_),
    .B1(_16201_),
    .B2(_16202_),
    .ZN(_18717_));
 OAI21_X2 _45596_ (.A(_15370_),
    .B1(_16205_),
    .B2(_16206_),
    .ZN(_18718_));
 AOI21_X2 _45597_ (.A(_16956_),
    .B1(_18717_),
    .B2(_18718_),
    .ZN(_18719_));
 OAI21_X2 _45598_ (.A(_17308_),
    .B1(_16211_),
    .B2(_16212_),
    .ZN(_18720_));
 NAND3_X2 _45599_ (.A1(_16214_),
    .A2(_16216_),
    .A3(_17236_),
    .ZN(_18721_));
 AOI21_X2 _45600_ (.A(_17517_),
    .B1(_18720_),
    .B2(_18721_),
    .ZN(_18722_));
 NOR2_X4 _45601_ (.A1(_18719_),
    .A2(_18722_),
    .ZN(_18723_));
 OAI21_X1 _45602_ (.A(_18716_),
    .B1(_18723_),
    .B2(_18706_),
    .ZN(_05108_));
 NAND2_X1 _45603_ (.A1(_18672_),
    .A2(\icache.lce.lce_cmd_inst.data_r [299]),
    .ZN(_18724_));
 OAI21_X4 _45604_ (.A(_15853_),
    .B1(_16223_),
    .B2(_16225_),
    .ZN(_18725_));
 NAND3_X2 _45605_ (.A1(_16232_),
    .A2(_16234_),
    .A3(_15911_),
    .ZN(_18726_));
 AOI21_X2 _45606_ (.A(_17300_),
    .B1(_18725_),
    .B2(_18726_),
    .ZN(_18727_));
 NAND3_X2 _45607_ (.A1(_16239_),
    .A2(_16241_),
    .A3(_15988_),
    .ZN(_18728_));
 NAND3_X2 _45608_ (.A1(_16244_),
    .A2(_16246_),
    .A3(_15464_),
    .ZN(_18729_));
 AOI21_X2 _45609_ (.A(_18531_),
    .B1(_18728_),
    .B2(_18729_),
    .ZN(_18730_));
 NOR2_X4 _45610_ (.A1(_18727_),
    .A2(_18730_),
    .ZN(_18731_));
 OAI21_X1 _45611_ (.A(_18724_),
    .B1(_18731_),
    .B2(_18706_),
    .ZN(_05109_));
 NAND2_X1 _45612_ (.A1(_18672_),
    .A2(\icache.lce.lce_cmd_inst.data_r [300]),
    .ZN(_18732_));
 NAND2_X1 _45613_ (.A1(_16261_),
    .A2(_17228_),
    .ZN(_18733_));
 NAND2_X1 _45614_ (.A1(_16255_),
    .A2(_18209_),
    .ZN(_18734_));
 NAND2_X1 _45615_ (.A1(_18733_),
    .A2(_18734_),
    .ZN(_18735_));
 NAND2_X1 _45616_ (.A1(_18735_),
    .A2(_17960_),
    .ZN(_18736_));
 NAND3_X2 _45617_ (.A1(_16268_),
    .A2(_16270_),
    .A3(_15754_),
    .ZN(_18737_));
 NAND3_X2 _45618_ (.A1(_16273_),
    .A2(_16275_),
    .A3(_15761_),
    .ZN(_18738_));
 NAND3_X2 _45619_ (.A1(_18737_),
    .A2(_18738_),
    .A3(_18460_),
    .ZN(_18739_));
 NAND2_X4 _45620_ (.A1(_18736_),
    .A2(_18739_),
    .ZN(_18740_));
 OAI21_X1 _45621_ (.A(_18732_),
    .B1(_18740_),
    .B2(_18706_),
    .ZN(_05112_));
 NAND2_X1 _45622_ (.A1(_18672_),
    .A2(\icache.lce.lce_cmd_inst.data_r [301]),
    .ZN(_18741_));
 NAND2_X1 _45623_ (.A1(_16282_),
    .A2(_16341_),
    .ZN(_18742_));
 NAND2_X1 _45624_ (.A1(_16286_),
    .A2(_15587_),
    .ZN(_18743_));
 NAND2_X2 _45625_ (.A1(_18742_),
    .A2(_18743_),
    .ZN(_18744_));
 NAND2_X1 _45626_ (.A1(_18744_),
    .A2(_17960_),
    .ZN(_18745_));
 OAI21_X4 _45627_ (.A(_16386_),
    .B1(_16289_),
    .B2(_16290_),
    .ZN(_18746_));
 BUF_X16 _45628_ (.A(_15644_),
    .Z(_18747_));
 NAND3_X4 _45629_ (.A1(_16292_),
    .A2(_16293_),
    .A3(_15433_),
    .ZN(_18748_));
 NAND3_X4 _45630_ (.A1(_18746_),
    .A2(_18747_),
    .A3(_18748_),
    .ZN(_18749_));
 NAND2_X4 _45631_ (.A1(_18745_),
    .A2(_18749_),
    .ZN(_18750_));
 OAI21_X1 _45632_ (.A(_18741_),
    .B1(_18750_),
    .B2(_18706_),
    .ZN(_05113_));
 NAND2_X1 _45633_ (.A1(_18672_),
    .A2(\icache.lce.lce_cmd_inst.data_r [302]),
    .ZN(_18751_));
 NAND2_X1 _45634_ (.A1(_16300_),
    .A2(_15395_),
    .ZN(_18752_));
 NAND2_X1 _45635_ (.A1(_16304_),
    .A2(_15406_),
    .ZN(_18753_));
 AOI21_X1 _45636_ (.A(_16049_),
    .B1(_18752_),
    .B2(_18753_),
    .ZN(_18754_));
 AOI21_X1 _45637_ (.A(_16307_),
    .B1(_16311_),
    .B2(_16312_),
    .ZN(_18755_));
 AOI21_X2 _45638_ (.A(_15664_),
    .B1(_16308_),
    .B2(_16309_),
    .ZN(_18756_));
 NOR3_X1 _45639_ (.A1(_18755_),
    .A2(_18756_),
    .A3(_16314_),
    .ZN(_18757_));
 OR2_X4 _45640_ (.A1(_18754_),
    .A2(_18757_),
    .ZN(_18758_));
 OAI21_X1 _45641_ (.A(_18751_),
    .B1(_18758_),
    .B2(_18706_),
    .ZN(_05114_));
 NAND2_X1 _45642_ (.A1(_18672_),
    .A2(\icache.lce.lce_cmd_inst.data_r [303]),
    .ZN(_18759_));
 OAI21_X1 _45643_ (.A(_16099_),
    .B1(_16318_),
    .B2(_16320_),
    .ZN(_18760_));
 NAND2_X1 _45644_ (.A1(_15589_),
    .A2(_15909_),
    .ZN(_18761_));
 OAI211_X4 _45645_ (.A(_18761_),
    .B(_18164_),
    .C1(_18116_),
    .C2(\icache.data_mems_6__data_mem.data_o [47]),
    .ZN(_18762_));
 AOI21_X2 _45646_ (.A(_17300_),
    .B1(_18760_),
    .B2(_18762_),
    .ZN(_18763_));
 OAI21_X2 _45647_ (.A(_17308_),
    .B1(_16328_),
    .B2(_16329_),
    .ZN(_18764_));
 NAND3_X4 _45648_ (.A1(_16331_),
    .A2(_16332_),
    .A3(_16230_),
    .ZN(_18765_));
 AOI21_X2 _45649_ (.A(_18531_),
    .B1(_18764_),
    .B2(_18765_),
    .ZN(_18766_));
 NOR2_X4 _45650_ (.A1(_18763_),
    .A2(_18766_),
    .ZN(_18767_));
 OAI21_X1 _45651_ (.A(_18759_),
    .B1(_18767_),
    .B2(_18706_),
    .ZN(_05115_));
 BUF_X8 _45652_ (.A(_18268_),
    .Z(_18768_));
 NAND2_X1 _45653_ (.A1(_18768_),
    .A2(\icache.lce.lce_cmd_inst.data_r [304]),
    .ZN(_18769_));
 NAND2_X1 _45654_ (.A1(_16340_),
    .A2(_17228_),
    .ZN(_18770_));
 NAND2_X1 _45655_ (.A1(_16346_),
    .A2(_18209_),
    .ZN(_18771_));
 NAND2_X1 _45656_ (.A1(_18770_),
    .A2(_18771_),
    .ZN(_18772_));
 NAND2_X1 _45657_ (.A1(_18772_),
    .A2(_17960_),
    .ZN(_18773_));
 OAI21_X2 _45658_ (.A(_15754_),
    .B1(_16351_),
    .B2(_16352_),
    .ZN(_18774_));
 NAND3_X2 _45659_ (.A1(_16354_),
    .A2(_16355_),
    .A3(_15901_),
    .ZN(_18775_));
 NAND3_X2 _45660_ (.A1(_18774_),
    .A2(_18747_),
    .A3(_18775_),
    .ZN(_18776_));
 NAND2_X4 _45661_ (.A1(_18773_),
    .A2(_18776_),
    .ZN(_18777_));
 OAI21_X1 _45662_ (.A(_18769_),
    .B1(_18777_),
    .B2(_18706_),
    .ZN(_05116_));
 NAND2_X1 _45663_ (.A1(_18768_),
    .A2(\icache.lce.lce_cmd_inst.data_r [305]),
    .ZN(_18778_));
 AND3_X1 _45664_ (.A1(_16361_),
    .A2(_16362_),
    .A3(_15432_),
    .ZN(_18779_));
 AOI21_X2 _45665_ (.A(_15477_),
    .B1(_16364_),
    .B2(_16365_),
    .ZN(_18780_));
 OAI21_X1 _45666_ (.A(_16631_),
    .B1(_18779_),
    .B2(_18780_),
    .ZN(_18781_));
 NAND2_X1 _45667_ (.A1(_16370_),
    .A2(_15379_),
    .ZN(_18782_));
 NAND3_X2 _45668_ (.A1(_16373_),
    .A2(_15406_),
    .A3(_16374_),
    .ZN(_18783_));
 NAND3_X1 _45669_ (.A1(_18782_),
    .A2(_16372_),
    .A3(_18783_),
    .ZN(_18784_));
 AND2_X2 _45670_ (.A1(_18781_),
    .A2(_18784_),
    .ZN(_18785_));
 OAI21_X1 _45671_ (.A(_18778_),
    .B1(_18785_),
    .B2(_18706_),
    .ZN(_05117_));
 NAND2_X1 _45672_ (.A1(_18768_),
    .A2(\icache.lce.lce_cmd_inst.data_r [306]),
    .ZN(_18786_));
 AND3_X1 _45673_ (.A1(_16382_),
    .A2(_17511_),
    .A3(_16383_),
    .ZN(_18787_));
 AOI21_X2 _45674_ (.A(_15938_),
    .B1(_16379_),
    .B2(_16380_),
    .ZN(_18788_));
 NOR3_X2 _45675_ (.A1(_18787_),
    .A2(_18788_),
    .A3(_18132_),
    .ZN(_18789_));
 NOR3_X2 _45676_ (.A1(_16387_),
    .A2(_16388_),
    .A3(_17459_),
    .ZN(_18790_));
 AOI21_X2 _45677_ (.A(_17511_),
    .B1(_16392_),
    .B2(_16395_),
    .ZN(_18791_));
 NOR3_X2 _45678_ (.A1(_18790_),
    .A2(_18791_),
    .A3(_15849_),
    .ZN(_18792_));
 NOR2_X4 _45679_ (.A1(_18789_),
    .A2(_18792_),
    .ZN(_18793_));
 BUF_X8 _45680_ (.A(_18294_),
    .Z(_18794_));
 OAI21_X1 _45681_ (.A(_18786_),
    .B1(_18793_),
    .B2(_18794_),
    .ZN(_05118_));
 NAND2_X1 _45682_ (.A1(_18768_),
    .A2(\icache.lce.lce_cmd_inst.data_r [307]),
    .ZN(_18795_));
 NOR2_X1 _45683_ (.A1(_16404_),
    .A2(_17264_),
    .ZN(_18796_));
 AOI21_X1 _45684_ (.A(_16643_),
    .B1(_16407_),
    .B2(_16409_),
    .ZN(_18797_));
 NOR3_X1 _45685_ (.A1(_18796_),
    .A2(_16265_),
    .A3(_18797_),
    .ZN(_18798_));
 OR3_X2 _45686_ (.A1(_16412_),
    .A2(_16413_),
    .A3(_15320_),
    .ZN(_18799_));
 NAND2_X1 _45687_ (.A1(_16417_),
    .A2(_15425_),
    .ZN(_18800_));
 AOI21_X1 _45688_ (.A(_15579_),
    .B1(_18799_),
    .B2(_18800_),
    .ZN(_18801_));
 OR2_X4 _45689_ (.A1(_18798_),
    .A2(_18801_),
    .ZN(_18802_));
 OAI21_X1 _45690_ (.A(_18795_),
    .B1(_18802_),
    .B2(_18794_),
    .ZN(_05119_));
 NAND2_X1 _45691_ (.A1(_18768_),
    .A2(\icache.lce.lce_cmd_inst.data_r [308]),
    .ZN(_18803_));
 OAI211_X2 _45692_ (.A(_16430_),
    .B(_17511_),
    .C1(_15721_),
    .C2(_15713_),
    .ZN(_18804_));
 BUF_X8 _45693_ (.A(_15502_),
    .Z(_18805_));
 NAND3_X1 _45694_ (.A1(_16432_),
    .A2(_17264_),
    .A3(_16433_),
    .ZN(_18806_));
 AND3_X1 _45695_ (.A1(_18804_),
    .A2(_18805_),
    .A3(_18806_),
    .ZN(_18807_));
 OAI21_X2 _45696_ (.A(_16256_),
    .B1(_16423_),
    .B2(_16424_),
    .ZN(_18808_));
 NAND2_X1 _45697_ (.A1(_15729_),
    .A2(_17839_),
    .ZN(_18809_));
 OAI211_X4 _45698_ (.A(_18809_),
    .B(_15545_),
    .C1(_18116_),
    .C2(\icache.data_mems_0__data_mem.data_o [52]),
    .ZN(_18810_));
 AOI21_X2 _45699_ (.A(_18531_),
    .B1(_18808_),
    .B2(_18810_),
    .ZN(_18811_));
 NOR2_X4 _45700_ (.A1(_18807_),
    .A2(_18811_),
    .ZN(_18812_));
 OAI21_X1 _45701_ (.A(_18803_),
    .B1(_18812_),
    .B2(_18794_),
    .ZN(_05120_));
 NAND2_X1 _45702_ (.A1(_18768_),
    .A2(\icache.lce.lce_cmd_inst.data_r [309]),
    .ZN(_18813_));
 AOI211_X2 _45703_ (.A(_16229_),
    .B(_16439_),
    .C1(_15679_),
    .C2(_15743_),
    .ZN(_18814_));
 AOI21_X4 _45704_ (.A(_15369_),
    .B1(_16441_),
    .B2(_16442_),
    .ZN(_18815_));
 OR3_X2 _45705_ (.A1(_18814_),
    .A2(_15597_),
    .A3(_18815_),
    .ZN(_18816_));
 NAND2_X1 _45706_ (.A1(_16451_),
    .A2(_15343_),
    .ZN(_18817_));
 NAND2_X1 _45707_ (.A1(_16447_),
    .A2(_15594_),
    .ZN(_18818_));
 NAND2_X2 _45708_ (.A1(_18817_),
    .A2(_18818_),
    .ZN(_18819_));
 NAND2_X1 _45709_ (.A1(_18819_),
    .A2(_15598_),
    .ZN(_18820_));
 NAND2_X4 _45710_ (.A1(_18816_),
    .A2(_18820_),
    .ZN(_18821_));
 OAI21_X1 _45711_ (.A(_18813_),
    .B1(_18821_),
    .B2(_18794_),
    .ZN(_05121_));
 NAND2_X1 _45712_ (.A1(_18768_),
    .A2(\icache.lce.lce_cmd_inst.data_r [310]),
    .ZN(_18822_));
 NAND2_X1 _45713_ (.A1(_16462_),
    .A2(_16021_),
    .ZN(_18823_));
 NAND2_X1 _45714_ (.A1(_16458_),
    .A2(_15804_),
    .ZN(_18824_));
 AND3_X1 _45715_ (.A1(_18823_),
    .A2(_18824_),
    .A3(_16562_),
    .ZN(_18825_));
 OAI21_X1 _45716_ (.A(_15812_),
    .B1(_16466_),
    .B2(_16467_),
    .ZN(_18826_));
 NAND3_X2 _45717_ (.A1(_16469_),
    .A2(_16470_),
    .A3(_15342_),
    .ZN(_18827_));
 AOI21_X2 _45718_ (.A(_17517_),
    .B1(_18826_),
    .B2(_18827_),
    .ZN(_18828_));
 NOR2_X4 _45719_ (.A1(_18825_),
    .A2(_18828_),
    .ZN(_18829_));
 OAI21_X1 _45720_ (.A(_18822_),
    .B1(_18829_),
    .B2(_18794_),
    .ZN(_05123_));
 NAND2_X1 _45721_ (.A1(_18768_),
    .A2(\icache.lce.lce_cmd_inst.data_r [311]),
    .ZN(_18830_));
 OAI21_X4 _45722_ (.A(_16099_),
    .B1(_16482_),
    .B2(_16483_),
    .ZN(_18831_));
 NAND3_X4 _45723_ (.A1(_16485_),
    .A2(_16486_),
    .A3(_16578_),
    .ZN(_18832_));
 NAND3_X1 _45724_ (.A1(_18831_),
    .A2(_17567_),
    .A3(_18832_),
    .ZN(_18833_));
 NAND3_X4 _45725_ (.A1(_16475_),
    .A2(_16476_),
    .A3(_16262_),
    .ZN(_18834_));
 NAND3_X4 _45726_ (.A1(_16478_),
    .A2(_16479_),
    .A3(_15994_),
    .ZN(_18835_));
 NAND3_X1 _45727_ (.A1(_18834_),
    .A2(_18835_),
    .A3(_18470_),
    .ZN(_18836_));
 NAND2_X2 _45728_ (.A1(_18833_),
    .A2(_18836_),
    .ZN(_18837_));
 OAI21_X1 _45729_ (.A(_18830_),
    .B1(_18837_),
    .B2(_18794_),
    .ZN(_05124_));
 NAND2_X1 _45730_ (.A1(_18768_),
    .A2(\icache.lce.lce_cmd_inst.data_r [312]),
    .ZN(_18838_));
 NAND2_X1 _45731_ (.A1(_16497_),
    .A2(_16021_),
    .ZN(_18839_));
 NAND2_X1 _45732_ (.A1(_16493_),
    .A2(_15804_),
    .ZN(_18840_));
 AND3_X1 _45733_ (.A1(_18839_),
    .A2(_18840_),
    .A3(_15940_),
    .ZN(_18841_));
 OAI21_X1 _45734_ (.A(_15812_),
    .B1(_16503_),
    .B2(_16504_),
    .ZN(_18842_));
 OAI21_X4 _45735_ (.A(_15445_),
    .B1(_16500_),
    .B2(_16501_),
    .ZN(_18843_));
 AOI21_X2 _45736_ (.A(_18531_),
    .B1(_18842_),
    .B2(_18843_),
    .ZN(_18844_));
 NOR2_X4 _45737_ (.A1(_18841_),
    .A2(_18844_),
    .ZN(_18845_));
 OAI21_X1 _45738_ (.A(_18838_),
    .B1(_18845_),
    .B2(_18794_),
    .ZN(_05125_));
 NAND2_X1 _45739_ (.A1(_18768_),
    .A2(\icache.lce.lce_cmd_inst.data_r [313]),
    .ZN(_18846_));
 NOR2_X1 _45740_ (.A1(_16511_),
    .A2(_15425_),
    .ZN(_18847_));
 AOI21_X1 _45741_ (.A(_16634_),
    .B1(_16514_),
    .B2(_16515_),
    .ZN(_18848_));
 NOR3_X1 _45742_ (.A1(_18847_),
    .A2(_15724_),
    .A3(_18848_),
    .ZN(_18849_));
 NAND2_X1 _45743_ (.A1(_16524_),
    .A2(_16195_),
    .ZN(_18850_));
 NAND2_X1 _45744_ (.A1(_16520_),
    .A2(_16541_),
    .ZN(_18851_));
 AOI21_X1 _45745_ (.A(_18419_),
    .B1(_18850_),
    .B2(_18851_),
    .ZN(_18852_));
 OR2_X4 _45746_ (.A1(_18849_),
    .A2(_18852_),
    .ZN(_18853_));
 OAI21_X1 _45747_ (.A(_18846_),
    .B1(_18853_),
    .B2(_18794_),
    .ZN(_05126_));
 BUF_X8 _45748_ (.A(_18268_),
    .Z(_18854_));
 NAND2_X1 _45749_ (.A1(_18854_),
    .A2(\icache.lce.lce_cmd_inst.data_r [292]),
    .ZN(_18855_));
 AOI21_X2 _45750_ (.A(_15379_),
    .B1(_16084_),
    .B2(_16086_),
    .ZN(_18856_));
 AOI21_X2 _45751_ (.A(_18164_),
    .B1(_16089_),
    .B2(_16091_),
    .ZN(_18857_));
 OAI21_X1 _45752_ (.A(_18324_),
    .B1(_18856_),
    .B2(_18857_),
    .ZN(_18858_));
 NAND3_X2 _45753_ (.A1(_16073_),
    .A2(_16075_),
    .A3(_15754_),
    .ZN(_18859_));
 NAND3_X2 _45754_ (.A1(_16078_),
    .A2(_16080_),
    .A3(_15761_),
    .ZN(_18860_));
 NAND3_X1 _45755_ (.A1(_18859_),
    .A2(_18860_),
    .A3(_18460_),
    .ZN(_18861_));
 NAND2_X2 _45756_ (.A1(_18858_),
    .A2(_18861_),
    .ZN(_18862_));
 OAI21_X1 _45757_ (.A(_18855_),
    .B1(_18862_),
    .B2(_18794_),
    .ZN(_05102_));
 NAND2_X1 _45758_ (.A1(_18854_),
    .A2(\icache.lce.lce_cmd_inst.data_r [293]),
    .ZN(_18863_));
 OAI21_X2 _45759_ (.A(_16099_),
    .B1(_16096_),
    .B2(_16097_),
    .ZN(_18864_));
 OAI21_X2 _45760_ (.A(_15370_),
    .B1(_16101_),
    .B2(_16102_),
    .ZN(_18865_));
 AOI21_X2 _45761_ (.A(_17300_),
    .B1(_18864_),
    .B2(_18865_),
    .ZN(_18866_));
 BUF_X16 _45762_ (.A(_15367_),
    .Z(_18867_));
 OAI21_X1 _45763_ (.A(_17308_),
    .B1(_16106_),
    .B2(_16107_),
    .ZN(_18868_));
 NAND3_X2 _45764_ (.A1(_16110_),
    .A2(_16113_),
    .A3(_16230_),
    .ZN(_18869_));
 AOI21_X1 _45765_ (.A(_18867_),
    .B1(_18868_),
    .B2(_18869_),
    .ZN(_18870_));
 NOR2_X2 _45766_ (.A1(_18866_),
    .A2(_18870_),
    .ZN(_18871_));
 OAI21_X1 _45767_ (.A(_18863_),
    .B1(_18871_),
    .B2(_18794_),
    .ZN(_05103_));
 NAND2_X1 _45768_ (.A1(_18854_),
    .A2(\icache.lce.lce_cmd_inst.data_r [294]),
    .ZN(_18872_));
 OR3_X1 _45769_ (.A1(_16126_),
    .A2(_16127_),
    .A3(_15320_),
    .ZN(_18873_));
 OR3_X1 _45770_ (.A1(_16130_),
    .A2(_16131_),
    .A3(_17068_),
    .ZN(_18874_));
 AOI21_X1 _45771_ (.A(_16049_),
    .B1(_18873_),
    .B2(_18874_),
    .ZN(_18875_));
 OAI21_X2 _45772_ (.A(_15812_),
    .B1(_16119_),
    .B2(_16120_),
    .ZN(_18876_));
 NAND2_X1 _45773_ (.A1(_16123_),
    .A2(_15751_),
    .ZN(_18877_));
 OAI211_X2 _45774_ (.A(_18877_),
    .B(_16226_),
    .C1(_16015_),
    .C2(\icache.data_mems_6__data_mem.data_o [38]),
    .ZN(_18878_));
 AND3_X1 _45775_ (.A1(_18876_),
    .A2(_15819_),
    .A3(_18878_),
    .ZN(_18879_));
 OR2_X4 _45776_ (.A1(_18875_),
    .A2(_18879_),
    .ZN(_18880_));
 BUF_X8 _45777_ (.A(_18294_),
    .Z(_18881_));
 OAI21_X1 _45778_ (.A(_18872_),
    .B1(_18880_),
    .B2(_18881_),
    .ZN(_05104_));
 NAND2_X1 _45779_ (.A1(_18854_),
    .A2(\icache.lce.lce_cmd_inst.data_r [215]),
    .ZN(_18882_));
 NAND2_X1 _45780_ (.A1(_17136_),
    .A2(_18662_),
    .ZN(_18883_));
 NAND3_X1 _45781_ (.A1(_17141_),
    .A2(_17146_),
    .A3(_18470_),
    .ZN(_18884_));
 NAND2_X2 _45782_ (.A1(_18883_),
    .A2(_18884_),
    .ZN(_18885_));
 OAI21_X1 _45783_ (.A(_18882_),
    .B1(_18885_),
    .B2(_18881_),
    .ZN(_05017_));
 NAND2_X1 _45784_ (.A1(_18854_),
    .A2(\icache.lce.lce_cmd_inst.data_r [216]),
    .ZN(_18886_));
 OAI21_X1 _45785_ (.A(_18324_),
    .B1(_17155_),
    .B2(_17160_),
    .ZN(_18887_));
 NAND3_X1 _45786_ (.A1(_17165_),
    .A2(_17169_),
    .A3(_18460_),
    .ZN(_18888_));
 NAND2_X2 _45787_ (.A1(_18887_),
    .A2(_18888_),
    .ZN(_18889_));
 OAI21_X1 _45788_ (.A(_18886_),
    .B1(_18889_),
    .B2(_18881_),
    .ZN(_05018_));
 NAND2_X1 _45789_ (.A1(_18854_),
    .A2(\icache.lce.lce_cmd_inst.data_r [217]),
    .ZN(_18890_));
 NAND2_X1 _45790_ (.A1(_17184_),
    .A2(_18662_),
    .ZN(_18891_));
 OAI21_X1 _45791_ (.A(_17971_),
    .B1(_17189_),
    .B2(_17193_),
    .ZN(_18892_));
 NAND2_X2 _45792_ (.A1(_18891_),
    .A2(_18892_),
    .ZN(_18893_));
 OAI21_X1 _45793_ (.A(_18890_),
    .B1(_18893_),
    .B2(_18881_),
    .ZN(_05019_));
 NAND2_X1 _45794_ (.A1(_18854_),
    .A2(\icache.lce.lce_cmd_inst.data_r [218]),
    .ZN(_18894_));
 AOI21_X1 _45795_ (.A(_16049_),
    .B1(_17199_),
    .B2(_17202_),
    .ZN(_18895_));
 AOI21_X1 _45796_ (.A(_16314_),
    .B1(_17208_),
    .B2(_17214_),
    .ZN(_18896_));
 OR2_X4 _45797_ (.A1(_18895_),
    .A2(_18896_),
    .ZN(_18897_));
 OAI21_X1 _45798_ (.A(_18894_),
    .B1(_18897_),
    .B2(_18881_),
    .ZN(_05020_));
 NAND2_X1 _45799_ (.A1(_18854_),
    .A2(\icache.lce.lce_cmd_inst.data_r [219]),
    .ZN(_18898_));
 NAND3_X2 _45800_ (.A1(_17222_),
    .A2(_15735_),
    .A3(_17226_),
    .ZN(_18899_));
 NAND3_X2 _45801_ (.A1(_17232_),
    .A2(_16823_),
    .A3(_17237_),
    .ZN(_18900_));
 NAND2_X4 _45802_ (.A1(_18899_),
    .A2(_18900_),
    .ZN(_18901_));
 OAI21_X1 _45803_ (.A(_18898_),
    .B1(_18901_),
    .B2(_18881_),
    .ZN(_05021_));
 NAND2_X1 _45804_ (.A1(_18854_),
    .A2(\icache.lce.lce_cmd_inst.data_r [220]),
    .ZN(_18902_));
 BUF_X16 _45805_ (.A(_15328_),
    .Z(_18903_));
 AOI21_X2 _45806_ (.A(_18903_),
    .B1(_17243_),
    .B2(_17248_),
    .ZN(_18904_));
 AOI21_X2 _45807_ (.A(_18867_),
    .B1(_17253_),
    .B2(_17257_),
    .ZN(_18905_));
 NOR2_X4 _45808_ (.A1(_18904_),
    .A2(_18905_),
    .ZN(_18906_));
 OAI21_X1 _45809_ (.A(_18902_),
    .B1(_18906_),
    .B2(_18881_),
    .ZN(_05023_));
 NAND2_X1 _45810_ (.A1(_18854_),
    .A2(\icache.lce.lce_cmd_inst.data_r [221]),
    .ZN(_18907_));
 NOR3_X1 _45811_ (.A1(_17265_),
    .A2(_16265_),
    .A3(_17268_),
    .ZN(_18908_));
 AOI21_X1 _45812_ (.A(_16314_),
    .B1(_17274_),
    .B2(_17278_),
    .ZN(_18909_));
 OR2_X4 _45813_ (.A1(_18908_),
    .A2(_18909_),
    .ZN(_18910_));
 OAI21_X1 _45814_ (.A(_18907_),
    .B1(_18910_),
    .B2(_18881_),
    .ZN(_05024_));
 BUF_X4 _45815_ (.A(_18268_),
    .Z(_18911_));
 NAND2_X1 _45816_ (.A1(_18911_),
    .A2(\icache.lce.lce_cmd_inst.data_r [222]),
    .ZN(_18912_));
 NOR2_X1 _45817_ (.A1(_17289_),
    .A2(_15354_),
    .ZN(_18913_));
 AOI21_X2 _45818_ (.A(_18867_),
    .B1(_17293_),
    .B2(_17296_),
    .ZN(_18914_));
 NOR2_X4 _45819_ (.A1(_18913_),
    .A2(_18914_),
    .ZN(_18915_));
 OAI21_X1 _45820_ (.A(_18912_),
    .B1(_18915_),
    .B2(_18881_),
    .ZN(_05025_));
 NAND2_X1 _45821_ (.A1(_18911_),
    .A2(\icache.lce.lce_cmd_inst.data_r [223]),
    .ZN(_18916_));
 NAND3_X2 _45822_ (.A1(_17303_),
    .A2(_15735_),
    .A3(_17306_),
    .ZN(_18917_));
 BUF_X16 _45823_ (.A(_16012_),
    .Z(_18918_));
 NAND3_X2 _45824_ (.A1(_17311_),
    .A2(_18918_),
    .A3(_17315_),
    .ZN(_18919_));
 NAND2_X4 _45825_ (.A1(_18917_),
    .A2(_18919_),
    .ZN(_18920_));
 OAI21_X1 _45826_ (.A(_18916_),
    .B1(_18920_),
    .B2(_18881_),
    .ZN(_05026_));
 NAND2_X1 _45827_ (.A1(_18911_),
    .A2(\icache.lce.lce_cmd_inst.data_r [224]),
    .ZN(_18921_));
 BUF_X8 _45828_ (.A(_15833_),
    .Z(_18922_));
 OAI21_X1 _45829_ (.A(_18922_),
    .B1(_17322_),
    .B2(_17325_),
    .ZN(_18923_));
 NAND3_X1 _45830_ (.A1(_17330_),
    .A2(_17334_),
    .A3(_15849_),
    .ZN(_18924_));
 AND2_X4 _45831_ (.A1(_18923_),
    .A2(_18924_),
    .ZN(_18925_));
 BUF_X4 _45832_ (.A(_18294_),
    .Z(_18926_));
 OAI21_X1 _45833_ (.A(_18921_),
    .B1(_18925_),
    .B2(_18926_),
    .ZN(_05027_));
 NAND2_X1 _45834_ (.A1(_18911_),
    .A2(\icache.lce.lce_cmd_inst.data_r [225]),
    .ZN(_18927_));
 AND3_X2 _45835_ (.A1(_17340_),
    .A2(_18805_),
    .A3(_17344_),
    .ZN(_18928_));
 AOI21_X2 _45836_ (.A(_18867_),
    .B1(_17348_),
    .B2(_17351_),
    .ZN(_18929_));
 NOR2_X4 _45837_ (.A1(_18928_),
    .A2(_18929_),
    .ZN(_18930_));
 OAI21_X1 _45838_ (.A(_18927_),
    .B1(_18930_),
    .B2(_18926_),
    .ZN(_05028_));
 NAND2_X1 _45839_ (.A1(_18911_),
    .A2(\icache.lce.lce_cmd_inst.data_r [226]),
    .ZN(_18931_));
 OAI21_X1 _45840_ (.A(_18922_),
    .B1(_17357_),
    .B2(_17360_),
    .ZN(_18932_));
 NAND3_X1 _45841_ (.A1(_17363_),
    .A2(_17415_),
    .A3(_17366_),
    .ZN(_18933_));
 AND2_X4 _45842_ (.A1(_18932_),
    .A2(_18933_),
    .ZN(_18934_));
 OAI21_X1 _45843_ (.A(_18931_),
    .B1(_18934_),
    .B2(_18926_),
    .ZN(_05029_));
 NAND2_X1 _45844_ (.A1(_18911_),
    .A2(\icache.lce.lce_cmd_inst.data_r [227]),
    .ZN(_18935_));
 NAND2_X1 _45845_ (.A1(_17379_),
    .A2(_17960_),
    .ZN(_18936_));
 OR3_X2 _45846_ (.A1(_17383_),
    .A2(_17386_),
    .A3(_15655_),
    .ZN(_18937_));
 NAND2_X4 _45847_ (.A1(_18936_),
    .A2(_18937_),
    .ZN(_18938_));
 OAI21_X1 _45848_ (.A(_18935_),
    .B1(_18938_),
    .B2(_18926_),
    .ZN(_05030_));
 NAND2_X1 _45849_ (.A1(_18911_),
    .A2(\icache.lce.lce_cmd_inst.data_r [228]),
    .ZN(_18939_));
 AOI21_X2 _45850_ (.A(_18351_),
    .B1(_17392_),
    .B2(_17394_),
    .ZN(_18940_));
 AND3_X1 _45851_ (.A1(_17398_),
    .A2(_15430_),
    .A3(_17401_),
    .ZN(_18941_));
 OR2_X4 _45852_ (.A1(_18940_),
    .A2(_18941_),
    .ZN(_18942_));
 OAI21_X1 _45853_ (.A(_18939_),
    .B1(_18942_),
    .B2(_18926_),
    .ZN(_05031_));
 NAND2_X1 _45854_ (.A1(_18911_),
    .A2(\icache.lce.lce_cmd_inst.data_r [229]),
    .ZN(_18943_));
 NAND3_X1 _45855_ (.A1(_17409_),
    .A2(_17413_),
    .A3(_15409_),
    .ZN(_18944_));
 OAI21_X1 _45856_ (.A(_16640_),
    .B1(_17418_),
    .B2(_17421_),
    .ZN(_18945_));
 AND2_X4 _45857_ (.A1(_18944_),
    .A2(_18945_),
    .ZN(_18946_));
 OAI21_X1 _45858_ (.A(_18943_),
    .B1(_18946_),
    .B2(_18926_),
    .ZN(_05032_));
 NAND2_X1 _45859_ (.A1(_18911_),
    .A2(\icache.lce.lce_cmd_inst.data_r [230]),
    .ZN(_18947_));
 OAI21_X1 _45860_ (.A(_18922_),
    .B1(_17428_),
    .B2(_17431_),
    .ZN(_18948_));
 NAND3_X1 _45861_ (.A1(_17436_),
    .A2(_17415_),
    .A3(_17439_),
    .ZN(_18949_));
 AND2_X4 _45862_ (.A1(_18948_),
    .A2(_18949_),
    .ZN(_18950_));
 OAI21_X1 _45863_ (.A(_18947_),
    .B1(_18950_),
    .B2(_18926_),
    .ZN(_05034_));
 NAND2_X1 _45864_ (.A1(_18911_),
    .A2(\icache.lce.lce_cmd_inst.data_r [231]),
    .ZN(_18951_));
 OAI21_X1 _45865_ (.A(_16631_),
    .B1(_17444_),
    .B2(_17447_),
    .ZN(_18952_));
 NAND3_X1 _45866_ (.A1(_17452_),
    .A2(_16372_),
    .A3(_17455_),
    .ZN(_18953_));
 AND2_X4 _45867_ (.A1(_18952_),
    .A2(_18953_),
    .ZN(_18954_));
 OAI21_X1 _45868_ (.A(_18951_),
    .B1(_18954_),
    .B2(_18926_),
    .ZN(_05035_));
 BUF_X8 _45869_ (.A(_18268_),
    .Z(_18955_));
 NAND2_X1 _45870_ (.A1(_18955_),
    .A2(\icache.lce.lce_cmd_inst.data_r [232]),
    .ZN(_18956_));
 OAI21_X1 _45871_ (.A(_18922_),
    .B1(_17462_),
    .B2(_17465_),
    .ZN(_18957_));
 NAND3_X1 _45872_ (.A1(_17469_),
    .A2(_17415_),
    .A3(_17471_),
    .ZN(_18958_));
 AND2_X2 _45873_ (.A1(_18957_),
    .A2(_18958_),
    .ZN(_18959_));
 OAI21_X1 _45874_ (.A(_18956_),
    .B1(_18959_),
    .B2(_18926_),
    .ZN(_05036_));
 NAND2_X1 _45875_ (.A1(_18955_),
    .A2(\icache.lce.lce_cmd_inst.data_r [233]),
    .ZN(_18960_));
 AOI21_X4 _45876_ (.A(_18903_),
    .B1(_17477_),
    .B2(_17480_),
    .ZN(_18961_));
 AND3_X1 _45877_ (.A1(_17484_),
    .A2(_15724_),
    .A3(_17486_),
    .ZN(_18962_));
 NOR2_X4 _45878_ (.A1(_18961_),
    .A2(_18962_),
    .ZN(_18963_));
 OAI21_X1 _45879_ (.A(_18960_),
    .B1(_18963_),
    .B2(_18926_),
    .ZN(_05037_));
 NAND2_X1 _45880_ (.A1(_18955_),
    .A2(\icache.lce.lce_cmd_inst.data_r [234]),
    .ZN(_18964_));
 AND3_X1 _45881_ (.A1(_17512_),
    .A2(_18805_),
    .A3(_17515_),
    .ZN(_18965_));
 AOI21_X2 _45882_ (.A(_18867_),
    .B1(_17520_),
    .B2(_17523_),
    .ZN(_18966_));
 NOR2_X4 _45883_ (.A1(_18965_),
    .A2(_18966_),
    .ZN(_18967_));
 BUF_X8 _45884_ (.A(_18294_),
    .Z(_18968_));
 OAI21_X1 _45885_ (.A(_18964_),
    .B1(_18967_),
    .B2(_18968_),
    .ZN(_05038_));
 NAND2_X1 _45886_ (.A1(_18955_),
    .A2(\icache.lce.lce_cmd_inst.data_r [235]),
    .ZN(_18969_));
 NAND2_X1 _45887_ (.A1(_17536_),
    .A2(_17960_),
    .ZN(_18970_));
 OAI21_X2 _45888_ (.A(_18376_),
    .B1(_17540_),
    .B2(_17543_),
    .ZN(_18971_));
 NAND2_X4 _45889_ (.A1(_18970_),
    .A2(_18971_),
    .ZN(_18972_));
 OAI21_X1 _45890_ (.A(_18969_),
    .B1(_18972_),
    .B2(_18968_),
    .ZN(_05039_));
 NAND2_X1 _45891_ (.A1(_18955_),
    .A2(\icache.lce.lce_cmd_inst.data_r [236]),
    .ZN(_18973_));
 AOI21_X2 _45892_ (.A(_18903_),
    .B1(_17557_),
    .B2(_17560_),
    .ZN(_18974_));
 AOI21_X2 _45893_ (.A(_18867_),
    .B1(_17549_),
    .B2(_17552_),
    .ZN(_18975_));
 NOR2_X4 _45894_ (.A1(_18974_),
    .A2(_18975_),
    .ZN(_18976_));
 OAI21_X1 _45895_ (.A(_18973_),
    .B1(_18976_),
    .B2(_18968_),
    .ZN(_05040_));
 NAND2_X1 _45896_ (.A1(_18955_),
    .A2(\icache.lce.lce_cmd_inst.data_r [237]),
    .ZN(_18977_));
 AND3_X1 _45897_ (.A1(_15508_),
    .A2(_18805_),
    .A3(_15515_),
    .ZN(_18978_));
 AOI21_X2 _45898_ (.A(_18867_),
    .B1(_15521_),
    .B2(_15528_),
    .ZN(_18979_));
 NOR2_X4 _45899_ (.A1(_18978_),
    .A2(_18979_),
    .ZN(_18980_));
 OAI21_X1 _45900_ (.A(_18977_),
    .B1(_18980_),
    .B2(_18968_),
    .ZN(_05041_));
 NAND2_X1 _45901_ (.A1(_18955_),
    .A2(\icache.lce.lce_cmd_inst.data_r [238]),
    .ZN(_18981_));
 AND3_X1 _45902_ (.A1(_15536_),
    .A2(_18805_),
    .A3(_15546_),
    .ZN(_18982_));
 AOI21_X2 _45903_ (.A(_18867_),
    .B1(_15552_),
    .B2(_15558_),
    .ZN(_18983_));
 NOR2_X4 _45904_ (.A1(_18982_),
    .A2(_18983_),
    .ZN(_18984_));
 OAI21_X1 _45905_ (.A(_18981_),
    .B1(_18984_),
    .B2(_18968_),
    .ZN(_05042_));
 NAND2_X1 _45906_ (.A1(_18955_),
    .A2(\icache.lce.lce_cmd_inst.data_r [239]),
    .ZN(_18985_));
 NAND2_X1 _45907_ (.A1(_15596_),
    .A2(_18662_),
    .ZN(_18986_));
 NAND2_X1 _45908_ (.A1(_15578_),
    .A2(_15598_),
    .ZN(_18987_));
 NAND2_X2 _45909_ (.A1(_18986_),
    .A2(_18987_),
    .ZN(_18988_));
 OAI21_X1 _45910_ (.A(_18985_),
    .B1(_18988_),
    .B2(_18968_),
    .ZN(_05043_));
 NAND2_X1 _45911_ (.A1(_18955_),
    .A2(\icache.lce.lce_cmd_inst.data_r [240]),
    .ZN(_18989_));
 AND3_X1 _45912_ (.A1(_15611_),
    .A2(_15620_),
    .A3(_15940_),
    .ZN(_18990_));
 AOI21_X2 _45913_ (.A(_18867_),
    .B1(_15626_),
    .B2(_15632_),
    .ZN(_18991_));
 NOR2_X4 _45914_ (.A1(_18990_),
    .A2(_18991_),
    .ZN(_18992_));
 OAI21_X1 _45915_ (.A(_18989_),
    .B1(_18992_),
    .B2(_18968_),
    .ZN(_05045_));
 NAND2_X1 _45916_ (.A1(_18955_),
    .A2(\icache.lce.lce_cmd_inst.data_r [241]),
    .ZN(_18993_));
 AOI21_X2 _45917_ (.A(_18903_),
    .B1(_15639_),
    .B2(_15643_),
    .ZN(_18994_));
 AOI21_X2 _45918_ (.A(_18867_),
    .B1(_15649_),
    .B2(_15654_),
    .ZN(_18995_));
 NOR2_X4 _45919_ (.A1(_18994_),
    .A2(_18995_),
    .ZN(_18996_));
 OAI21_X1 _45920_ (.A(_18993_),
    .B1(_18996_),
    .B2(_18968_),
    .ZN(_05046_));
 BUF_X8 _45921_ (.A(_18268_),
    .Z(_18997_));
 NAND2_X1 _45922_ (.A1(_18997_),
    .A2(\icache.lce.lce_cmd_inst.data_r [242]),
    .ZN(_18998_));
 AND3_X1 _45923_ (.A1(_15676_),
    .A2(_15681_),
    .A3(_15940_),
    .ZN(_18999_));
 BUF_X16 _45924_ (.A(_15367_),
    .Z(_19000_));
 AOI21_X2 _45925_ (.A(_19000_),
    .B1(_15663_),
    .B2(_15668_),
    .ZN(_19001_));
 NOR2_X4 _45926_ (.A1(_18999_),
    .A2(_19001_),
    .ZN(_19002_));
 OAI21_X1 _45927_ (.A(_18998_),
    .B1(_19002_),
    .B2(_18968_),
    .ZN(_05047_));
 NAND2_X1 _45928_ (.A1(_18997_),
    .A2(\icache.lce.lce_cmd_inst.data_r [243]),
    .ZN(_19003_));
 AND3_X1 _45929_ (.A1(_15690_),
    .A2(_15474_),
    .A3(_15694_),
    .ZN(_19004_));
 BUF_X16 _45930_ (.A(_15833_),
    .Z(_19005_));
 AOI21_X2 _45931_ (.A(_19005_),
    .B1(_15698_),
    .B2(_15704_),
    .ZN(_19006_));
 NOR2_X4 _45932_ (.A1(_19004_),
    .A2(_19006_),
    .ZN(_19007_));
 OAI21_X1 _45933_ (.A(_19003_),
    .B1(_19007_),
    .B2(_18968_),
    .ZN(_05048_));
 NAND2_X1 _45934_ (.A1(_18997_),
    .A2(\icache.lce.lce_cmd_inst.data_r [244]),
    .ZN(_19008_));
 AOI21_X2 _45935_ (.A(_16956_),
    .B1(_15711_),
    .B2(_15717_),
    .ZN(_19009_));
 AND3_X1 _45936_ (.A1(_15723_),
    .A2(_16265_),
    .A3(_15730_),
    .ZN(_19010_));
 NOR2_X4 _45937_ (.A1(_19009_),
    .A2(_19010_),
    .ZN(_19011_));
 BUF_X8 _45938_ (.A(_18294_),
    .Z(_19012_));
 OAI21_X1 _45939_ (.A(_19008_),
    .B1(_19011_),
    .B2(_19012_),
    .ZN(_05049_));
 NAND2_X1 _45940_ (.A1(_18997_),
    .A2(\icache.lce.lce_cmd_inst.data_r [245]),
    .ZN(_19013_));
 OAI21_X2 _45941_ (.A(_18324_),
    .B1(_15741_),
    .B2(_15745_),
    .ZN(_19014_));
 NAND3_X2 _45942_ (.A1(_15755_),
    .A2(_15762_),
    .A3(_18460_),
    .ZN(_19015_));
 NAND2_X4 _45943_ (.A1(_19014_),
    .A2(_19015_),
    .ZN(_19016_));
 OAI21_X1 _45944_ (.A(_19013_),
    .B1(_19016_),
    .B2(_19012_),
    .ZN(_05050_));
 NAND2_X1 _45945_ (.A1(_18997_),
    .A2(\icache.lce.lce_cmd_inst.data_r [246]),
    .ZN(_19017_));
 AND3_X1 _45946_ (.A1(_15771_),
    .A2(_15780_),
    .A3(_16562_),
    .ZN(_19018_));
 AOI21_X1 _45947_ (.A(_19005_),
    .B1(_15786_),
    .B2(_15790_),
    .ZN(_19019_));
 NOR2_X2 _45948_ (.A1(_19018_),
    .A2(_19019_),
    .ZN(_19020_));
 OAI21_X1 _45949_ (.A(_19017_),
    .B1(_19020_),
    .B2(_19012_),
    .ZN(_05051_));
 NAND2_X1 _45950_ (.A1(_18997_),
    .A2(\icache.lce.lce_cmd_inst.data_r [247]),
    .ZN(_19021_));
 AND3_X1 _45951_ (.A1(_15798_),
    .A2(_15805_),
    .A3(_15503_),
    .ZN(_19022_));
 AOI21_X2 _45952_ (.A(_19000_),
    .B1(_15813_),
    .B2(_15818_),
    .ZN(_19023_));
 NOR2_X2 _45953_ (.A1(_19022_),
    .A2(_19023_),
    .ZN(_19024_));
 OAI21_X1 _45954_ (.A(_19021_),
    .B1(_19024_),
    .B2(_19012_),
    .ZN(_05052_));
 NAND2_X1 _45955_ (.A1(_18997_),
    .A2(\icache.lce.lce_cmd_inst.data_r [248]),
    .ZN(_19025_));
 AOI21_X1 _45956_ (.A(_18351_),
    .B1(_15827_),
    .B2(_15832_),
    .ZN(_19026_));
 AOI21_X1 _45957_ (.A(_18419_),
    .B1(_15842_),
    .B2(_15848_),
    .ZN(_19027_));
 OR2_X2 _45958_ (.A1(_19026_),
    .A2(_19027_),
    .ZN(_19028_));
 OAI21_X1 _45959_ (.A(_19025_),
    .B1(_19028_),
    .B2(_19012_),
    .ZN(_05053_));
 NAND2_X1 _45960_ (.A1(_18997_),
    .A2(\icache.lce.lce_cmd_inst.data_r [249]),
    .ZN(_19029_));
 AOI21_X2 _45961_ (.A(_16956_),
    .B1(_15856_),
    .B2(_15861_),
    .ZN(_19030_));
 AOI21_X2 _45962_ (.A(_19005_),
    .B1(_15866_),
    .B2(_15870_),
    .ZN(_19031_));
 NOR2_X4 _45963_ (.A1(_19030_),
    .A2(_19031_),
    .ZN(_19032_));
 OAI21_X1 _45964_ (.A(_19029_),
    .B1(_19032_),
    .B2(_19012_),
    .ZN(_05054_));
 NAND2_X1 _45965_ (.A1(_18997_),
    .A2(\icache.lce.lce_cmd_inst.data_r [250]),
    .ZN(_19033_));
 BUF_X16 _45966_ (.A(_15670_),
    .Z(_19034_));
 NAND2_X1 _45967_ (.A1(_15883_),
    .A2(_19034_),
    .ZN(_19035_));
 NAND2_X1 _45968_ (.A1(_15897_),
    .A2(_17567_),
    .ZN(_19036_));
 NAND2_X4 _45969_ (.A1(_19035_),
    .A2(_19036_),
    .ZN(_19037_));
 OAI21_X1 _45970_ (.A(_19033_),
    .B1(_19037_),
    .B2(_19012_),
    .ZN(_05056_));
 NAND2_X1 _45971_ (.A1(_18997_),
    .A2(\icache.lce.lce_cmd_inst.data_r [251]),
    .ZN(_19038_));
 NAND2_X2 _45972_ (.A1(_17498_),
    .A2(_18662_),
    .ZN(_19039_));
 OAI21_X2 _45973_ (.A(_17971_),
    .B1(_17503_),
    .B2(_17506_),
    .ZN(_19040_));
 NAND2_X4 _45974_ (.A1(_19039_),
    .A2(_19040_),
    .ZN(_19041_));
 OAI21_X1 _45975_ (.A(_19038_),
    .B1(_19041_),
    .B2(_19012_),
    .ZN(_05057_));
 BUF_X16 _45976_ (.A(_15301_),
    .Z(_19042_));
 BUF_X4 _45977_ (.A(_19042_),
    .Z(_19043_));
 NAND2_X1 _45978_ (.A1(_19043_),
    .A2(\icache.lce.lce_cmd_inst.data_r [252]),
    .ZN(_19044_));
 AOI21_X1 _45979_ (.A(_18351_),
    .B1(_15473_),
    .B2(_15481_),
    .ZN(_19045_));
 AND3_X1 _45980_ (.A1(_15490_),
    .A2(_15430_),
    .A3(_15498_),
    .ZN(_19046_));
 OR2_X4 _45981_ (.A1(_19045_),
    .A2(_19046_),
    .ZN(_19047_));
 OAI21_X1 _45982_ (.A(_19044_),
    .B1(_19047_),
    .B2(_19012_),
    .ZN(_05058_));
 NAND2_X1 _45983_ (.A1(_19043_),
    .A2(\icache.lce.lce_cmd_inst.data_r [253]),
    .ZN(_19048_));
 NAND3_X2 _45984_ (.A1(_15440_),
    .A2(_15735_),
    .A3(_15447_),
    .ZN(_19049_));
 NAND3_X2 _45985_ (.A1(_15456_),
    .A2(_18918_),
    .A3(_15465_),
    .ZN(_19050_));
 NAND2_X4 _45986_ (.A1(_19049_),
    .A2(_19050_),
    .ZN(_19051_));
 OAI21_X1 _45987_ (.A(_19048_),
    .B1(_19051_),
    .B2(_19012_),
    .ZN(_05059_));
 NAND2_X1 _45988_ (.A1(_19043_),
    .A2(\icache.lce.lce_cmd_inst.data_r [254]),
    .ZN(_19052_));
 AOI21_X2 _45989_ (.A(_16406_),
    .B1(_15396_),
    .B2(_15407_),
    .ZN(_19053_));
 AOI21_X1 _45990_ (.A(_16314_),
    .B1(_15416_),
    .B2(_15426_),
    .ZN(_19054_));
 OR2_X4 _45991_ (.A1(_19053_),
    .A2(_19054_),
    .ZN(_19055_));
 BUF_X16 _45992_ (.A(_15302_),
    .Z(_19056_));
 BUF_X4 _45993_ (.A(_19056_),
    .Z(_19057_));
 OAI21_X1 _45994_ (.A(_19052_),
    .B1(_19055_),
    .B2(_19057_),
    .ZN(_05060_));
 NAND2_X1 _45995_ (.A1(_19043_),
    .A2(\icache.lce.lce_cmd_inst.data_r [255]),
    .ZN(_19058_));
 AOI21_X2 _45996_ (.A(_18903_),
    .B1(_15377_),
    .B2(_15383_),
    .ZN(_19059_));
 AOI21_X2 _45997_ (.A(_19000_),
    .B1(_15357_),
    .B2(_15364_),
    .ZN(_19060_));
 NOR2_X4 _45998_ (.A1(_19059_),
    .A2(_19060_),
    .ZN(_19061_));
 OAI21_X1 _45999_ (.A(_19058_),
    .B1(_19061_),
    .B2(_19057_),
    .ZN(_05061_));
 NAND2_X1 _46000_ (.A1(_19043_),
    .A2(\icache.lce.lce_cmd_inst.data_r [256]),
    .ZN(_19062_));
 AND3_X1 _46001_ (.A1(_15312_),
    .A2(_18805_),
    .A3(_15326_),
    .ZN(_19063_));
 AOI21_X2 _46002_ (.A(_19000_),
    .B1(_15340_),
    .B2(_15348_),
    .ZN(_19064_));
 NOR2_X4 _46003_ (.A1(_19063_),
    .A2(_19064_),
    .ZN(_19065_));
 OAI21_X1 _46004_ (.A(_19062_),
    .B1(_19065_),
    .B2(_19057_),
    .ZN(_05062_));
 NAND2_X1 _46005_ (.A1(_19043_),
    .A2(\icache.lce.lce_cmd_inst.data_r [257]),
    .ZN(_19066_));
 NAND2_X1 _46006_ (.A1(_18593_),
    .A2(_16341_),
    .ZN(_19067_));
 NAND2_X1 _46007_ (.A1(_18597_),
    .A2(_15587_),
    .ZN(_19068_));
 NAND2_X1 _46008_ (.A1(_19067_),
    .A2(_19068_),
    .ZN(_19069_));
 NAND2_X1 _46009_ (.A1(_19069_),
    .A2(_19034_),
    .ZN(_19070_));
 AND3_X1 _46010_ (.A1(_18603_),
    .A2(_16418_),
    .A3(_18604_),
    .ZN(_19071_));
 AOI21_X2 _46011_ (.A(_16227_),
    .B1(_18600_),
    .B2(_18601_),
    .ZN(_19072_));
 OAI21_X2 _46012_ (.A(_18376_),
    .B1(_19071_),
    .B2(_19072_),
    .ZN(_19073_));
 NAND2_X4 _46013_ (.A1(_19070_),
    .A2(_19073_),
    .ZN(_19074_));
 OAI21_X1 _46014_ (.A(_19066_),
    .B1(_19074_),
    .B2(_19057_),
    .ZN(_05063_));
 NAND2_X1 _46015_ (.A1(_19043_),
    .A2(\icache.lce.lce_cmd_inst.data_r [258]),
    .ZN(_19075_));
 NOR3_X2 _46016_ (.A1(_18609_),
    .A2(_18610_),
    .A3(_16195_),
    .ZN(_19076_));
 AOI21_X2 _46017_ (.A(_15938_),
    .B1(_18612_),
    .B2(_18613_),
    .ZN(_19077_));
 OAI21_X2 _46018_ (.A(_18324_),
    .B1(_19076_),
    .B2(_19077_),
    .ZN(_19078_));
 OAI21_X2 _46019_ (.A(_15860_),
    .B1(_18616_),
    .B2(_18617_),
    .ZN(_19079_));
 NAND3_X2 _46020_ (.A1(_18619_),
    .A2(_18620_),
    .A3(_15994_),
    .ZN(_19080_));
 NAND3_X2 _46021_ (.A1(_19079_),
    .A2(_18747_),
    .A3(_19080_),
    .ZN(_19081_));
 NAND2_X4 _46022_ (.A1(_19078_),
    .A2(_19081_),
    .ZN(_19082_));
 OAI21_X1 _46023_ (.A(_19075_),
    .B1(_19082_),
    .B2(_19057_),
    .ZN(_05064_));
 NAND2_X1 _46024_ (.A1(_19043_),
    .A2(\icache.lce.lce_cmd_inst.data_r [259]),
    .ZN(_19083_));
 NAND2_X1 _46025_ (.A1(_15967_),
    .A2(\icache.data_mems_1__data_mem.data_o [3]),
    .ZN(_19084_));
 AOI21_X1 _46026_ (.A(_16307_),
    .B1(_18632_),
    .B2(_19084_),
    .ZN(_19085_));
 AOI21_X1 _46027_ (.A(_15812_),
    .B1(_18634_),
    .B2(_18635_),
    .ZN(_19086_));
 OR3_X1 _46028_ (.A1(_19085_),
    .A2(_19086_),
    .A3(_15655_),
    .ZN(_19087_));
 BUF_X16 _46029_ (.A(_16012_),
    .Z(_19088_));
 NOR3_X2 _46030_ (.A1(_18625_),
    .A2(_18626_),
    .A3(_15311_),
    .ZN(_19089_));
 AOI21_X2 _46031_ (.A(_16053_),
    .B1(_18628_),
    .B2(_18629_),
    .ZN(_19090_));
 OAI21_X2 _46032_ (.A(_19088_),
    .B1(_19089_),
    .B2(_19090_),
    .ZN(_19091_));
 NAND2_X4 _46033_ (.A1(_19087_),
    .A2(_19091_),
    .ZN(_19092_));
 OAI21_X1 _46034_ (.A(_19083_),
    .B1(_19092_),
    .B2(_19057_),
    .ZN(_05065_));
 NAND2_X1 _46035_ (.A1(_19043_),
    .A2(\icache.lce.lce_cmd_inst.data_r [260]),
    .ZN(_19093_));
 NOR3_X2 _46036_ (.A1(_18646_),
    .A2(_18647_),
    .A3(_17273_),
    .ZN(_19094_));
 AOI21_X2 _46037_ (.A(_17988_),
    .B1(_18649_),
    .B2(_18650_),
    .ZN(_19095_));
 OAI21_X2 _46038_ (.A(_17827_),
    .B1(_19094_),
    .B2(_19095_),
    .ZN(_19096_));
 OAI21_X2 _46039_ (.A(_15860_),
    .B1(_18640_),
    .B2(_18641_),
    .ZN(_19097_));
 NAND2_X1 _46040_ (.A1(_16727_),
    .A2(_17839_),
    .ZN(_19098_));
 OAI211_X2 _46041_ (.A(_19098_),
    .B(_17981_),
    .C1(_15324_),
    .C2(\icache.data_mems_6__data_mem.data_o [4]),
    .ZN(_19099_));
 NAND3_X2 _46042_ (.A1(_19097_),
    .A2(_19099_),
    .A3(_18470_),
    .ZN(_19100_));
 NAND2_X4 _46043_ (.A1(_19096_),
    .A2(_19100_),
    .ZN(_19101_));
 OAI21_X1 _46044_ (.A(_19093_),
    .B1(_19101_),
    .B2(_19057_),
    .ZN(_05067_));
 NAND2_X1 _46045_ (.A1(_19043_),
    .A2(\icache.lce.lce_cmd_inst.data_r [261]),
    .ZN(_19102_));
 OR3_X2 _46046_ (.A1(_18655_),
    .A2(_18656_),
    .A3(_15405_),
    .ZN(_19103_));
 NAND3_X2 _46047_ (.A1(_18658_),
    .A2(_15932_),
    .A3(_18659_),
    .ZN(_19104_));
 NAND3_X1 _46048_ (.A1(_19103_),
    .A2(_16438_),
    .A3(_19104_),
    .ZN(_19105_));
 AND3_X2 _46049_ (.A1(_18667_),
    .A2(_18668_),
    .A3(_16634_),
    .ZN(_19106_));
 AOI21_X1 _46050_ (.A(_15727_),
    .B1(_18664_),
    .B2(_18665_),
    .ZN(_19107_));
 OAI21_X1 _46051_ (.A(_18366_),
    .B1(_19106_),
    .B2(_19107_),
    .ZN(_19108_));
 AND2_X4 _46052_ (.A1(_19105_),
    .A2(_19108_),
    .ZN(_19109_));
 OAI21_X1 _46053_ (.A(_19102_),
    .B1(_19109_),
    .B2(_19057_),
    .ZN(_05068_));
 BUF_X4 _46054_ (.A(_19042_),
    .Z(_19110_));
 NAND2_X1 _46055_ (.A1(_19110_),
    .A2(\icache.lce.lce_cmd_inst.data_r [262]),
    .ZN(_19111_));
 NOR2_X1 _46056_ (.A1(_18676_),
    .A2(_17511_),
    .ZN(_19112_));
 AOI21_X1 _46057_ (.A(_15586_),
    .B1(_18678_),
    .B2(_18679_),
    .ZN(_19113_));
 OR3_X1 _46058_ (.A1(_19112_),
    .A2(_15597_),
    .A3(_19113_),
    .ZN(_19114_));
 AOI21_X1 _46059_ (.A(_16307_),
    .B1(_18685_),
    .B2(_18686_),
    .ZN(_19115_));
 AOI21_X2 _46060_ (.A(_15497_),
    .B1(_18682_),
    .B2(_18683_),
    .ZN(_19116_));
 OR3_X2 _46061_ (.A1(_19115_),
    .A2(_19116_),
    .A3(_15699_),
    .ZN(_19117_));
 NAND2_X4 _46062_ (.A1(_19114_),
    .A2(_19117_),
    .ZN(_19118_));
 OAI21_X1 _46063_ (.A(_19111_),
    .B1(_19118_),
    .B2(_19057_),
    .ZN(_05069_));
 NAND2_X1 _46064_ (.A1(_19110_),
    .A2(\icache.lce.lce_cmd_inst.data_r [263]),
    .ZN(_19119_));
 OR3_X1 _46065_ (.A1(_17898_),
    .A2(_17899_),
    .A3(_15544_),
    .ZN(_19120_));
 NAND2_X1 _46066_ (.A1(_17903_),
    .A2(_18209_),
    .ZN(_19121_));
 NAND2_X1 _46067_ (.A1(_19120_),
    .A2(_19121_),
    .ZN(_19122_));
 NAND2_X1 _46068_ (.A1(_19122_),
    .A2(_19034_),
    .ZN(_19123_));
 AOI21_X2 _46069_ (.A(_16014_),
    .B1(_17906_),
    .B2(_17907_),
    .ZN(_19124_));
 AOI21_X2 _46070_ (.A(_16227_),
    .B1(_17909_),
    .B2(_17910_),
    .ZN(_19125_));
 OAI21_X2 _46071_ (.A(_18376_),
    .B1(_19124_),
    .B2(_19125_),
    .ZN(_19126_));
 NAND2_X4 _46072_ (.A1(_19123_),
    .A2(_19126_),
    .ZN(_19127_));
 OAI21_X1 _46073_ (.A(_19119_),
    .B1(_19127_),
    .B2(_19057_),
    .ZN(_05070_));
 NAND2_X1 _46074_ (.A1(_19110_),
    .A2(\icache.lce.lce_cmd_inst.data_r [264]),
    .ZN(_19128_));
 NOR2_X1 _46075_ (.A1(_17917_),
    .A2(_15545_),
    .ZN(_19129_));
 AOI21_X1 _46076_ (.A(_16056_),
    .B1(_17919_),
    .B2(_17920_),
    .ZN(_19130_));
 OAI21_X1 _46077_ (.A(_16631_),
    .B1(_19129_),
    .B2(_19130_),
    .ZN(_19131_));
 AND3_X1 _46078_ (.A1(_17923_),
    .A2(_17924_),
    .A3(_16634_),
    .ZN(_19132_));
 AOI21_X1 _46079_ (.A(_15727_),
    .B1(_17926_),
    .B2(_17927_),
    .ZN(_19133_));
 OAI21_X1 _46080_ (.A(_16640_),
    .B1(_19132_),
    .B2(_19133_),
    .ZN(_19134_));
 AND2_X4 _46081_ (.A1(_19131_),
    .A2(_19134_),
    .ZN(_19135_));
 BUF_X4 _46082_ (.A(_19056_),
    .Z(_19136_));
 OAI21_X1 _46083_ (.A(_19128_),
    .B1(_19135_),
    .B2(_19136_),
    .ZN(_05071_));
 NAND2_X1 _46084_ (.A1(_19110_),
    .A2(\icache.lce.lce_cmd_inst.data_r [265]),
    .ZN(_19137_));
 NAND3_X2 _46085_ (.A1(_17933_),
    .A2(_17934_),
    .A3(_16099_),
    .ZN(_19138_));
 NAND3_X2 _46086_ (.A1(_17936_),
    .A2(_17937_),
    .A3(_16578_),
    .ZN(_19139_));
 NAND3_X2 _46087_ (.A1(_19138_),
    .A2(_19139_),
    .A3(_16143_),
    .ZN(_19140_));
 NAND3_X1 _46088_ (.A1(_17940_),
    .A2(_17941_),
    .A3(_16262_),
    .ZN(_19141_));
 NAND3_X1 _46089_ (.A1(_17943_),
    .A2(_17944_),
    .A3(_15610_),
    .ZN(_19142_));
 NAND3_X2 _46090_ (.A1(_19141_),
    .A2(_19142_),
    .A3(_18460_),
    .ZN(_19143_));
 NAND2_X4 _46091_ (.A1(_19140_),
    .A2(_19143_),
    .ZN(_19144_));
 OAI21_X1 _46092_ (.A(_19137_),
    .B1(_19144_),
    .B2(_19136_),
    .ZN(_05072_));
 NAND2_X1 _46093_ (.A1(_19110_),
    .A2(\icache.lce.lce_cmd_inst.data_r [266]),
    .ZN(_19145_));
 NOR3_X2 _46094_ (.A1(_17572_),
    .A2(_17573_),
    .A3(_15938_),
    .ZN(_19146_));
 AOI21_X2 _46095_ (.A(_17264_),
    .B1(_17575_),
    .B2(_17576_),
    .ZN(_19147_));
 NOR3_X2 _46096_ (.A1(_19146_),
    .A2(_19147_),
    .A3(_18132_),
    .ZN(_19148_));
 NOR3_X2 _46097_ (.A1(_17564_),
    .A2(_17565_),
    .A3(_17511_),
    .ZN(_19149_));
 AOI21_X2 _46098_ (.A(_17459_),
    .B1(_17568_),
    .B2(_17569_),
    .ZN(_19150_));
 NOR3_X2 _46099_ (.A1(_19149_),
    .A2(_19150_),
    .A3(_16033_),
    .ZN(_19151_));
 NOR2_X4 _46100_ (.A1(_19148_),
    .A2(_19151_),
    .ZN(_19152_));
 OAI21_X1 _46101_ (.A(_19145_),
    .B1(_19152_),
    .B2(_19136_),
    .ZN(_05073_));
 NAND2_X1 _46102_ (.A1(_19110_),
    .A2(\icache.lce.lce_cmd_inst.data_r [267]),
    .ZN(_19153_));
 AND3_X1 _46103_ (.A1(_17594_),
    .A2(_17595_),
    .A3(_15586_),
    .ZN(_19154_));
 AOI21_X2 _46104_ (.A(_15727_),
    .B1(_17591_),
    .B2(_17592_),
    .ZN(_19155_));
 NOR2_X4 _46105_ (.A1(_19154_),
    .A2(_19155_),
    .ZN(_19156_));
 NOR2_X1 _46106_ (.A1(_19156_),
    .A2(_16200_),
    .ZN(_19157_));
 NAND3_X4 _46107_ (.A1(_17583_),
    .A2(_17584_),
    .A3(_15988_),
    .ZN(_19158_));
 NAND3_X4 _46108_ (.A1(_17587_),
    .A2(_17588_),
    .A3(_15464_),
    .ZN(_19159_));
 AOI21_X2 _46109_ (.A(_19005_),
    .B1(_19158_),
    .B2(_19159_),
    .ZN(_19160_));
 NOR2_X4 _46110_ (.A1(_19157_),
    .A2(_19160_),
    .ZN(_19161_));
 OAI21_X1 _46111_ (.A(_19153_),
    .B1(_19161_),
    .B2(_19136_),
    .ZN(_05074_));
 NAND2_X1 _46112_ (.A1(_19110_),
    .A2(\icache.lce.lce_cmd_inst.data_r [268]),
    .ZN(_19162_));
 OR3_X1 _46113_ (.A1(_17600_),
    .A2(_17601_),
    .A3(_15544_),
    .ZN(_19163_));
 NAND3_X2 _46114_ (.A1(_17603_),
    .A2(_15545_),
    .A3(_17604_),
    .ZN(_19164_));
 NAND3_X1 _46115_ (.A1(_19163_),
    .A2(_16360_),
    .A3(_19164_),
    .ZN(_19165_));
 AND3_X1 _46116_ (.A1(_17607_),
    .A2(_17608_),
    .A3(_16643_),
    .ZN(_19166_));
 AOI21_X1 _46117_ (.A(_16324_),
    .B1(_17610_),
    .B2(_17611_),
    .ZN(_19167_));
 OAI21_X1 _46118_ (.A(_16640_),
    .B1(_19166_),
    .B2(_19167_),
    .ZN(_19168_));
 AND2_X4 _46119_ (.A1(_19165_),
    .A2(_19168_),
    .ZN(_19169_));
 OAI21_X1 _46120_ (.A(_19162_),
    .B1(_19169_),
    .B2(_19136_),
    .ZN(_05075_));
 NAND2_X1 _46121_ (.A1(_19110_),
    .A2(\icache.lce.lce_cmd_inst.data_r [269]),
    .ZN(_19170_));
 NAND2_X1 _46122_ (.A1(_17618_),
    .A2(_15770_),
    .ZN(_19171_));
 NAND2_X1 _46123_ (.A1(_17622_),
    .A2(_15514_),
    .ZN(_19172_));
 AOI21_X1 _46124_ (.A(_18351_),
    .B1(_19171_),
    .B2(_19172_),
    .ZN(_19173_));
 NAND2_X1 _46125_ (.A1(_17628_),
    .A2(_17273_),
    .ZN(_19174_));
 NAND3_X1 _46126_ (.A1(_17630_),
    .A2(_15673_),
    .A3(_17631_),
    .ZN(_19175_));
 AOI21_X1 _46127_ (.A(_18419_),
    .B1(_19174_),
    .B2(_19175_),
    .ZN(_19176_));
 OR2_X4 _46128_ (.A1(_19173_),
    .A2(_19176_),
    .ZN(_19177_));
 OAI21_X1 _46129_ (.A(_19170_),
    .B1(_19177_),
    .B2(_19136_),
    .ZN(_05076_));
 NAND2_X1 _46130_ (.A1(_19110_),
    .A2(\icache.lce.lce_cmd_inst.data_r [270]),
    .ZN(_19178_));
 BUF_X8 _46131_ (.A(_15408_),
    .Z(_19179_));
 NOR2_X1 _46132_ (.A1(_17640_),
    .A2(_16512_),
    .ZN(_19180_));
 AOI21_X1 _46133_ (.A(_15477_),
    .B1(_17642_),
    .B2(_17643_),
    .ZN(_19181_));
 OAI21_X1 _46134_ (.A(_19179_),
    .B1(_19180_),
    .B2(_19181_),
    .ZN(_19182_));
 BUF_X8 _46135_ (.A(_15314_),
    .Z(_19183_));
 NAND2_X1 _46136_ (.A1(_15443_),
    .A2(\icache.data_mems_3__data_mem.data_o [14]),
    .ZN(_19184_));
 AOI21_X1 _46137_ (.A(_17511_),
    .B1(_17646_),
    .B2(_19184_),
    .ZN(_19185_));
 AOI21_X1 _46138_ (.A(_15727_),
    .B1(_17648_),
    .B2(_17649_),
    .ZN(_19186_));
 OAI21_X1 _46139_ (.A(_19183_),
    .B1(_19185_),
    .B2(_19186_),
    .ZN(_19187_));
 AND2_X4 _46140_ (.A1(_19182_),
    .A2(_19187_),
    .ZN(_19188_));
 OAI21_X1 _46141_ (.A(_19178_),
    .B1(_19188_),
    .B2(_19136_),
    .ZN(_05078_));
 NAND2_X1 _46142_ (.A1(_19110_),
    .A2(\icache.lce.lce_cmd_inst.data_r [271]),
    .ZN(_19189_));
 AOI21_X2 _46143_ (.A(_15343_),
    .B1(_17661_),
    .B2(_17662_),
    .ZN(_19190_));
 AOI21_X2 _46144_ (.A(_17710_),
    .B1(_17664_),
    .B2(_17665_),
    .ZN(_19191_));
 OAI21_X2 _46145_ (.A(_18324_),
    .B1(_19190_),
    .B2(_19191_),
    .ZN(_19192_));
 NAND3_X2 _46146_ (.A1(_17654_),
    .A2(_17655_),
    .A3(_15754_),
    .ZN(_19193_));
 NAND3_X2 _46147_ (.A1(_17657_),
    .A2(_17658_),
    .A3(_15853_),
    .ZN(_19194_));
 NAND3_X2 _46148_ (.A1(_19193_),
    .A2(_19194_),
    .A3(_18460_),
    .ZN(_19195_));
 NAND2_X4 _46149_ (.A1(_19192_),
    .A2(_19195_),
    .ZN(_19196_));
 OAI21_X1 _46150_ (.A(_19189_),
    .B1(_19196_),
    .B2(_19136_),
    .ZN(_05079_));
 BUF_X4 _46151_ (.A(_19042_),
    .Z(_19197_));
 NAND2_X1 _46152_ (.A1(_19197_),
    .A2(\icache.lce.lce_cmd_inst.data_r [272]),
    .ZN(_19198_));
 OR3_X1 _46153_ (.A1(_17670_),
    .A2(_17671_),
    .A3(_15320_),
    .ZN(_19199_));
 NAND2_X1 _46154_ (.A1(_17675_),
    .A2(_15804_),
    .ZN(_19200_));
 AOI21_X1 _46155_ (.A(_16406_),
    .B1(_19199_),
    .B2(_19200_),
    .ZN(_19201_));
 AND3_X1 _46156_ (.A1(_17682_),
    .A2(_17683_),
    .A3(_15463_),
    .ZN(_19202_));
 AOI21_X1 _46157_ (.A(_15484_),
    .B1(_17679_),
    .B2(_17680_),
    .ZN(_19203_));
 NOR3_X1 _46158_ (.A1(_19202_),
    .A2(_19203_),
    .A3(_16314_),
    .ZN(_19204_));
 OR2_X4 _46159_ (.A1(_19201_),
    .A2(_19204_),
    .ZN(_19205_));
 OAI21_X1 _46160_ (.A(_19198_),
    .B1(_19205_),
    .B2(_19136_),
    .ZN(_05080_));
 NAND2_X1 _46161_ (.A1(_19197_),
    .A2(\icache.lce.lce_cmd_inst.data_r [273]),
    .ZN(_19206_));
 OR3_X1 _46162_ (.A1(_17688_),
    .A2(_17689_),
    .A3(_15544_),
    .ZN(_19207_));
 NAND2_X1 _46163_ (.A1(_17693_),
    .A2(_15567_),
    .ZN(_19208_));
 NAND2_X2 _46164_ (.A1(_19207_),
    .A2(_19208_),
    .ZN(_19209_));
 NAND2_X1 _46165_ (.A1(_19209_),
    .A2(_18662_),
    .ZN(_19210_));
 OAI21_X2 _46166_ (.A(_15761_),
    .B1(_17697_),
    .B2(_17698_),
    .ZN(_19211_));
 NAND3_X2 _46167_ (.A1(_17700_),
    .A2(_17701_),
    .A3(_15433_),
    .ZN(_19212_));
 NAND3_X4 _46168_ (.A1(_19211_),
    .A2(_18918_),
    .A3(_19212_),
    .ZN(_19213_));
 NAND2_X4 _46169_ (.A1(_19210_),
    .A2(_19213_),
    .ZN(_19214_));
 OAI21_X1 _46170_ (.A(_19206_),
    .B1(_19214_),
    .B2(_19136_),
    .ZN(_05081_));
 NAND2_X1 _46171_ (.A1(_19197_),
    .A2(\icache.lce.lce_cmd_inst.data_r [274]),
    .ZN(_19215_));
 AND3_X1 _46172_ (.A1(_17718_),
    .A2(_17719_),
    .A3(_15497_),
    .ZN(_19216_));
 AOI21_X1 _46173_ (.A(_15678_),
    .B1(_17715_),
    .B2(_17716_),
    .ZN(_19217_));
 NOR2_X2 _46174_ (.A1(_19216_),
    .A2(_19217_),
    .ZN(_19218_));
 NOR2_X1 _46175_ (.A1(_19218_),
    .A2(_15354_),
    .ZN(_19219_));
 NAND3_X2 _46176_ (.A1(_17707_),
    .A2(_17708_),
    .A3(_16578_),
    .ZN(_19220_));
 NAND3_X2 _46177_ (.A1(_17711_),
    .A2(_17712_),
    .A3(_17236_),
    .ZN(_19221_));
 AOI21_X2 _46178_ (.A(_19000_),
    .B1(_19220_),
    .B2(_19221_),
    .ZN(_19222_));
 NOR2_X4 _46179_ (.A1(_19219_),
    .A2(_19222_),
    .ZN(_19223_));
 BUF_X4 _46180_ (.A(_19056_),
    .Z(_19224_));
 OAI21_X1 _46181_ (.A(_19215_),
    .B1(_19223_),
    .B2(_19224_),
    .ZN(_05082_));
 NAND2_X1 _46182_ (.A1(_19197_),
    .A2(\icache.lce.lce_cmd_inst.data_r [275]),
    .ZN(_19225_));
 OR3_X1 _46183_ (.A1(_17724_),
    .A2(_17725_),
    .A3(_15424_),
    .ZN(_19226_));
 NAND3_X1 _46184_ (.A1(_17727_),
    .A2(_15425_),
    .A3(_17728_),
    .ZN(_19227_));
 AND3_X1 _46185_ (.A1(_19226_),
    .A2(_15474_),
    .A3(_19227_),
    .ZN(_19228_));
 NAND3_X2 _46186_ (.A1(_17733_),
    .A2(_17734_),
    .A3(_15988_),
    .ZN(_19229_));
 NAND3_X2 _46187_ (.A1(_17736_),
    .A2(_17737_),
    .A3(_15464_),
    .ZN(_19230_));
 AOI21_X4 _46188_ (.A(_19005_),
    .B1(_19229_),
    .B2(_19230_),
    .ZN(_19231_));
 NOR2_X4 _46189_ (.A1(_19228_),
    .A2(_19231_),
    .ZN(_19232_));
 OAI21_X1 _46190_ (.A(_19225_),
    .B1(_19232_),
    .B2(_19224_),
    .ZN(_05083_));
 NAND2_X1 _46191_ (.A1(_19197_),
    .A2(\icache.lce.lce_cmd_inst.data_r [276]),
    .ZN(_19233_));
 NOR2_X1 _46192_ (.A1(_17744_),
    .A2(_17459_),
    .ZN(_19234_));
 AOI21_X1 _46193_ (.A(_15331_),
    .B1(_17746_),
    .B2(_17747_),
    .ZN(_19235_));
 OR3_X1 _46194_ (.A1(_19234_),
    .A2(_16012_),
    .A3(_19235_),
    .ZN(_19236_));
 OAI21_X2 _46195_ (.A(_15754_),
    .B1(_17750_),
    .B2(_17751_),
    .ZN(_19237_));
 NAND2_X1 _46196_ (.A1(_17079_),
    .A2(_15479_),
    .ZN(_19238_));
 OAI211_X4 _46197_ (.A(_19238_),
    .B(_16578_),
    .C1(_18116_),
    .C2(\icache.data_mems_6__data_mem.data_o [20]),
    .ZN(_19239_));
 NAND3_X2 _46198_ (.A1(_19237_),
    .A2(_19239_),
    .A3(_18470_),
    .ZN(_19240_));
 NAND2_X4 _46199_ (.A1(_19236_),
    .A2(_19240_),
    .ZN(_19241_));
 OAI21_X1 _46200_ (.A(_19233_),
    .B1(_19241_),
    .B2(_19224_),
    .ZN(_05084_));
 NAND2_X1 _46201_ (.A1(_19197_),
    .A2(\icache.lce.lce_cmd_inst.data_r [277]),
    .ZN(_19242_));
 OAI21_X2 _46202_ (.A(_15660_),
    .B1(_17765_),
    .B2(_17766_),
    .ZN(_19243_));
 NAND2_X1 _46203_ (.A1(_17088_),
    .A2(_15421_),
    .ZN(_19244_));
 OAI211_X2 _46204_ (.A(_19244_),
    .B(_15378_),
    .C1(_15318_),
    .C2(\icache.data_mems_4__data_mem.data_o [21]),
    .ZN(_19245_));
 AND3_X1 _46205_ (.A1(_19243_),
    .A2(_19245_),
    .A3(_15522_),
    .ZN(_19246_));
 NAND3_X1 _46206_ (.A1(_17761_),
    .A2(_17459_),
    .A3(_17762_),
    .ZN(_19247_));
 NAND2_X1 _46207_ (.A1(_16253_),
    .A2(\icache.data_mems_1__data_mem.data_o [21]),
    .ZN(_19248_));
 OAI211_X2 _46208_ (.A(_19248_),
    .B(_15678_),
    .C1(_15909_),
    .C2(_17103_),
    .ZN(_19249_));
 AOI21_X1 _46209_ (.A(_18419_),
    .B1(_19247_),
    .B2(_19249_),
    .ZN(_19250_));
 OR2_X4 _46210_ (.A1(_19246_),
    .A2(_19250_),
    .ZN(_19251_));
 OAI21_X1 _46211_ (.A(_19242_),
    .B1(_19251_),
    .B2(_19224_),
    .ZN(_05085_));
 NAND2_X1 _46212_ (.A1(_19197_),
    .A2(\icache.lce.lce_cmd_inst.data_r [278]),
    .ZN(_19252_));
 NAND2_X1 _46213_ (.A1(_17779_),
    .A2(_16578_),
    .ZN(_19253_));
 NAND2_X1 _46214_ (.A1(_17775_),
    .A2(_15594_),
    .ZN(_19254_));
 NAND3_X1 _46215_ (.A1(_19253_),
    .A2(_19254_),
    .A3(_15409_),
    .ZN(_19255_));
 AOI21_X1 _46216_ (.A(_15673_),
    .B1(_17783_),
    .B2(_17784_),
    .ZN(_19256_));
 AOI21_X1 _46217_ (.A(_15678_),
    .B1(_17786_),
    .B2(_17787_),
    .ZN(_19257_));
 OAI21_X1 _46218_ (.A(_19183_),
    .B1(_19256_),
    .B2(_19257_),
    .ZN(_19258_));
 AND2_X4 _46219_ (.A1(_19255_),
    .A2(_19258_),
    .ZN(_19259_));
 OAI21_X1 _46220_ (.A(_19252_),
    .B1(_19259_),
    .B2(_19224_),
    .ZN(_05086_));
 NAND2_X1 _46221_ (.A1(_19197_),
    .A2(\icache.lce.lce_cmd_inst.data_r [279]),
    .ZN(_19260_));
 NOR3_X1 _46222_ (.A1(_17801_),
    .A2(_17802_),
    .A3(_16512_),
    .ZN(_19261_));
 AOI21_X2 _46223_ (.A(_17710_),
    .B1(_17804_),
    .B2(_17805_),
    .ZN(_19262_));
 OAI21_X2 _46224_ (.A(_17827_),
    .B1(_19261_),
    .B2(_19262_),
    .ZN(_19263_));
 AND3_X4 _46225_ (.A1(_17796_),
    .A2(_16418_),
    .A3(_17797_),
    .ZN(_19264_));
 AOI21_X4 _46226_ (.A(_16227_),
    .B1(_17793_),
    .B2(_17794_),
    .ZN(_19265_));
 OAI21_X2 _46227_ (.A(_19088_),
    .B1(_19264_),
    .B2(_19265_),
    .ZN(_19266_));
 NAND2_X4 _46228_ (.A1(_19263_),
    .A2(_19266_),
    .ZN(_19267_));
 OAI21_X1 _46229_ (.A(_19260_),
    .B1(_19267_),
    .B2(_19224_),
    .ZN(_05087_));
 NAND2_X1 _46230_ (.A1(_19197_),
    .A2(\icache.lce.lce_cmd_inst.data_r [280]),
    .ZN(_19268_));
 AOI21_X2 _46231_ (.A(_15379_),
    .B1(_17818_),
    .B2(_17819_),
    .ZN(_19269_));
 AOI21_X2 _46232_ (.A(_18164_),
    .B1(_17821_),
    .B2(_17822_),
    .ZN(_19270_));
 OAI21_X2 _46233_ (.A(_17827_),
    .B1(_19269_),
    .B2(_19270_),
    .ZN(_19271_));
 OAI21_X2 _46234_ (.A(_15754_),
    .B1(_17813_),
    .B2(_17814_),
    .ZN(_19272_));
 OAI21_X2 _46235_ (.A(_15761_),
    .B1(_17810_),
    .B2(_17811_),
    .ZN(_19273_));
 NAND3_X2 _46236_ (.A1(_19272_),
    .A2(_19273_),
    .A3(_18470_),
    .ZN(_19274_));
 NAND2_X4 _46237_ (.A1(_19271_),
    .A2(_19274_),
    .ZN(_19275_));
 OAI21_X1 _46238_ (.A(_19268_),
    .B1(_19275_),
    .B2(_19224_),
    .ZN(_05089_));
 NAND2_X1 _46239_ (.A1(_19197_),
    .A2(\icache.lce.lce_cmd_inst.data_r [281]),
    .ZN(_19276_));
 OAI21_X2 _46240_ (.A(_16256_),
    .B1(_17835_),
    .B2(_17836_),
    .ZN(_19277_));
 NAND3_X2 _46241_ (.A1(_17838_),
    .A2(_17840_),
    .A3(_17236_),
    .ZN(_19278_));
 AOI21_X2 _46242_ (.A(_18903_),
    .B1(_19277_),
    .B2(_19278_),
    .ZN(_19279_));
 OAI21_X2 _46243_ (.A(_16256_),
    .B1(_17828_),
    .B2(_17829_),
    .ZN(_19280_));
 NAND3_X2 _46244_ (.A1(_17831_),
    .A2(_17832_),
    .A3(_17236_),
    .ZN(_19281_));
 AOI21_X2 _46245_ (.A(_19000_),
    .B1(_19280_),
    .B2(_19281_),
    .ZN(_19282_));
 NOR2_X4 _46246_ (.A1(_19279_),
    .A2(_19282_),
    .ZN(_19283_));
 OAI21_X1 _46247_ (.A(_19276_),
    .B1(_19283_),
    .B2(_19224_),
    .ZN(_05090_));
 BUF_X8 _46248_ (.A(_19042_),
    .Z(_19284_));
 NAND2_X1 _46249_ (.A1(_19284_),
    .A2(\icache.lce.lce_cmd_inst.data_r [282]),
    .ZN(_19285_));
 AND3_X2 _46250_ (.A1(_17849_),
    .A2(_17459_),
    .A3(_17850_),
    .ZN(_19286_));
 AOI21_X2 _46251_ (.A(_17264_),
    .B1(_17846_),
    .B2(_17847_),
    .ZN(_19287_));
 OAI21_X2 _46252_ (.A(_18324_),
    .B1(_19286_),
    .B2(_19287_),
    .ZN(_19288_));
 OAI21_X2 _46253_ (.A(_17308_),
    .B1(_17853_),
    .B2(_17854_),
    .ZN(_19289_));
 NAND3_X2 _46254_ (.A1(_17856_),
    .A2(_17857_),
    .A3(_16230_),
    .ZN(_19290_));
 NAND3_X2 _46255_ (.A1(_19289_),
    .A2(_18747_),
    .A3(_19290_),
    .ZN(_19291_));
 NAND2_X4 _46256_ (.A1(_19288_),
    .A2(_19291_),
    .ZN(_19292_));
 OAI21_X1 _46257_ (.A(_19285_),
    .B1(_19292_),
    .B2(_19224_),
    .ZN(_05091_));
 NAND2_X1 _46258_ (.A1(_19284_),
    .A2(\icache.lce.lce_cmd_inst.data_r [283]),
    .ZN(_19293_));
 NOR3_X2 _46259_ (.A1(_17862_),
    .A2(_17863_),
    .A3(_16195_),
    .ZN(_19294_));
 AOI21_X2 _46260_ (.A(_15938_),
    .B1(_17865_),
    .B2(_17866_),
    .ZN(_19295_));
 NOR3_X2 _46261_ (.A1(_19294_),
    .A2(_19295_),
    .A3(_18132_),
    .ZN(_19296_));
 OAI21_X2 _46262_ (.A(_17308_),
    .B1(_17869_),
    .B2(_17870_),
    .ZN(_19297_));
 NAND3_X2 _46263_ (.A1(_17872_),
    .A2(_17873_),
    .A3(_16230_),
    .ZN(_19298_));
 AOI21_X2 _46264_ (.A(_19000_),
    .B1(_19297_),
    .B2(_19298_),
    .ZN(_19299_));
 NOR2_X4 _46265_ (.A1(_19296_),
    .A2(_19299_),
    .ZN(_19300_));
 OAI21_X1 _46266_ (.A(_19293_),
    .B1(_19300_),
    .B2(_19224_),
    .ZN(_05092_));
 NAND2_X1 _46267_ (.A1(_19284_),
    .A2(\icache.lce.lce_cmd_inst.data_r [284]),
    .ZN(_19301_));
 NAND2_X1 _46268_ (.A1(_17885_),
    .A2(_17228_),
    .ZN(_19302_));
 NAND2_X1 _46269_ (.A1(_17881_),
    .A2(_15567_),
    .ZN(_19303_));
 NAND2_X1 _46270_ (.A1(_19302_),
    .A2(_19303_),
    .ZN(_19304_));
 NAND2_X1 _46271_ (.A1(_19304_),
    .A2(_19034_),
    .ZN(_19305_));
 NAND2_X1 _46272_ (.A1(_17890_),
    .A2(_15343_),
    .ZN(_19306_));
 NAND3_X1 _46273_ (.A1(_17892_),
    .A2(_15395_),
    .A3(_17893_),
    .ZN(_19307_));
 NAND2_X1 _46274_ (.A1(_19306_),
    .A2(_19307_),
    .ZN(_19308_));
 NAND2_X1 _46275_ (.A1(_19308_),
    .A2(_17567_),
    .ZN(_19309_));
 NAND2_X4 _46276_ (.A1(_19305_),
    .A2(_19309_),
    .ZN(_19310_));
 BUF_X16 _46277_ (.A(_19056_),
    .Z(_19311_));
 OAI21_X1 _46278_ (.A(_19301_),
    .B1(_19310_),
    .B2(_19311_),
    .ZN(_05093_));
 NAND2_X1 _46279_ (.A1(_19284_),
    .A2(\icache.lce.lce_cmd_inst.data_r [285]),
    .ZN(_19312_));
 NOR3_X2 _46280_ (.A1(_15902_),
    .A2(_15903_),
    .A3(_16512_),
    .ZN(_19313_));
 AOI21_X1 _46281_ (.A(_17710_),
    .B1(_15907_),
    .B2(_15910_),
    .ZN(_19314_));
 OAI21_X2 _46282_ (.A(_18324_),
    .B1(_19313_),
    .B2(_19314_),
    .ZN(_19315_));
 NOR3_X4 _46283_ (.A1(_15915_),
    .A2(_15917_),
    .A3(_15779_),
    .ZN(_19316_));
 AOI21_X2 _46284_ (.A(_16227_),
    .B1(_15920_),
    .B2(_15923_),
    .ZN(_19317_));
 OAI21_X2 _46285_ (.A(_18376_),
    .B1(_19316_),
    .B2(_19317_),
    .ZN(_19318_));
 NAND2_X4 _46286_ (.A1(_19315_),
    .A2(_19318_),
    .ZN(_19319_));
 OAI21_X1 _46287_ (.A(_19312_),
    .B1(_19319_),
    .B2(_19311_),
    .ZN(_05094_));
 NAND2_X1 _46288_ (.A1(_19284_),
    .A2(\icache.lce.lce_cmd_inst.data_r [286]),
    .ZN(_19320_));
 NAND2_X1 _46289_ (.A1(_15937_),
    .A2(_17228_),
    .ZN(_19321_));
 NAND2_X1 _46290_ (.A1(_15931_),
    .A2(_15567_),
    .ZN(_19322_));
 NAND2_X1 _46291_ (.A1(_19321_),
    .A2(_19322_),
    .ZN(_19323_));
 NAND2_X1 _46292_ (.A1(_19323_),
    .A2(_19034_),
    .ZN(_19324_));
 NOR3_X2 _46293_ (.A1(_15942_),
    .A2(_15943_),
    .A3(_15779_),
    .ZN(_19325_));
 AOI21_X2 _46294_ (.A(_16227_),
    .B1(_15945_),
    .B2(_15947_),
    .ZN(_19326_));
 OAI21_X2 _46295_ (.A(_18376_),
    .B1(_19325_),
    .B2(_19326_),
    .ZN(_19327_));
 NAND2_X4 _46296_ (.A1(_19324_),
    .A2(_19327_),
    .ZN(_19328_));
 OAI21_X1 _46297_ (.A(_19320_),
    .B1(_19328_),
    .B2(_19311_),
    .ZN(_05095_));
 NAND2_X1 _46298_ (.A1(_19284_),
    .A2(\icache.lce.lce_cmd_inst.data_r [287]),
    .ZN(_19329_));
 AOI21_X2 _46299_ (.A(_18164_),
    .B1(_15953_),
    .B2(_15956_),
    .ZN(_19330_));
 AOI21_X2 _46300_ (.A(_15425_),
    .B1(_15959_),
    .B2(_15961_),
    .ZN(_19331_));
 NOR3_X2 _46301_ (.A1(_19330_),
    .A2(_19331_),
    .A3(_18132_),
    .ZN(_19332_));
 NAND2_X1 _46302_ (.A1(_15965_),
    .A2(_15909_),
    .ZN(_19333_));
 OAI211_X2 _46303_ (.A(_19333_),
    .B(_15395_),
    .C1(_18116_),
    .C2(\icache.data_mems_0__data_mem.data_o [31]),
    .ZN(_19334_));
 NAND2_X1 _46304_ (.A1(_17312_),
    .A2(_16001_),
    .ZN(_19335_));
 OAI211_X4 _46305_ (.A(_19335_),
    .B(_17981_),
    .C1(_15324_),
    .C2(\icache.data_mems_2__data_mem.data_o [31]),
    .ZN(_19336_));
 AOI21_X2 _46306_ (.A(_19000_),
    .B1(_19334_),
    .B2(_19336_),
    .ZN(_19337_));
 NOR2_X4 _46307_ (.A1(_19332_),
    .A2(_19337_),
    .ZN(_19338_));
 OAI21_X1 _46308_ (.A(_19329_),
    .B1(_19338_),
    .B2(_19311_),
    .ZN(_05096_));
 NAND2_X1 _46309_ (.A1(_19284_),
    .A2(\icache.lce.lce_cmd_inst.data_r [288]),
    .ZN(_19339_));
 NOR3_X2 _46310_ (.A1(_15974_),
    .A2(_15975_),
    .A3(_15619_),
    .ZN(_19340_));
 AOI21_X2 _46311_ (.A(_18164_),
    .B1(_15977_),
    .B2(_15979_),
    .ZN(_19341_));
 OAI21_X2 _46312_ (.A(_18324_),
    .B1(_19340_),
    .B2(_19341_),
    .ZN(_19342_));
 AOI21_X2 _46313_ (.A(_16583_),
    .B1(_15983_),
    .B2(_15987_),
    .ZN(_19343_));
 AOI21_X4 _46314_ (.A(_16227_),
    .B1(_15991_),
    .B2(_15993_),
    .ZN(_19344_));
 OAI21_X2 _46315_ (.A(_18376_),
    .B1(_19343_),
    .B2(_19344_),
    .ZN(_19345_));
 NAND2_X4 _46316_ (.A1(_19342_),
    .A2(_19345_),
    .ZN(_19346_));
 OAI21_X1 _46317_ (.A(_19339_),
    .B1(_19346_),
    .B2(_19311_),
    .ZN(_05097_));
 NAND2_X1 _46318_ (.A1(_19284_),
    .A2(\icache.lce.lce_cmd_inst.data_r [289]),
    .ZN(_19347_));
 BUF_X16 _46319_ (.A(_15819_),
    .Z(_19348_));
 OAI21_X2 _46320_ (.A(_16396_),
    .B1(_16002_),
    .B2(_16003_),
    .ZN(_19349_));
 NAND3_X2 _46321_ (.A1(_16006_),
    .A2(_16009_),
    .A3(_15446_),
    .ZN(_19350_));
 AOI21_X2 _46322_ (.A(_19348_),
    .B1(_19349_),
    .B2(_19350_),
    .ZN(_19351_));
 NAND3_X2 _46323_ (.A1(_16016_),
    .A2(_16019_),
    .A3(_15988_),
    .ZN(_19352_));
 NAND3_X4 _46324_ (.A1(_16023_),
    .A2(_16025_),
    .A3(_15464_),
    .ZN(_19353_));
 AOI21_X2 _46325_ (.A(_19005_),
    .B1(_19352_),
    .B2(_19353_),
    .ZN(_19354_));
 NOR2_X4 _46326_ (.A1(_19351_),
    .A2(_19354_),
    .ZN(_19355_));
 OAI21_X1 _46327_ (.A(_19347_),
    .B1(_19355_),
    .B2(_19311_),
    .ZN(_05098_));
 NAND2_X1 _46328_ (.A1(_19284_),
    .A2(\icache.lce.lce_cmd_inst.data_r [290]),
    .ZN(_19356_));
 OAI21_X2 _46329_ (.A(_16396_),
    .B1(_16039_),
    .B2(_16040_),
    .ZN(_19357_));
 OAI21_X2 _46330_ (.A(_15712_),
    .B1(_16043_),
    .B2(_16044_),
    .ZN(_19358_));
 AOI21_X2 _46331_ (.A(_19348_),
    .B1(_19357_),
    .B2(_19358_),
    .ZN(_19359_));
 OAI21_X2 _46332_ (.A(_16341_),
    .B1(_16030_),
    .B2(_16031_),
    .ZN(_19360_));
 NAND2_X1 _46333_ (.A1(_16036_),
    .A2(_17839_),
    .ZN(_19361_));
 OAI211_X4 _46334_ (.A(_19361_),
    .B(_15932_),
    .C1(_18116_),
    .C2(\icache.data_mems_6__data_mem.data_o [34]),
    .ZN(_19362_));
 AOI21_X2 _46335_ (.A(_19005_),
    .B1(_19360_),
    .B2(_19362_),
    .ZN(_19363_));
 NOR2_X4 _46336_ (.A1(_19359_),
    .A2(_19363_),
    .ZN(_19364_));
 OAI21_X1 _46337_ (.A(_19356_),
    .B1(_19364_),
    .B2(_19311_),
    .ZN(_05100_));
 NAND2_X1 _46338_ (.A1(_19284_),
    .A2(\icache.lce.lce_cmd_inst.data_r [291]),
    .ZN(_19365_));
 BUF_X16 _46339_ (.A(_15597_),
    .Z(_19366_));
 NOR3_X2 _46340_ (.A1(_16060_),
    .A2(_16062_),
    .A3(_15938_),
    .ZN(_19367_));
 AOI21_X2 _46341_ (.A(_17264_),
    .B1(_16065_),
    .B2(_16068_),
    .ZN(_19368_));
 OAI21_X1 _46342_ (.A(_19366_),
    .B1(_19367_),
    .B2(_19368_),
    .ZN(_19369_));
 OAI21_X2 _46343_ (.A(_15446_),
    .B1(_16051_),
    .B2(_16052_),
    .ZN(_19370_));
 NAND2_X1 _46344_ (.A1(_16057_),
    .A2(_16001_),
    .ZN(_19371_));
 OAI211_X4 _46345_ (.A(_19371_),
    .B(_15779_),
    .C1(_15324_),
    .C2(\icache.data_mems_0__data_mem.data_o [35]),
    .ZN(_19372_));
 NAND3_X2 _46346_ (.A1(_19370_),
    .A2(_19372_),
    .A3(_18460_),
    .ZN(_19373_));
 NAND2_X4 _46347_ (.A1(_19369_),
    .A2(_19373_),
    .ZN(_19374_));
 OAI21_X1 _46348_ (.A(_19365_),
    .B1(_19374_),
    .B2(_19311_),
    .ZN(_05101_));
 BUF_X8 _46349_ (.A(_19042_),
    .Z(_19375_));
 NAND2_X1 _46350_ (.A1(_19375_),
    .A2(\icache.lce.lce_cmd_inst.data_r [196]),
    .ZN(_19376_));
 AOI21_X2 _46351_ (.A(_19348_),
    .B1(_16730_),
    .B2(_16734_),
    .ZN(_19377_));
 AOI21_X1 _46352_ (.A(_19005_),
    .B1(_16739_),
    .B2(_16744_),
    .ZN(_19378_));
 NOR2_X2 _46353_ (.A1(_19377_),
    .A2(_19378_),
    .ZN(_19379_));
 OAI21_X1 _46354_ (.A(_19376_),
    .B1(_19379_),
    .B2(_19311_),
    .ZN(_04995_));
 NAND2_X1 _46355_ (.A1(_19375_),
    .A2(\icache.lce.lce_cmd_inst.data_r [197]),
    .ZN(_19380_));
 AND3_X1 _46356_ (.A1(_16750_),
    .A2(_15474_),
    .A3(_16756_),
    .ZN(_19381_));
 AOI21_X1 _46357_ (.A(_19005_),
    .B1(_16760_),
    .B2(_16764_),
    .ZN(_19382_));
 NOR2_X2 _46358_ (.A1(_19381_),
    .A2(_19382_),
    .ZN(_19383_));
 OAI21_X1 _46359_ (.A(_19380_),
    .B1(_19383_),
    .B2(_19311_),
    .ZN(_04996_));
 NAND2_X1 _46360_ (.A1(_19375_),
    .A2(\icache.lce.lce_cmd_inst.data_r [198]),
    .ZN(_19384_));
 NAND2_X2 _46361_ (.A1(_16774_),
    .A2(_18662_),
    .ZN(_19385_));
 OAI21_X1 _46362_ (.A(_19088_),
    .B1(_16778_),
    .B2(_16782_),
    .ZN(_19386_));
 NAND2_X2 _46363_ (.A1(_19385_),
    .A2(_19386_),
    .ZN(_19387_));
 BUF_X8 _46364_ (.A(_19056_),
    .Z(_19388_));
 OAI21_X1 _46365_ (.A(_19384_),
    .B1(_19387_),
    .B2(_19388_),
    .ZN(_04997_));
 NAND2_X1 _46366_ (.A1(_19375_),
    .A2(\icache.lce.lce_cmd_inst.data_r [199]),
    .ZN(_19389_));
 AOI21_X1 _46367_ (.A(_19348_),
    .B1(_16791_),
    .B2(_16795_),
    .ZN(_19390_));
 AOI21_X1 _46368_ (.A(_19005_),
    .B1(_16801_),
    .B2(_16807_),
    .ZN(_19391_));
 NOR2_X2 _46369_ (.A1(_19390_),
    .A2(_19391_),
    .ZN(_19392_));
 OAI21_X1 _46370_ (.A(_19389_),
    .B1(_19392_),
    .B2(_19388_),
    .ZN(_04998_));
 NAND2_X1 _46371_ (.A1(_19375_),
    .A2(\icache.lce.lce_cmd_inst.data_r [200]),
    .ZN(_19393_));
 OAI21_X2 _46372_ (.A(_19366_),
    .B1(_16813_),
    .B2(_16818_),
    .ZN(_19394_));
 NAND3_X2 _46373_ (.A1(_16822_),
    .A2(_18747_),
    .A3(_16827_),
    .ZN(_19395_));
 NAND2_X4 _46374_ (.A1(_19394_),
    .A2(_19395_),
    .ZN(_19396_));
 OAI21_X1 _46375_ (.A(_19393_),
    .B1(_19396_),
    .B2(_19388_),
    .ZN(_05001_));
 NAND2_X1 _46376_ (.A1(_19375_),
    .A2(\icache.lce.lce_cmd_inst.data_r [201]),
    .ZN(_19397_));
 AOI21_X2 _46377_ (.A(_19348_),
    .B1(_16834_),
    .B2(_16838_),
    .ZN(_19398_));
 BUF_X16 _46378_ (.A(_15833_),
    .Z(_19399_));
 AOI21_X2 _46379_ (.A(_19399_),
    .B1(_16844_),
    .B2(_16849_),
    .ZN(_19400_));
 NOR2_X4 _46380_ (.A1(_19398_),
    .A2(_19400_),
    .ZN(_19401_));
 OAI21_X1 _46381_ (.A(_19397_),
    .B1(_19401_),
    .B2(_19388_),
    .ZN(_05002_));
 NAND2_X1 _46382_ (.A1(_19375_),
    .A2(\icache.lce.lce_cmd_inst.data_r [202]),
    .ZN(_19402_));
 AND3_X1 _46383_ (.A1(_16857_),
    .A2(_16863_),
    .A3(_15503_),
    .ZN(_19403_));
 AOI21_X2 _46384_ (.A(_19000_),
    .B1(_16870_),
    .B2(_16874_),
    .ZN(_19404_));
 NOR2_X4 _46385_ (.A1(_19403_),
    .A2(_19404_),
    .ZN(_19405_));
 OAI21_X1 _46386_ (.A(_19402_),
    .B1(_19405_),
    .B2(_19388_),
    .ZN(_05003_));
 NAND2_X1 _46387_ (.A1(_19375_),
    .A2(\icache.lce.lce_cmd_inst.data_r [203]),
    .ZN(_19406_));
 AND3_X1 _46388_ (.A1(_16881_),
    .A2(_15474_),
    .A3(_16884_),
    .ZN(_19407_));
 AOI21_X2 _46389_ (.A(_19399_),
    .B1(_16888_),
    .B2(_16893_),
    .ZN(_19408_));
 NOR2_X4 _46390_ (.A1(_19407_),
    .A2(_19408_),
    .ZN(_19409_));
 OAI21_X1 _46391_ (.A(_19406_),
    .B1(_19409_),
    .B2(_19388_),
    .ZN(_05004_));
 NAND2_X1 _46392_ (.A1(_19375_),
    .A2(\icache.lce.lce_cmd_inst.data_r [204]),
    .ZN(_19410_));
 AOI21_X1 _46393_ (.A(_16406_),
    .B1(_16899_),
    .B2(_16902_),
    .ZN(_19411_));
 AND3_X1 _46394_ (.A1(_16906_),
    .A2(_15819_),
    .A3(_16911_),
    .ZN(_19412_));
 OR2_X4 _46395_ (.A1(_19411_),
    .A2(_19412_),
    .ZN(_19413_));
 OAI21_X1 _46396_ (.A(_19410_),
    .B1(_19413_),
    .B2(_19388_),
    .ZN(_05005_));
 NAND2_X1 _46397_ (.A1(_19375_),
    .A2(\icache.lce.lce_cmd_inst.data_r [205]),
    .ZN(_19414_));
 AOI21_X2 _46398_ (.A(_18903_),
    .B1(_16917_),
    .B2(_16922_),
    .ZN(_19415_));
 AOI21_X2 _46399_ (.A(_19000_),
    .B1(_16927_),
    .B2(_16932_),
    .ZN(_19416_));
 NOR2_X4 _46400_ (.A1(_19415_),
    .A2(_19416_),
    .ZN(_19417_));
 OAI21_X1 _46401_ (.A(_19414_),
    .B1(_19417_),
    .B2(_19388_),
    .ZN(_05006_));
 BUF_X4 _46402_ (.A(_19042_),
    .Z(_19418_));
 NAND2_X1 _46403_ (.A1(_19418_),
    .A2(\icache.lce.lce_cmd_inst.data_r [206]),
    .ZN(_19419_));
 NAND2_X1 _46404_ (.A1(_16944_),
    .A2(_19034_),
    .ZN(_19420_));
 NAND3_X2 _46405_ (.A1(_16948_),
    .A2(_18747_),
    .A3(_16952_),
    .ZN(_19421_));
 NAND2_X4 _46406_ (.A1(_19420_),
    .A2(_19421_),
    .ZN(_19422_));
 OAI21_X1 _46407_ (.A(_19419_),
    .B1(_19422_),
    .B2(_19388_),
    .ZN(_05007_));
 NAND2_X1 _46408_ (.A1(_19418_),
    .A2(\icache.lce.lce_cmd_inst.data_r [207]),
    .ZN(_19423_));
 AOI21_X2 _46409_ (.A(_18903_),
    .B1(_16960_),
    .B2(_16964_),
    .ZN(_19424_));
 BUF_X16 _46410_ (.A(_15367_),
    .Z(_19425_));
 AOI21_X2 _46411_ (.A(_19425_),
    .B1(_16969_),
    .B2(_16974_),
    .ZN(_19426_));
 NOR2_X4 _46412_ (.A1(_19424_),
    .A2(_19426_),
    .ZN(_19427_));
 OAI21_X1 _46413_ (.A(_19423_),
    .B1(_19427_),
    .B2(_19388_),
    .ZN(_05008_));
 NAND2_X1 _46414_ (.A1(_19418_),
    .A2(\icache.lce.lce_cmd_inst.data_r [208]),
    .ZN(_19428_));
 AOI21_X1 _46415_ (.A(_19348_),
    .B1(_16980_),
    .B2(_16985_),
    .ZN(_19429_));
 AOI21_X1 _46416_ (.A(_19399_),
    .B1(_16990_),
    .B2(_16994_),
    .ZN(_19430_));
 NOR2_X2 _46417_ (.A1(_19429_),
    .A2(_19430_),
    .ZN(_19431_));
 BUF_X4 _46418_ (.A(_19056_),
    .Z(_19432_));
 OAI21_X1 _46419_ (.A(_19428_),
    .B1(_19431_),
    .B2(_19432_),
    .ZN(_05009_));
 NAND2_X1 _46420_ (.A1(_19418_),
    .A2(\icache.lce.lce_cmd_inst.data_r [209]),
    .ZN(_19433_));
 NAND2_X1 _46421_ (.A1(_17010_),
    .A2(_19034_),
    .ZN(_19434_));
 OAI21_X2 _46422_ (.A(_18376_),
    .B1(_17015_),
    .B2(_17020_),
    .ZN(_19435_));
 NAND2_X2 _46423_ (.A1(_19434_),
    .A2(_19435_),
    .ZN(_19436_));
 OAI21_X1 _46424_ (.A(_19433_),
    .B1(_19436_),
    .B2(_19432_),
    .ZN(_05010_));
 NAND2_X1 _46425_ (.A1(_19418_),
    .A2(\icache.lce.lce_cmd_inst.data_r [210]),
    .ZN(_19437_));
 AOI21_X1 _46426_ (.A(_19348_),
    .B1(_17026_),
    .B2(_17031_),
    .ZN(_19438_));
 AOI21_X1 _46427_ (.A(_19399_),
    .B1(_17036_),
    .B2(_17041_),
    .ZN(_19439_));
 NOR2_X2 _46428_ (.A1(_19438_),
    .A2(_19439_),
    .ZN(_19440_));
 OAI21_X1 _46429_ (.A(_19437_),
    .B1(_19440_),
    .B2(_19432_),
    .ZN(_05012_));
 NAND2_X1 _46430_ (.A1(_19418_),
    .A2(\icache.lce.lce_cmd_inst.data_r [211]),
    .ZN(_19441_));
 AOI21_X1 _46431_ (.A(_18903_),
    .B1(_17047_),
    .B2(_17051_),
    .ZN(_19442_));
 AOI21_X2 _46432_ (.A(_19425_),
    .B1(_17057_),
    .B2(_17062_),
    .ZN(_19443_));
 NOR2_X2 _46433_ (.A1(_19442_),
    .A2(_19443_),
    .ZN(_19444_));
 OAI21_X1 _46434_ (.A(_19441_),
    .B1(_19444_),
    .B2(_19432_),
    .ZN(_05013_));
 NAND2_X1 _46435_ (.A1(_19418_),
    .A2(\icache.lce.lce_cmd_inst.data_r [212]),
    .ZN(_19445_));
 NAND3_X1 _46436_ (.A1(_17069_),
    .A2(_16360_),
    .A3(_17072_),
    .ZN(_19446_));
 NAND3_X1 _46437_ (.A1(_17078_),
    .A2(_17084_),
    .A3(_15315_),
    .ZN(_19447_));
 AND2_X4 _46438_ (.A1(_19446_),
    .A2(_19447_),
    .ZN(_19448_));
 OAI21_X1 _46439_ (.A(_19445_),
    .B1(_19448_),
    .B2(_19432_),
    .ZN(_05014_));
 NAND2_X1 _46440_ (.A1(_19418_),
    .A2(\icache.lce.lce_cmd_inst.data_r [213]),
    .ZN(_19449_));
 NAND2_X1 _46441_ (.A1(_17097_),
    .A2(_18662_),
    .ZN(_19450_));
 NAND3_X1 _46442_ (.A1(_17101_),
    .A2(_18918_),
    .A3(_17105_),
    .ZN(_19451_));
 NAND2_X2 _46443_ (.A1(_19450_),
    .A2(_19451_),
    .ZN(_19452_));
 OAI21_X1 _46444_ (.A(_19449_),
    .B1(_19452_),
    .B2(_19432_),
    .ZN(_05015_));
 NAND2_X1 _46445_ (.A1(_19418_),
    .A2(\icache.lce.lce_cmd_inst.data_r [214]),
    .ZN(_19453_));
 AOI21_X1 _46446_ (.A(_18903_),
    .B1(_17111_),
    .B2(_17114_),
    .ZN(_19454_));
 AOI21_X1 _46447_ (.A(_19425_),
    .B1(_17119_),
    .B2(_17123_),
    .ZN(_19455_));
 NOR2_X2 _46448_ (.A1(_19454_),
    .A2(_19455_),
    .ZN(_19456_));
 OAI21_X1 _46449_ (.A(_19453_),
    .B1(_19456_),
    .B2(_19432_),
    .ZN(_05016_));
 NAND2_X1 _46450_ (.A1(_19418_),
    .A2(\icache.lce.lce_cmd_inst.data_r [193]),
    .ZN(_19457_));
 AND3_X1 _46451_ (.A1(_16670_),
    .A2(_15621_),
    .A3(_16673_),
    .ZN(_19458_));
 AOI21_X2 _46452_ (.A(_19399_),
    .B1(_16677_),
    .B2(_16681_),
    .ZN(_19459_));
 NOR2_X4 _46453_ (.A1(_19458_),
    .A2(_19459_),
    .ZN(_19460_));
 OAI21_X1 _46454_ (.A(_19457_),
    .B1(_19460_),
    .B2(_19432_),
    .ZN(_04992_));
 BUF_X16 _46455_ (.A(_19042_),
    .Z(_19461_));
 NAND2_X1 _46456_ (.A1(_19461_),
    .A2(\icache.lce.lce_cmd_inst.data_r [194]),
    .ZN(_19462_));
 AOI21_X2 _46457_ (.A(_18351_),
    .B1(_16688_),
    .B2(_16691_),
    .ZN(_19463_));
 AND3_X1 _46458_ (.A1(_16696_),
    .A2(_15430_),
    .A3(_16700_),
    .ZN(_19464_));
 OR2_X4 _46459_ (.A1(_19463_),
    .A2(_19464_),
    .ZN(_19465_));
 OAI21_X1 _46460_ (.A(_19462_),
    .B1(_19465_),
    .B2(_19432_),
    .ZN(_04993_));
 NAND2_X1 _46461_ (.A1(_19461_),
    .A2(\icache.lce.lce_cmd_inst.data_r [195]),
    .ZN(_19466_));
 AOI21_X1 _46462_ (.A(_16406_),
    .B1(_16707_),
    .B2(_16712_),
    .ZN(_19467_));
 AND3_X1 _46463_ (.A1(_16717_),
    .A2(_16721_),
    .A3(_15819_),
    .ZN(_19468_));
 OR2_X4 _46464_ (.A1(_19467_),
    .A2(_19468_),
    .ZN(_19469_));
 OAI21_X1 _46465_ (.A(_19466_),
    .B1(_19469_),
    .B2(_19432_),
    .ZN(_04994_));
 NAND2_X1 _46466_ (.A1(_19461_),
    .A2(\icache.lce.lce_cmd_inst.data_r [116]),
    .ZN(_19470_));
 AOI21_X1 _46467_ (.A(_16406_),
    .B1(_18474_),
    .B2(_18475_),
    .ZN(_19471_));
 AND3_X1 _46468_ (.A1(_18478_),
    .A2(_18480_),
    .A3(_15819_),
    .ZN(_19472_));
 OR2_X2 _46469_ (.A1(_19471_),
    .A2(_19472_),
    .ZN(_19473_));
 BUF_X8 _46470_ (.A(_19056_),
    .Z(_19474_));
 OAI21_X1 _46471_ (.A(_19470_),
    .B1(_19473_),
    .B2(_19474_),
    .ZN(_04907_));
 NAND2_X1 _46472_ (.A1(_19461_),
    .A2(\icache.lce.lce_cmd_inst.data_r [117]),
    .ZN(_19475_));
 OAI21_X2 _46473_ (.A(_17827_),
    .B1(_18485_),
    .B2(_18486_),
    .ZN(_19476_));
 NAND3_X2 _46474_ (.A1(_18488_),
    .A2(_18918_),
    .A3(_18489_),
    .ZN(_19477_));
 NAND2_X4 _46475_ (.A1(_19476_),
    .A2(_19477_),
    .ZN(_19478_));
 OAI21_X1 _46476_ (.A(_19475_),
    .B1(_19478_),
    .B2(_19474_),
    .ZN(_04908_));
 NAND2_X1 _46477_ (.A1(_19461_),
    .A2(\icache.lce.lce_cmd_inst.data_r [118]),
    .ZN(_19479_));
 AND3_X1 _46478_ (.A1(_18493_),
    .A2(_18494_),
    .A3(_16562_),
    .ZN(_19480_));
 AOI21_X1 _46479_ (.A(_19399_),
    .B1(_18496_),
    .B2(_18497_),
    .ZN(_19481_));
 NOR2_X2 _46480_ (.A1(_19480_),
    .A2(_19481_),
    .ZN(_19482_));
 OAI21_X1 _46481_ (.A(_19479_),
    .B1(_19482_),
    .B2(_19474_),
    .ZN(_04909_));
 NAND2_X1 _46482_ (.A1(_19461_),
    .A2(\icache.lce.lce_cmd_inst.data_r [119]),
    .ZN(_19483_));
 NAND2_X2 _46483_ (.A1(_18503_),
    .A2(_19034_),
    .ZN(_19484_));
 OAI21_X2 _46484_ (.A(_18376_),
    .B1(_18505_),
    .B2(_18506_),
    .ZN(_19485_));
 NAND2_X4 _46485_ (.A1(_19484_),
    .A2(_19485_),
    .ZN(_19486_));
 OAI21_X1 _46486_ (.A(_19483_),
    .B1(_19486_),
    .B2(_19474_),
    .ZN(_04910_));
 NAND2_X1 _46487_ (.A1(_19461_),
    .A2(\icache.lce.lce_cmd_inst.data_r [120]),
    .ZN(_19487_));
 NAND2_X1 _46488_ (.A1(_18512_),
    .A2(_19034_),
    .ZN(_19488_));
 NAND2_X1 _46489_ (.A1(_18516_),
    .A2(_17567_),
    .ZN(_19489_));
 NAND2_X2 _46490_ (.A1(_19488_),
    .A2(_19489_),
    .ZN(_19490_));
 OAI21_X1 _46491_ (.A(_19487_),
    .B1(_19490_),
    .B2(_19474_),
    .ZN(_04912_));
 NAND2_X1 _46492_ (.A1(_19461_),
    .A2(\icache.lce.lce_cmd_inst.data_r [121]),
    .ZN(_19491_));
 NOR3_X2 _46493_ (.A1(_18520_),
    .A2(_18521_),
    .A3(_18085_),
    .ZN(_19492_));
 AOI21_X2 _46494_ (.A(_19399_),
    .B1(_18523_),
    .B2(_18524_),
    .ZN(_19493_));
 NOR2_X4 _46495_ (.A1(_19492_),
    .A2(_19493_),
    .ZN(_19494_));
 OAI21_X1 _46496_ (.A(_19491_),
    .B1(_19494_),
    .B2(_19474_),
    .ZN(_04913_));
 NAND2_X1 _46497_ (.A1(_19461_),
    .A2(\icache.lce.lce_cmd_inst.data_r [122]),
    .ZN(_19495_));
 AND3_X1 _46498_ (.A1(_18528_),
    .A2(_18529_),
    .A3(_16562_),
    .ZN(_19496_));
 AOI21_X4 _46499_ (.A(_19399_),
    .B1(_18532_),
    .B2(_18533_),
    .ZN(_19497_));
 NOR2_X4 _46500_ (.A1(_19496_),
    .A2(_19497_),
    .ZN(_19498_));
 OAI21_X1 _46501_ (.A(_19495_),
    .B1(_19498_),
    .B2(_19474_),
    .ZN(_04914_));
 NAND2_X1 _46502_ (.A1(_19461_),
    .A2(\icache.lce.lce_cmd_inst.data_r [123]),
    .ZN(_19499_));
 AND3_X1 _46503_ (.A1(_18537_),
    .A2(_18538_),
    .A3(_16562_),
    .ZN(_19500_));
 AOI21_X2 _46504_ (.A(_19399_),
    .B1(_18540_),
    .B2(_18541_),
    .ZN(_19501_));
 NOR2_X4 _46505_ (.A1(_19500_),
    .A2(_19501_),
    .ZN(_19502_));
 OAI21_X1 _46506_ (.A(_19499_),
    .B1(_19502_),
    .B2(_19474_),
    .ZN(_04915_));
 BUF_X8 _46507_ (.A(_19042_),
    .Z(_19503_));
 NAND2_X1 _46508_ (.A1(_19503_),
    .A2(\icache.lce.lce_cmd_inst.data_r [124]),
    .ZN(_19504_));
 BUF_X16 _46509_ (.A(_15328_),
    .Z(_19505_));
 AOI21_X1 _46510_ (.A(_19505_),
    .B1(_18546_),
    .B2(_18548_),
    .ZN(_19506_));
 AOI21_X1 _46511_ (.A(_19425_),
    .B1(_18550_),
    .B2(_18551_),
    .ZN(_19507_));
 NOR2_X2 _46512_ (.A1(_19506_),
    .A2(_19507_),
    .ZN(_19508_));
 OAI21_X1 _46513_ (.A(_19504_),
    .B1(_19508_),
    .B2(_19474_),
    .ZN(_04916_));
 NAND2_X1 _46514_ (.A1(_19503_),
    .A2(\icache.lce.lce_cmd_inst.data_r [125]),
    .ZN(_19509_));
 BUF_X16 _46515_ (.A(_15734_),
    .Z(_19510_));
 OAI21_X1 _46516_ (.A(_19510_),
    .B1(_18555_),
    .B2(_18556_),
    .ZN(_19511_));
 NAND3_X2 _46517_ (.A1(_18558_),
    .A2(_18918_),
    .A3(_18559_),
    .ZN(_19512_));
 NAND2_X4 _46518_ (.A1(_19511_),
    .A2(_19512_),
    .ZN(_19513_));
 OAI21_X1 _46519_ (.A(_19509_),
    .B1(_19513_),
    .B2(_19474_),
    .ZN(_04917_));
 NAND2_X1 _46520_ (.A1(_19503_),
    .A2(\icache.lce.lce_cmd_inst.data_r [126]),
    .ZN(_19514_));
 NAND2_X1 _46521_ (.A1(_18569_),
    .A2(_18662_),
    .ZN(_19515_));
 NAND2_X1 _46522_ (.A1(_18565_),
    .A2(_15598_),
    .ZN(_19516_));
 NAND2_X2 _46523_ (.A1(_19515_),
    .A2(_19516_),
    .ZN(_19517_));
 BUF_X16 _46524_ (.A(_19056_),
    .Z(_19518_));
 OAI21_X1 _46525_ (.A(_19514_),
    .B1(_19517_),
    .B2(_19518_),
    .ZN(_04918_));
 NAND2_X1 _46526_ (.A1(_19503_),
    .A2(\icache.lce.lce_cmd_inst.data_r [127]),
    .ZN(_19519_));
 AND3_X1 _46527_ (.A1(_18574_),
    .A2(_18575_),
    .A3(_16562_),
    .ZN(_19520_));
 AOI21_X2 _46528_ (.A(_19399_),
    .B1(_18577_),
    .B2(_18578_),
    .ZN(_19521_));
 NOR2_X4 _46529_ (.A1(_19520_),
    .A2(_19521_),
    .ZN(_19522_));
 OAI21_X1 _46530_ (.A(_19519_),
    .B1(_19522_),
    .B2(_19518_),
    .ZN(_04919_));
 NAND2_X1 _46531_ (.A1(_19503_),
    .A2(\icache.lce.lce_cmd_inst.data_r [128]),
    .ZN(_19523_));
 AOI21_X2 _46532_ (.A(_19348_),
    .B1(_18582_),
    .B2(_18584_),
    .ZN(_19524_));
 BUF_X16 _46533_ (.A(_15833_),
    .Z(_19525_));
 AOI21_X2 _46534_ (.A(_19525_),
    .B1(_18586_),
    .B2(_18587_),
    .ZN(_19526_));
 NOR2_X4 _46535_ (.A1(_19524_),
    .A2(_19526_),
    .ZN(_19527_));
 OAI21_X1 _46536_ (.A(_19523_),
    .B1(_19527_),
    .B2(_19518_),
    .ZN(_04920_));
 NAND2_X1 _46537_ (.A1(_19503_),
    .A2(\icache.lce.lce_cmd_inst.data_r [129]),
    .ZN(_19528_));
 AOI21_X1 _46538_ (.A(_16406_),
    .B1(_18594_),
    .B2(_18598_),
    .ZN(_19529_));
 NOR3_X1 _46539_ (.A1(_18602_),
    .A2(_18605_),
    .A3(_15734_),
    .ZN(_19530_));
 OR2_X4 _46540_ (.A1(_19529_),
    .A2(_19530_),
    .ZN(_19531_));
 OAI21_X1 _46541_ (.A(_19528_),
    .B1(_19531_),
    .B2(_19518_),
    .ZN(_04921_));
 NAND2_X1 _46542_ (.A1(_19503_),
    .A2(\icache.lce.lce_cmd_inst.data_r [130]),
    .ZN(_19532_));
 AOI21_X2 _46543_ (.A(_19505_),
    .B1(_18618_),
    .B2(_18621_),
    .ZN(_19533_));
 AOI21_X2 _46544_ (.A(_19425_),
    .B1(_18611_),
    .B2(_18614_),
    .ZN(_19534_));
 NOR2_X4 _46545_ (.A1(_19533_),
    .A2(_19534_),
    .ZN(_19535_));
 OAI21_X1 _46546_ (.A(_19532_),
    .B1(_19535_),
    .B2(_19518_),
    .ZN(_04923_));
 NAND2_X1 _46547_ (.A1(_19503_),
    .A2(\icache.lce.lce_cmd_inst.data_r [131]),
    .ZN(_19536_));
 AND3_X1 _46548_ (.A1(_18633_),
    .A2(_18805_),
    .A3(_18636_),
    .ZN(_19537_));
 AOI21_X2 _46549_ (.A(_19425_),
    .B1(_18627_),
    .B2(_18630_),
    .ZN(_19538_));
 NOR2_X4 _46550_ (.A1(_19537_),
    .A2(_19538_),
    .ZN(_19539_));
 OAI21_X1 _46551_ (.A(_19536_),
    .B1(_19539_),
    .B2(_19518_),
    .ZN(_04924_));
 NAND2_X1 _46552_ (.A1(_19503_),
    .A2(\icache.lce.lce_cmd_inst.data_r [132]),
    .ZN(_19540_));
 AND3_X1 _46553_ (.A1(_18642_),
    .A2(_15621_),
    .A3(_18644_),
    .ZN(_19541_));
 AOI21_X2 _46554_ (.A(_19525_),
    .B1(_18648_),
    .B2(_18651_),
    .ZN(_19542_));
 NOR2_X4 _46555_ (.A1(_19541_),
    .A2(_19542_),
    .ZN(_19543_));
 OAI21_X1 _46556_ (.A(_19540_),
    .B1(_19543_),
    .B2(_19518_),
    .ZN(_04925_));
 NAND2_X1 _46557_ (.A1(_19503_),
    .A2(\icache.lce.lce_cmd_inst.data_r [133]),
    .ZN(_19544_));
 NAND2_X1 _46558_ (.A1(_18661_),
    .A2(_19034_),
    .ZN(_19545_));
 OAI21_X2 _46559_ (.A(_18376_),
    .B1(_18666_),
    .B2(_18669_),
    .ZN(_19546_));
 NAND2_X4 _46560_ (.A1(_19545_),
    .A2(_19546_),
    .ZN(_19547_));
 OAI21_X1 _46561_ (.A(_19544_),
    .B1(_19547_),
    .B2(_19518_),
    .ZN(_04926_));
 BUF_X4 _46562_ (.A(_19042_),
    .Z(_19548_));
 NAND2_X1 _46563_ (.A1(_19548_),
    .A2(\icache.lce.lce_cmd_inst.data_r [134]),
    .ZN(_19549_));
 OAI21_X1 _46564_ (.A(_19179_),
    .B1(_18677_),
    .B2(_18680_),
    .ZN(_19550_));
 OAI21_X1 _46565_ (.A(_19183_),
    .B1(_18684_),
    .B2(_18687_),
    .ZN(_19551_));
 AND2_X4 _46566_ (.A1(_19550_),
    .A2(_19551_),
    .ZN(_19552_));
 OAI21_X1 _46567_ (.A(_19549_),
    .B1(_19552_),
    .B2(_19518_),
    .ZN(_04927_));
 NAND2_X1 _46568_ (.A1(_19548_),
    .A2(\icache.lce.lce_cmd_inst.data_r [135]),
    .ZN(_19553_));
 AND3_X1 _46569_ (.A1(_17900_),
    .A2(_15621_),
    .A3(_17904_),
    .ZN(_19554_));
 AOI21_X2 _46570_ (.A(_19525_),
    .B1(_17908_),
    .B2(_17911_),
    .ZN(_19555_));
 NOR2_X4 _46571_ (.A1(_19554_),
    .A2(_19555_),
    .ZN(_19556_));
 OAI21_X1 _46572_ (.A(_19553_),
    .B1(_19556_),
    .B2(_19518_),
    .ZN(_04928_));
 NAND2_X1 _46573_ (.A1(_19548_),
    .A2(\icache.lce.lce_cmd_inst.data_r [136]),
    .ZN(_19557_));
 OAI21_X1 _46574_ (.A(_18922_),
    .B1(_17918_),
    .B2(_17921_),
    .ZN(_19558_));
 OAI21_X2 _46575_ (.A(_18366_),
    .B1(_17925_),
    .B2(_17928_),
    .ZN(_19559_));
 AND2_X4 _46576_ (.A1(_19558_),
    .A2(_19559_),
    .ZN(_19560_));
 BUF_X4 _46577_ (.A(_19056_),
    .Z(_19561_));
 OAI21_X1 _46578_ (.A(_19557_),
    .B1(_19560_),
    .B2(_19561_),
    .ZN(_04929_));
 NAND2_X1 _46579_ (.A1(_19548_),
    .A2(\icache.lce.lce_cmd_inst.data_r [137]),
    .ZN(_19562_));
 OAI21_X1 _46580_ (.A(_19510_),
    .B1(_17935_),
    .B2(_17938_),
    .ZN(_19563_));
 OAI21_X2 _46581_ (.A(_19088_),
    .B1(_17942_),
    .B2(_17945_),
    .ZN(_19564_));
 NAND2_X4 _46582_ (.A1(_19563_),
    .A2(_19564_),
    .ZN(_19565_));
 OAI21_X1 _46583_ (.A(_19562_),
    .B1(_19565_),
    .B2(_19561_),
    .ZN(_04930_));
 NAND2_X1 _46584_ (.A1(_19548_),
    .A2(\icache.lce.lce_cmd_inst.data_r [138]),
    .ZN(_19566_));
 AOI21_X2 _46585_ (.A(_19505_),
    .B1(_17566_),
    .B2(_17570_),
    .ZN(_19567_));
 AOI21_X2 _46586_ (.A(_19425_),
    .B1(_17574_),
    .B2(_17577_),
    .ZN(_19568_));
 NOR2_X4 _46587_ (.A1(_19567_),
    .A2(_19568_),
    .ZN(_19569_));
 OAI21_X1 _46588_ (.A(_19566_),
    .B1(_19569_),
    .B2(_19561_),
    .ZN(_04931_));
 NAND2_X1 _46589_ (.A1(_19548_),
    .A2(\icache.lce.lce_cmd_inst.data_r [139]),
    .ZN(_19570_));
 OAI21_X2 _46590_ (.A(_19510_),
    .B1(_17585_),
    .B2(_17589_),
    .ZN(_19571_));
 OAI21_X2 _46591_ (.A(_19088_),
    .B1(_17593_),
    .B2(_17596_),
    .ZN(_19572_));
 NAND2_X4 _46592_ (.A1(_19571_),
    .A2(_19572_),
    .ZN(_19573_));
 OAI21_X1 _46593_ (.A(_19570_),
    .B1(_19573_),
    .B2(_19561_),
    .ZN(_04932_));
 NAND2_X1 _46594_ (.A1(_19548_),
    .A2(\icache.lce.lce_cmd_inst.data_r [140]),
    .ZN(_19574_));
 NAND3_X1 _46595_ (.A1(_17602_),
    .A2(_16438_),
    .A3(_17605_),
    .ZN(_19575_));
 OAI21_X1 _46596_ (.A(_18366_),
    .B1(_17609_),
    .B2(_17612_),
    .ZN(_19576_));
 AND2_X4 _46597_ (.A1(_19575_),
    .A2(_19576_),
    .ZN(_19577_));
 OAI21_X1 _46598_ (.A(_19574_),
    .B1(_19577_),
    .B2(_19561_),
    .ZN(_04934_));
 NAND2_X1 _46599_ (.A1(_19548_),
    .A2(\icache.lce.lce_cmd_inst.data_r [141]),
    .ZN(_19578_));
 BUF_X16 _46600_ (.A(_15579_),
    .Z(_19579_));
 NAND2_X1 _46601_ (.A1(_17624_),
    .A2(_19579_),
    .ZN(_19580_));
 NAND2_X1 _46602_ (.A1(_17633_),
    .A2(_15598_),
    .ZN(_19581_));
 NAND2_X4 _46603_ (.A1(_19580_),
    .A2(_19581_),
    .ZN(_19582_));
 OAI21_X1 _46604_ (.A(_19578_),
    .B1(_19582_),
    .B2(_19561_),
    .ZN(_04935_));
 NAND2_X1 _46605_ (.A1(_19548_),
    .A2(\icache.lce.lce_cmd_inst.data_r [142]),
    .ZN(_19583_));
 OAI21_X1 _46606_ (.A(_18922_),
    .B1(_17641_),
    .B2(_17644_),
    .ZN(_19584_));
 NAND3_X1 _46607_ (.A1(_17647_),
    .A2(_17415_),
    .A3(_17650_),
    .ZN(_19585_));
 AND2_X4 _46608_ (.A1(_19584_),
    .A2(_19585_),
    .ZN(_19586_));
 OAI21_X1 _46609_ (.A(_19583_),
    .B1(_19586_),
    .B2(_19561_),
    .ZN(_04936_));
 NAND2_X1 _46610_ (.A1(_19548_),
    .A2(\icache.lce.lce_cmd_inst.data_r [143]),
    .ZN(_19587_));
 OAI21_X2 _46611_ (.A(_19366_),
    .B1(_17656_),
    .B2(_17659_),
    .ZN(_19588_));
 NAND3_X2 _46612_ (.A1(_17663_),
    .A2(_17666_),
    .A3(_18460_),
    .ZN(_19589_));
 NAND2_X4 _46613_ (.A1(_19588_),
    .A2(_19589_),
    .ZN(_19590_));
 OAI21_X1 _46614_ (.A(_19587_),
    .B1(_19590_),
    .B2(_19561_),
    .ZN(_04937_));
 BUF_X4 _46615_ (.A(_19042_),
    .Z(_19591_));
 NAND2_X1 _46616_ (.A1(_19591_),
    .A2(\icache.lce.lce_cmd_inst.data_r [144]),
    .ZN(_19592_));
 BUF_X16 _46617_ (.A(_15670_),
    .Z(_19593_));
 NAND2_X1 _46618_ (.A1(_17677_),
    .A2(_19593_),
    .ZN(_19594_));
 BUF_X16 _46619_ (.A(_15644_),
    .Z(_19595_));
 OAI21_X2 _46620_ (.A(_19595_),
    .B1(_17681_),
    .B2(_17684_),
    .ZN(_19596_));
 NAND2_X4 _46621_ (.A1(_19594_),
    .A2(_19596_),
    .ZN(_19597_));
 OAI21_X1 _46622_ (.A(_19592_),
    .B1(_19597_),
    .B2(_19561_),
    .ZN(_04938_));
 NAND2_X1 _46623_ (.A1(_19591_),
    .A2(\icache.lce.lce_cmd_inst.data_r [145]),
    .ZN(_19598_));
 NAND2_X1 _46624_ (.A1(_17695_),
    .A2(_19593_),
    .ZN(_19599_));
 OAI21_X2 _46625_ (.A(_19595_),
    .B1(_17699_),
    .B2(_17702_),
    .ZN(_19600_));
 NAND2_X4 _46626_ (.A1(_19599_),
    .A2(_19600_),
    .ZN(_19601_));
 OAI21_X1 _46627_ (.A(_19598_),
    .B1(_19601_),
    .B2(_19561_),
    .ZN(_04939_));
 NAND2_X1 _46628_ (.A1(_19591_),
    .A2(\icache.lce.lce_cmd_inst.data_r [146]),
    .ZN(_19602_));
 OAI21_X2 _46629_ (.A(_19366_),
    .B1(_17709_),
    .B2(_17713_),
    .ZN(_19603_));
 OAI21_X2 _46630_ (.A(_19595_),
    .B1(_17717_),
    .B2(_17720_),
    .ZN(_19604_));
 NAND2_X4 _46631_ (.A1(_19603_),
    .A2(_19604_),
    .ZN(_19605_));
 BUF_X4 _46632_ (.A(_19056_),
    .Z(_19606_));
 OAI21_X1 _46633_ (.A(_19602_),
    .B1(_19605_),
    .B2(_19606_),
    .ZN(_04940_));
 NAND2_X1 _46634_ (.A1(_19591_),
    .A2(\icache.lce.lce_cmd_inst.data_r [147]),
    .ZN(_19607_));
 NAND2_X1 _46635_ (.A1(_17730_),
    .A2(_19593_),
    .ZN(_19608_));
 OAI21_X2 _46636_ (.A(_19595_),
    .B1(_17735_),
    .B2(_17738_),
    .ZN(_19609_));
 NAND2_X4 _46637_ (.A1(_19608_),
    .A2(_19609_),
    .ZN(_19610_));
 OAI21_X1 _46638_ (.A(_19607_),
    .B1(_19610_),
    .B2(_19606_),
    .ZN(_04941_));
 NAND2_X1 _46639_ (.A1(_19591_),
    .A2(\icache.lce.lce_cmd_inst.data_r [148]),
    .ZN(_19611_));
 OAI21_X1 _46640_ (.A(_19179_),
    .B1(_17745_),
    .B2(_17748_),
    .ZN(_19612_));
 NAND3_X1 _46641_ (.A1(_17752_),
    .A2(_16372_),
    .A3(_17754_),
    .ZN(_19613_));
 AND2_X4 _46642_ (.A1(_19612_),
    .A2(_19613_),
    .ZN(_19614_));
 OAI21_X1 _46643_ (.A(_19611_),
    .B1(_19614_),
    .B2(_19606_),
    .ZN(_04942_));
 NAND2_X1 _46644_ (.A1(_19591_),
    .A2(\icache.lce.lce_cmd_inst.data_r [149]),
    .ZN(_19615_));
 NOR3_X1 _46645_ (.A1(_17760_),
    .A2(_15724_),
    .A3(_17763_),
    .ZN(_19616_));
 AOI21_X2 _46646_ (.A(_18419_),
    .B1(_17767_),
    .B2(_17769_),
    .ZN(_19617_));
 OR2_X4 _46647_ (.A1(_19616_),
    .A2(_19617_),
    .ZN(_19618_));
 OAI21_X1 _46648_ (.A(_19615_),
    .B1(_19618_),
    .B2(_19606_),
    .ZN(_04943_));
 NAND2_X1 _46649_ (.A1(_19591_),
    .A2(\icache.lce.lce_cmd_inst.data_r [150]),
    .ZN(_19619_));
 NAND2_X1 _46650_ (.A1(_17781_),
    .A2(_19579_),
    .ZN(_19620_));
 NAND2_X1 _46651_ (.A1(_17789_),
    .A2(_15905_),
    .ZN(_19621_));
 NAND2_X4 _46652_ (.A1(_19620_),
    .A2(_19621_),
    .ZN(_19622_));
 OAI21_X1 _46653_ (.A(_19619_),
    .B1(_19622_),
    .B2(_19606_),
    .ZN(_04945_));
 NAND2_X1 _46654_ (.A1(_19591_),
    .A2(\icache.lce.lce_cmd_inst.data_r [151]),
    .ZN(_19623_));
 NOR2_X1 _46655_ (.A1(_17799_),
    .A2(_16200_),
    .ZN(_19624_));
 AOI21_X2 _46656_ (.A(_19525_),
    .B1(_17803_),
    .B2(_17806_),
    .ZN(_19625_));
 NOR2_X4 _46657_ (.A1(_19624_),
    .A2(_19625_),
    .ZN(_19626_));
 OAI21_X1 _46658_ (.A(_19623_),
    .B1(_19626_),
    .B2(_19606_),
    .ZN(_04946_));
 NAND2_X1 _46659_ (.A1(_19591_),
    .A2(\icache.lce.lce_cmd_inst.data_r [152]),
    .ZN(_19627_));
 AOI21_X2 _46660_ (.A(_19348_),
    .B1(_17812_),
    .B2(_17815_),
    .ZN(_19628_));
 AOI21_X2 _46661_ (.A(_19525_),
    .B1(_17820_),
    .B2(_17823_),
    .ZN(_19629_));
 NOR2_X4 _46662_ (.A1(_19628_),
    .A2(_19629_),
    .ZN(_19630_));
 OAI21_X1 _46663_ (.A(_19627_),
    .B1(_19630_),
    .B2(_19606_),
    .ZN(_04947_));
 NAND2_X1 _46664_ (.A1(_19591_),
    .A2(\icache.lce.lce_cmd_inst.data_r [153]),
    .ZN(_19631_));
 OAI21_X1 _46665_ (.A(_19510_),
    .B1(_17837_),
    .B2(_17841_),
    .ZN(_19632_));
 OAI21_X2 _46666_ (.A(_19088_),
    .B1(_17830_),
    .B2(_17833_),
    .ZN(_19633_));
 NAND2_X4 _46667_ (.A1(_19632_),
    .A2(_19633_),
    .ZN(_19634_));
 OAI21_X1 _46668_ (.A(_19631_),
    .B1(_19634_),
    .B2(_19606_),
    .ZN(_04948_));
 BUF_X8 _46669_ (.A(_15301_),
    .Z(_19635_));
 BUF_X4 _46670_ (.A(_19635_),
    .Z(_19636_));
 NAND2_X1 _46671_ (.A1(_19636_),
    .A2(\icache.lce.lce_cmd_inst.data_r [154]),
    .ZN(_19637_));
 OR3_X2 _46672_ (.A1(_17848_),
    .A2(_17851_),
    .A3(_15655_),
    .ZN(_19638_));
 NAND3_X2 _46673_ (.A1(_17855_),
    .A2(_18918_),
    .A3(_17858_),
    .ZN(_19639_));
 NAND2_X4 _46674_ (.A1(_19638_),
    .A2(_19639_),
    .ZN(_19640_));
 OAI21_X1 _46675_ (.A(_19637_),
    .B1(_19640_),
    .B2(_19606_),
    .ZN(_04949_));
 NAND2_X1 _46676_ (.A1(_19636_),
    .A2(\icache.lce.lce_cmd_inst.data_r [155]),
    .ZN(_19641_));
 AOI21_X2 _46677_ (.A(_19505_),
    .B1(_17871_),
    .B2(_17874_),
    .ZN(_19642_));
 AOI21_X2 _46678_ (.A(_19425_),
    .B1(_17864_),
    .B2(_17867_),
    .ZN(_19643_));
 NOR2_X4 _46679_ (.A1(_19642_),
    .A2(_19643_),
    .ZN(_19644_));
 OAI21_X1 _46680_ (.A(_19641_),
    .B1(_19644_),
    .B2(_19606_),
    .ZN(_04950_));
 NAND2_X1 _46681_ (.A1(_19636_),
    .A2(\icache.lce.lce_cmd_inst.data_r [156]),
    .ZN(_19645_));
 AOI21_X1 _46682_ (.A(_16406_),
    .B1(_17882_),
    .B2(_17886_),
    .ZN(_19646_));
 AOI21_X1 _46683_ (.A(_16314_),
    .B1(_17891_),
    .B2(_17894_),
    .ZN(_19647_));
 OR2_X4 _46684_ (.A1(_19646_),
    .A2(_19647_),
    .ZN(_19648_));
 BUF_X16 _46685_ (.A(_15302_),
    .Z(_19649_));
 BUF_X4 _46686_ (.A(_19649_),
    .Z(_19650_));
 OAI21_X1 _46687_ (.A(_19645_),
    .B1(_19648_),
    .B2(_19650_),
    .ZN(_04951_));
 NAND2_X1 _46688_ (.A1(_19636_),
    .A2(\icache.lce.lce_cmd_inst.data_r [157]),
    .ZN(_19651_));
 AOI21_X2 _46689_ (.A(_19348_),
    .B1(_15904_),
    .B2(_15912_),
    .ZN(_19652_));
 AOI21_X2 _46690_ (.A(_19525_),
    .B1(_15918_),
    .B2(_15924_),
    .ZN(_19653_));
 NOR2_X4 _46691_ (.A1(_19652_),
    .A2(_19653_),
    .ZN(_19654_));
 OAI21_X1 _46692_ (.A(_19651_),
    .B1(_19654_),
    .B2(_19650_),
    .ZN(_04952_));
 NAND2_X1 _46693_ (.A1(_19636_),
    .A2(\icache.lce.lce_cmd_inst.data_r [158]),
    .ZN(_19655_));
 AND3_X1 _46694_ (.A1(_15944_),
    .A2(_15522_),
    .A3(_15948_),
    .ZN(_19656_));
 AOI21_X1 _46695_ (.A(_18419_),
    .B1(_15933_),
    .B2(_15939_),
    .ZN(_19657_));
 OR2_X4 _46696_ (.A1(_19656_),
    .A2(_19657_),
    .ZN(_19658_));
 OAI21_X1 _46697_ (.A(_19655_),
    .B1(_19658_),
    .B2(_19650_),
    .ZN(_04953_));
 NAND2_X1 _46698_ (.A1(_19636_),
    .A2(\icache.lce.lce_cmd_inst.data_r [159]),
    .ZN(_19659_));
 AND3_X1 _46699_ (.A1(_15966_),
    .A2(_15970_),
    .A3(_15503_),
    .ZN(_19660_));
 AOI21_X2 _46700_ (.A(_19425_),
    .B1(_15957_),
    .B2(_15962_),
    .ZN(_19661_));
 NOR2_X4 _46701_ (.A1(_19660_),
    .A2(_19661_),
    .ZN(_19662_));
 OAI21_X1 _46702_ (.A(_19659_),
    .B1(_19662_),
    .B2(_19650_),
    .ZN(_04954_));
 NAND2_X1 _46703_ (.A1(_19636_),
    .A2(\icache.lce.lce_cmd_inst.data_r [160]),
    .ZN(_19663_));
 AOI21_X2 _46704_ (.A(_15368_),
    .B1(_15976_),
    .B2(_15980_),
    .ZN(_19664_));
 AOI21_X2 _46705_ (.A(_19525_),
    .B1(_15989_),
    .B2(_15995_),
    .ZN(_19665_));
 NOR2_X4 _46706_ (.A1(_19664_),
    .A2(_19665_),
    .ZN(_19666_));
 OAI21_X1 _46707_ (.A(_19663_),
    .B1(_19666_),
    .B2(_19650_),
    .ZN(_04956_));
 NAND2_X1 _46708_ (.A1(_19636_),
    .A2(\icache.lce.lce_cmd_inst.data_r [161]),
    .ZN(_19667_));
 OAI21_X2 _46709_ (.A(_19366_),
    .B1(_16004_),
    .B2(_16010_),
    .ZN(_19668_));
 OAI21_X2 _46710_ (.A(_19595_),
    .B1(_16020_),
    .B2(_16026_),
    .ZN(_19669_));
 NAND2_X4 _46711_ (.A1(_19668_),
    .A2(_19669_),
    .ZN(_19670_));
 OAI21_X1 _46712_ (.A(_19667_),
    .B1(_19670_),
    .B2(_19650_),
    .ZN(_04957_));
 NAND2_X1 _46713_ (.A1(_19636_),
    .A2(\icache.lce.lce_cmd_inst.data_r [162]),
    .ZN(_19671_));
 AND3_X2 _46714_ (.A1(_16032_),
    .A2(_15621_),
    .A3(_16037_),
    .ZN(_19672_));
 AOI21_X2 _46715_ (.A(_19525_),
    .B1(_16041_),
    .B2(_16045_),
    .ZN(_19673_));
 NOR2_X4 _46716_ (.A1(_19672_),
    .A2(_19673_),
    .ZN(_19674_));
 OAI21_X1 _46717_ (.A(_19671_),
    .B1(_19674_),
    .B2(_19650_),
    .ZN(_04958_));
 NAND2_X1 _46718_ (.A1(_19636_),
    .A2(\icache.lce.lce_cmd_inst.data_r [163]),
    .ZN(_19675_));
 AND3_X1 _46719_ (.A1(_16054_),
    .A2(_18805_),
    .A3(_16058_),
    .ZN(_19676_));
 AOI21_X2 _46720_ (.A(_19425_),
    .B1(_16063_),
    .B2(_16069_),
    .ZN(_19677_));
 NOR2_X4 _46721_ (.A1(_19676_),
    .A2(_19677_),
    .ZN(_19678_));
 OAI21_X1 _46722_ (.A(_19675_),
    .B1(_19678_),
    .B2(_19650_),
    .ZN(_04959_));
 BUF_X4 _46723_ (.A(_19635_),
    .Z(_19679_));
 NAND2_X1 _46724_ (.A1(_19679_),
    .A2(\icache.lce.lce_cmd_inst.data_r [164]),
    .ZN(_19680_));
 AOI21_X2 _46725_ (.A(_19505_),
    .B1(_16076_),
    .B2(_16081_),
    .ZN(_19681_));
 BUF_X16 _46726_ (.A(_15367_),
    .Z(_19682_));
 AOI21_X2 _46727_ (.A(_19682_),
    .B1(_16087_),
    .B2(_16092_),
    .ZN(_19683_));
 NOR2_X4 _46728_ (.A1(_19681_),
    .A2(_19683_),
    .ZN(_19684_));
 OAI21_X1 _46729_ (.A(_19680_),
    .B1(_19684_),
    .B2(_19650_),
    .ZN(_04960_));
 NAND2_X1 _46730_ (.A1(_19679_),
    .A2(\icache.lce.lce_cmd_inst.data_r [165]),
    .ZN(_19685_));
 AOI21_X2 _46731_ (.A(_15368_),
    .B1(_16098_),
    .B2(_16103_),
    .ZN(_19686_));
 AOI21_X2 _46732_ (.A(_19525_),
    .B1(_16108_),
    .B2(_16114_),
    .ZN(_19687_));
 NOR2_X4 _46733_ (.A1(_19686_),
    .A2(_19687_),
    .ZN(_19688_));
 OAI21_X1 _46734_ (.A(_19685_),
    .B1(_19688_),
    .B2(_19650_),
    .ZN(_04961_));
 NAND2_X1 _46735_ (.A1(_19679_),
    .A2(\icache.lce.lce_cmd_inst.data_r [166]),
    .ZN(_19689_));
 AND3_X1 _46736_ (.A1(_16121_),
    .A2(_15621_),
    .A3(_16124_),
    .ZN(_19690_));
 AOI21_X2 _46737_ (.A(_19525_),
    .B1(_16128_),
    .B2(_16132_),
    .ZN(_19691_));
 NOR2_X4 _46738_ (.A1(_19690_),
    .A2(_19691_),
    .ZN(_19692_));
 BUF_X4 _46739_ (.A(_19649_),
    .Z(_19693_));
 OAI21_X1 _46740_ (.A(_19689_),
    .B1(_19692_),
    .B2(_19693_),
    .ZN(_04962_));
 NAND2_X1 _46741_ (.A1(_19679_),
    .A2(\icache.lce.lce_cmd_inst.data_r [167]),
    .ZN(_19694_));
 AOI21_X2 _46742_ (.A(_15368_),
    .B1(_16138_),
    .B2(_16142_),
    .ZN(_19695_));
 BUF_X16 _46743_ (.A(_15833_),
    .Z(_19696_));
 AOI21_X2 _46744_ (.A(_19696_),
    .B1(_16147_),
    .B2(_16151_),
    .ZN(_19697_));
 NOR2_X4 _46745_ (.A1(_19695_),
    .A2(_19697_),
    .ZN(_19698_));
 OAI21_X1 _46746_ (.A(_19694_),
    .B1(_19698_),
    .B2(_19693_),
    .ZN(_04963_));
 NAND2_X1 _46747_ (.A1(_19679_),
    .A2(\icache.lce.lce_cmd_inst.data_r [168]),
    .ZN(_19699_));
 NAND3_X2 _46748_ (.A1(_16158_),
    .A2(_16161_),
    .A3(_15645_),
    .ZN(_19700_));
 NAND3_X2 _46749_ (.A1(_16165_),
    .A2(_18918_),
    .A3(_16171_),
    .ZN(_19701_));
 NAND2_X4 _46750_ (.A1(_19700_),
    .A2(_19701_),
    .ZN(_19702_));
 OAI21_X1 _46751_ (.A(_19699_),
    .B1(_19702_),
    .B2(_19693_),
    .ZN(_04964_));
 NAND2_X1 _46752_ (.A1(_19679_),
    .A2(\icache.lce.lce_cmd_inst.data_r [169]),
    .ZN(_19703_));
 AND3_X1 _46753_ (.A1(_16189_),
    .A2(_16196_),
    .A3(_15503_),
    .ZN(_19704_));
 AOI21_X2 _46754_ (.A(_19682_),
    .B1(_16178_),
    .B2(_16183_),
    .ZN(_19705_));
 NOR2_X4 _46755_ (.A1(_19704_),
    .A2(_19705_),
    .ZN(_19706_));
 OAI21_X1 _46756_ (.A(_19703_),
    .B1(_19706_),
    .B2(_19693_),
    .ZN(_04965_));
 NAND2_X1 _46757_ (.A1(_19679_),
    .A2(\icache.lce.lce_cmd_inst.data_r [170]),
    .ZN(_19707_));
 AOI21_X2 _46758_ (.A(_19505_),
    .B1(_16203_),
    .B2(_16207_),
    .ZN(_19708_));
 AOI21_X2 _46759_ (.A(_19682_),
    .B1(_16213_),
    .B2(_16218_),
    .ZN(_19709_));
 NOR2_X4 _46760_ (.A1(_19708_),
    .A2(_19709_),
    .ZN(_19710_));
 OAI21_X1 _46761_ (.A(_19707_),
    .B1(_19710_),
    .B2(_19693_),
    .ZN(_04967_));
 NAND2_X1 _46762_ (.A1(_19679_),
    .A2(\icache.lce.lce_cmd_inst.data_r [171]),
    .ZN(_19711_));
 OAI21_X2 _46763_ (.A(_19510_),
    .B1(_16228_),
    .B2(_16235_),
    .ZN(_19712_));
 OAI21_X2 _46764_ (.A(_19088_),
    .B1(_16242_),
    .B2(_16247_),
    .ZN(_19713_));
 NAND2_X4 _46765_ (.A1(_19712_),
    .A2(_19713_),
    .ZN(_19714_));
 OAI21_X1 _46766_ (.A(_19711_),
    .B1(_19714_),
    .B2(_19693_),
    .ZN(_04968_));
 NAND2_X1 _46767_ (.A1(_19679_),
    .A2(\icache.lce.lce_cmd_inst.data_r [172]),
    .ZN(_19715_));
 NAND2_X1 _46768_ (.A1(_16264_),
    .A2(_19579_),
    .ZN(_19716_));
 OAI21_X4 _46769_ (.A(_19088_),
    .B1(_16271_),
    .B2(_16276_),
    .ZN(_19717_));
 NAND2_X4 _46770_ (.A1(_19716_),
    .A2(_19717_),
    .ZN(_19718_));
 OAI21_X1 _46771_ (.A(_19715_),
    .B1(_19718_),
    .B2(_19693_),
    .ZN(_04969_));
 NAND2_X1 _46772_ (.A1(_19679_),
    .A2(\icache.lce.lce_cmd_inst.data_r [173]),
    .ZN(_19719_));
 AND3_X1 _46773_ (.A1(_16283_),
    .A2(_16287_),
    .A3(_16562_),
    .ZN(_19720_));
 AOI21_X2 _46774_ (.A(_19696_),
    .B1(_16291_),
    .B2(_16294_),
    .ZN(_19721_));
 NOR2_X4 _46775_ (.A1(_19720_),
    .A2(_19721_),
    .ZN(_19722_));
 OAI21_X1 _46776_ (.A(_19719_),
    .B1(_19722_),
    .B2(_19693_),
    .ZN(_04970_));
 BUF_X4 _46777_ (.A(_19635_),
    .Z(_19723_));
 NAND2_X1 _46778_ (.A1(_19723_),
    .A2(\icache.lce.lce_cmd_inst.data_r [174]),
    .ZN(_19724_));
 NAND3_X1 _46779_ (.A1(_16301_),
    .A2(_16305_),
    .A3(_15409_),
    .ZN(_19725_));
 OAI21_X1 _46780_ (.A(_19183_),
    .B1(_16310_),
    .B2(_16313_),
    .ZN(_19726_));
 AND2_X2 _46781_ (.A1(_19725_),
    .A2(_19726_),
    .ZN(_19727_));
 OAI21_X1 _46782_ (.A(_19724_),
    .B1(_19727_),
    .B2(_19693_),
    .ZN(_04971_));
 NAND2_X1 _46783_ (.A1(_19723_),
    .A2(\icache.lce.lce_cmd_inst.data_r [175]),
    .ZN(_19728_));
 AND3_X1 _46784_ (.A1(_16322_),
    .A2(_15621_),
    .A3(_16325_),
    .ZN(_19729_));
 AOI21_X2 _46785_ (.A(_19696_),
    .B1(_16330_),
    .B2(_16333_),
    .ZN(_19730_));
 NOR2_X4 _46786_ (.A1(_19729_),
    .A2(_19730_),
    .ZN(_19731_));
 OAI21_X1 _46787_ (.A(_19728_),
    .B1(_19731_),
    .B2(_19693_),
    .ZN(_04972_));
 NAND2_X1 _46788_ (.A1(_19723_),
    .A2(\icache.lce.lce_cmd_inst.data_r [176]),
    .ZN(_19732_));
 NAND2_X1 _46789_ (.A1(_16349_),
    .A2(_19579_),
    .ZN(_19733_));
 OAI21_X2 _46790_ (.A(_19088_),
    .B1(_16353_),
    .B2(_16356_),
    .ZN(_19734_));
 NAND2_X4 _46791_ (.A1(_19733_),
    .A2(_19734_),
    .ZN(_19735_));
 BUF_X4 _46792_ (.A(_19649_),
    .Z(_19736_));
 OAI21_X1 _46793_ (.A(_19732_),
    .B1(_19735_),
    .B2(_19736_),
    .ZN(_04973_));
 NAND2_X1 _46794_ (.A1(_19723_),
    .A2(\icache.lce.lce_cmd_inst.data_r [177]),
    .ZN(_19737_));
 NOR3_X1 _46795_ (.A1(_16363_),
    .A2(_16366_),
    .A3(_16265_),
    .ZN(_19738_));
 AOI21_X1 _46796_ (.A(_16314_),
    .B1(_16371_),
    .B2(_16375_),
    .ZN(_19739_));
 OR2_X2 _46797_ (.A1(_19738_),
    .A2(_19739_),
    .ZN(_19740_));
 OAI21_X1 _46798_ (.A(_19737_),
    .B1(_19740_),
    .B2(_19736_),
    .ZN(_04974_));
 NAND2_X1 _46799_ (.A1(_19723_),
    .A2(\icache.lce.lce_cmd_inst.data_r [178]),
    .ZN(_19741_));
 OR3_X1 _46800_ (.A1(_16381_),
    .A2(_16012_),
    .A3(_16384_),
    .ZN(_19742_));
 NAND3_X2 _46801_ (.A1(_16389_),
    .A2(_18918_),
    .A3(_16397_),
    .ZN(_19743_));
 NAND2_X4 _46802_ (.A1(_19742_),
    .A2(_19743_),
    .ZN(_19744_));
 OAI21_X1 _46803_ (.A(_19741_),
    .B1(_19744_),
    .B2(_19736_),
    .ZN(_04975_));
 NAND2_X1 _46804_ (.A1(_19723_),
    .A2(\icache.lce.lce_cmd_inst.data_r [179]),
    .ZN(_19745_));
 OAI21_X1 _46805_ (.A(_19179_),
    .B1(_16405_),
    .B2(_16410_),
    .ZN(_19746_));
 NAND3_X1 _46806_ (.A1(_16414_),
    .A2(_16372_),
    .A3(_16419_),
    .ZN(_19747_));
 AND2_X4 _46807_ (.A1(_19746_),
    .A2(_19747_),
    .ZN(_19748_));
 OAI21_X1 _46808_ (.A(_19745_),
    .B1(_19748_),
    .B2(_19736_),
    .ZN(_04976_));
 NAND2_X1 _46809_ (.A1(_19723_),
    .A2(\icache.lce.lce_cmd_inst.data_r [180]),
    .ZN(_19749_));
 NAND3_X1 _46810_ (.A1(_16425_),
    .A2(_16360_),
    .A3(_16428_),
    .ZN(_19750_));
 NAND3_X1 _46811_ (.A1(_16431_),
    .A2(_16640_),
    .A3(_16434_),
    .ZN(_19751_));
 AND2_X4 _46812_ (.A1(_19750_),
    .A2(_19751_),
    .ZN(_19752_));
 OAI21_X1 _46813_ (.A(_19749_),
    .B1(_19752_),
    .B2(_19736_),
    .ZN(_04978_));
 NAND2_X1 _46814_ (.A1(_19723_),
    .A2(\icache.lce.lce_cmd_inst.data_r [181]),
    .ZN(_19753_));
 OAI21_X1 _46815_ (.A(_19179_),
    .B1(_16440_),
    .B2(_16443_),
    .ZN(_19754_));
 NAND3_X1 _46816_ (.A1(_16448_),
    .A2(_16452_),
    .A3(_15315_),
    .ZN(_19755_));
 AND2_X4 _46817_ (.A1(_19754_),
    .A2(_19755_),
    .ZN(_19756_));
 OAI21_X1 _46818_ (.A(_19753_),
    .B1(_19756_),
    .B2(_19736_),
    .ZN(_04979_));
 NAND2_X1 _46819_ (.A1(_19723_),
    .A2(\icache.lce.lce_cmd_inst.data_r [182]),
    .ZN(_19757_));
 NAND2_X1 _46820_ (.A1(_16464_),
    .A2(_19593_),
    .ZN(_19758_));
 OAI21_X2 _46821_ (.A(_19595_),
    .B1(_16468_),
    .B2(_16471_),
    .ZN(_19759_));
 NAND2_X4 _46822_ (.A1(_19758_),
    .A2(_19759_),
    .ZN(_19760_));
 OAI21_X1 _46823_ (.A(_19757_),
    .B1(_19760_),
    .B2(_19736_),
    .ZN(_04980_));
 NAND2_X1 _46824_ (.A1(_19723_),
    .A2(\icache.lce.lce_cmd_inst.data_r [183]),
    .ZN(_19761_));
 OAI21_X2 _46825_ (.A(_19510_),
    .B1(_16477_),
    .B2(_16480_),
    .ZN(_19762_));
 NAND3_X2 _46826_ (.A1(_16484_),
    .A2(_18918_),
    .A3(_16487_),
    .ZN(_19763_));
 NAND2_X4 _46827_ (.A1(_19762_),
    .A2(_19763_),
    .ZN(_19764_));
 OAI21_X1 _46828_ (.A(_19761_),
    .B1(_19764_),
    .B2(_19736_),
    .ZN(_04981_));
 BUF_X16 _46829_ (.A(_19635_),
    .Z(_19765_));
 NAND2_X1 _46830_ (.A1(_19765_),
    .A2(\icache.lce.lce_cmd_inst.data_r [184]),
    .ZN(_19766_));
 AND3_X1 _46831_ (.A1(_16494_),
    .A2(_16498_),
    .A3(_15686_),
    .ZN(_19767_));
 AOI21_X2 _46832_ (.A(_19696_),
    .B1(_16502_),
    .B2(_16505_),
    .ZN(_19768_));
 NOR2_X4 _46833_ (.A1(_19767_),
    .A2(_19768_),
    .ZN(_19769_));
 OAI21_X1 _46834_ (.A(_19766_),
    .B1(_19769_),
    .B2(_19736_),
    .ZN(_04982_));
 NAND2_X1 _46835_ (.A1(_19765_),
    .A2(\icache.lce.lce_cmd_inst.data_r [185]),
    .ZN(_19770_));
 OAI21_X1 _46836_ (.A(_18922_),
    .B1(_16513_),
    .B2(_16516_),
    .ZN(_19771_));
 NAND3_X1 _46837_ (.A1(_16521_),
    .A2(_16525_),
    .A3(_15849_),
    .ZN(_19772_));
 AND2_X4 _46838_ (.A1(_19771_),
    .A2(_19772_),
    .ZN(_19773_));
 OAI21_X1 _46839_ (.A(_19770_),
    .B1(_19773_),
    .B2(_19736_),
    .ZN(_04983_));
 NAND2_X1 _46840_ (.A1(_19765_),
    .A2(\icache.lce.lce_cmd_inst.data_r [186]),
    .ZN(_19774_));
 NAND2_X1 _46841_ (.A1(_16538_),
    .A2(_19579_),
    .ZN(_19775_));
 OAI21_X2 _46842_ (.A(_19088_),
    .B1(_16543_),
    .B2(_16547_),
    .ZN(_19776_));
 NAND2_X4 _46843_ (.A1(_19775_),
    .A2(_19776_),
    .ZN(_19777_));
 BUF_X16 _46844_ (.A(_19649_),
    .Z(_19778_));
 OAI21_X1 _46845_ (.A(_19774_),
    .B1(_19777_),
    .B2(_19778_),
    .ZN(_04984_));
 NAND2_X1 _46846_ (.A1(_19765_),
    .A2(\icache.lce.lce_cmd_inst.data_r [187]),
    .ZN(_19779_));
 AND3_X1 _46847_ (.A1(_16555_),
    .A2(_16561_),
    .A3(_15503_),
    .ZN(_19780_));
 AOI21_X2 _46848_ (.A(_19682_),
    .B1(_16568_),
    .B2(_16572_),
    .ZN(_19781_));
 NOR2_X4 _46849_ (.A1(_19780_),
    .A2(_19781_),
    .ZN(_19782_));
 OAI21_X1 _46850_ (.A(_19779_),
    .B1(_19782_),
    .B2(_19778_),
    .ZN(_04985_));
 NAND2_X1 _46851_ (.A1(_19765_),
    .A2(\icache.lce.lce_cmd_inst.data_r [188]),
    .ZN(_19783_));
 AOI21_X2 _46852_ (.A(_19505_),
    .B1(_16588_),
    .B2(_16592_),
    .ZN(_19784_));
 AOI21_X2 _46853_ (.A(_19682_),
    .B1(_16579_),
    .B2(_16584_),
    .ZN(_19785_));
 NOR2_X4 _46854_ (.A1(_19784_),
    .A2(_19785_),
    .ZN(_19786_));
 OAI21_X1 _46855_ (.A(_19783_),
    .B1(_19786_),
    .B2(_19778_),
    .ZN(_04986_));
 NAND2_X1 _46856_ (.A1(_19765_),
    .A2(\icache.lce.lce_cmd_inst.data_r [189]),
    .ZN(_19787_));
 AND3_X1 _46857_ (.A1(_16599_),
    .A2(_15621_),
    .A3(_16603_),
    .ZN(_19788_));
 AOI21_X2 _46858_ (.A(_19696_),
    .B1(_16607_),
    .B2(_16610_),
    .ZN(_19789_));
 NOR2_X2 _46859_ (.A1(_19788_),
    .A2(_19789_),
    .ZN(_19790_));
 OAI21_X1 _46860_ (.A(_19787_),
    .B1(_19790_),
    .B2(_19778_),
    .ZN(_04987_));
 NAND2_X1 _46861_ (.A1(_19765_),
    .A2(\icache.lce.lce_cmd_inst.data_r [190]),
    .ZN(_19791_));
 OAI21_X1 _46862_ (.A(_19366_),
    .B1(_16616_),
    .B2(_16619_),
    .ZN(_19792_));
 NAND3_X1 _46863_ (.A1(_16624_),
    .A2(_18747_),
    .A3(_16627_),
    .ZN(_19793_));
 NAND2_X2 _46864_ (.A1(_19792_),
    .A2(_19793_),
    .ZN(_19794_));
 OAI21_X1 _46865_ (.A(_19791_),
    .B1(_19794_),
    .B2(_19778_),
    .ZN(_04989_));
 NAND2_X1 _46866_ (.A1(_19765_),
    .A2(\icache.lce.lce_cmd_inst.data_r [191]),
    .ZN(_19795_));
 OAI21_X1 _46867_ (.A(_19179_),
    .B1(_16644_),
    .B2(_16647_),
    .ZN(_19796_));
 OAI21_X1 _46868_ (.A(_19183_),
    .B1(_16635_),
    .B2(_16638_),
    .ZN(_19797_));
 AND2_X4 _46869_ (.A1(_19796_),
    .A2(_19797_),
    .ZN(_19798_));
 OAI21_X1 _46870_ (.A(_19795_),
    .B1(_19798_),
    .B2(_19778_),
    .ZN(_04990_));
 NAND2_X1 _46871_ (.A1(_19765_),
    .A2(\icache.lce.lce_cmd_inst.data_r [192]),
    .ZN(_19799_));
 AND3_X1 _46872_ (.A1(_16653_),
    .A2(_16656_),
    .A3(_15522_),
    .ZN(_19800_));
 AOI21_X2 _46873_ (.A(_18419_),
    .B1(_16660_),
    .B2(_16663_),
    .ZN(_19801_));
 OR2_X4 _46874_ (.A1(_19800_),
    .A2(_19801_),
    .ZN(_19802_));
 OAI21_X1 _46875_ (.A(_19799_),
    .B1(_19802_),
    .B2(_19778_),
    .ZN(_04991_));
 NAND2_X1 _46876_ (.A1(_19765_),
    .A2(\icache.lce.lce_cmd_inst.data_r [97]),
    .ZN(_19803_));
 NAND2_X1 _46877_ (.A1(_18299_),
    .A2(_19593_),
    .ZN(_19804_));
 NAND3_X2 _46878_ (.A1(_18301_),
    .A2(_18747_),
    .A3(_18302_),
    .ZN(_19805_));
 NAND2_X4 _46879_ (.A1(_19804_),
    .A2(_19805_),
    .ZN(_19806_));
 OAI21_X1 _46880_ (.A(_19803_),
    .B1(_19806_),
    .B2(_19778_),
    .ZN(_05397_));
 BUF_X4 _46881_ (.A(_19635_),
    .Z(_19807_));
 NAND2_X1 _46882_ (.A1(_19807_),
    .A2(\icache.lce.lce_cmd_inst.data_r [98]),
    .ZN(_19808_));
 OAI21_X1 _46883_ (.A(_19179_),
    .B1(_18307_),
    .B2(_18308_),
    .ZN(_19809_));
 NAND3_X1 _46884_ (.A1(_18310_),
    .A2(_16640_),
    .A3(_18312_),
    .ZN(_19810_));
 AND2_X4 _46885_ (.A1(_19809_),
    .A2(_19810_),
    .ZN(_19811_));
 OAI21_X1 _46886_ (.A(_19808_),
    .B1(_19811_),
    .B2(_19778_),
    .ZN(_05398_));
 NAND2_X1 _46887_ (.A1(_19807_),
    .A2(\icache.lce.lce_cmd_inst.data_r [99]),
    .ZN(_19812_));
 AOI21_X1 _46888_ (.A(_18351_),
    .B1(_18316_),
    .B2(_18317_),
    .ZN(_19813_));
 NOR3_X2 _46889_ (.A1(_18319_),
    .A2(_18320_),
    .A3(_15597_),
    .ZN(_19814_));
 OR2_X4 _46890_ (.A1(_19813_),
    .A2(_19814_),
    .ZN(_19815_));
 OAI21_X1 _46891_ (.A(_19812_),
    .B1(_19815_),
    .B2(_19778_),
    .ZN(_05399_));
 NAND2_X1 _46892_ (.A1(_19807_),
    .A2(\icache.lce.lce_cmd_inst.data_r [100]),
    .ZN(_19816_));
 OAI21_X2 _46893_ (.A(_19510_),
    .B1(_18325_),
    .B2(_18326_),
    .ZN(_19817_));
 NAND3_X2 _46894_ (.A1(_18328_),
    .A2(_18330_),
    .A3(_18470_),
    .ZN(_19818_));
 NAND2_X4 _46895_ (.A1(_19817_),
    .A2(_19818_),
    .ZN(_19819_));
 BUF_X8 _46896_ (.A(_19649_),
    .Z(_19820_));
 OAI21_X1 _46897_ (.A(_19816_),
    .B1(_19819_),
    .B2(_19820_),
    .ZN(_04890_));
 NAND2_X1 _46898_ (.A1(_19807_),
    .A2(\icache.lce.lce_cmd_inst.data_r [101]),
    .ZN(_19821_));
 NAND2_X1 _46899_ (.A1(_18336_),
    .A2(_19593_),
    .ZN(_19822_));
 OAI21_X2 _46900_ (.A(_19595_),
    .B1(_18338_),
    .B2(_18339_),
    .ZN(_19823_));
 NAND2_X4 _46901_ (.A1(_19822_),
    .A2(_19823_),
    .ZN(_19824_));
 OAI21_X1 _46902_ (.A(_19821_),
    .B1(_19824_),
    .B2(_19820_),
    .ZN(_04891_));
 NAND2_X1 _46903_ (.A1(_19807_),
    .A2(\icache.lce.lce_cmd_inst.data_r [102]),
    .ZN(_19825_));
 NOR3_X1 _46904_ (.A1(_18343_),
    .A2(_16265_),
    .A3(_18344_),
    .ZN(_19826_));
 AOI21_X1 _46905_ (.A(_16314_),
    .B1(_18346_),
    .B2(_18347_),
    .ZN(_19827_));
 OR2_X2 _46906_ (.A1(_19826_),
    .A2(_19827_),
    .ZN(_19828_));
 OAI21_X1 _46907_ (.A(_19825_),
    .B1(_19828_),
    .B2(_19820_),
    .ZN(_04892_));
 NAND2_X1 _46908_ (.A1(_19807_),
    .A2(\icache.lce.lce_cmd_inst.data_r [103]),
    .ZN(_19829_));
 NAND3_X1 _46909_ (.A1(_18352_),
    .A2(_16438_),
    .A3(_18353_),
    .ZN(_19830_));
 NAND3_X1 _46910_ (.A1(_18355_),
    .A2(_17415_),
    .A3(_18357_),
    .ZN(_19831_));
 AND2_X2 _46911_ (.A1(_19830_),
    .A2(_19831_),
    .ZN(_19832_));
 OAI21_X1 _46912_ (.A(_19829_),
    .B1(_19832_),
    .B2(_19820_),
    .ZN(_04893_));
 NAND2_X1 _46913_ (.A1(_19807_),
    .A2(\icache.lce.lce_cmd_inst.data_r [104]),
    .ZN(_19833_));
 OAI21_X1 _46914_ (.A(_19179_),
    .B1(_18363_),
    .B2(_18364_),
    .ZN(_19834_));
 OAI21_X1 _46915_ (.A(_19183_),
    .B1(_18367_),
    .B2(_18368_),
    .ZN(_19835_));
 AND2_X2 _46916_ (.A1(_19834_),
    .A2(_19835_),
    .ZN(_19836_));
 OAI21_X1 _46917_ (.A(_19833_),
    .B1(_19836_),
    .B2(_19820_),
    .ZN(_04894_));
 NAND2_X1 _46918_ (.A1(_19807_),
    .A2(\icache.lce.lce_cmd_inst.data_r [105]),
    .ZN(_19837_));
 OR3_X1 _46919_ (.A1(_18377_),
    .A2(_18378_),
    .A3(_15314_),
    .ZN(_19838_));
 OAI21_X1 _46920_ (.A(_19183_),
    .B1(_18373_),
    .B2(_18374_),
    .ZN(_19839_));
 AND2_X2 _46921_ (.A1(_19838_),
    .A2(_19839_),
    .ZN(_19840_));
 OAI21_X1 _46922_ (.A(_19837_),
    .B1(_19840_),
    .B2(_19820_),
    .ZN(_04895_));
 NAND2_X1 _46923_ (.A1(_19807_),
    .A2(\icache.lce.lce_cmd_inst.data_r [106]),
    .ZN(_19841_));
 OR3_X1 _46924_ (.A1(_18382_),
    .A2(_18384_),
    .A3(_15699_),
    .ZN(_19842_));
 OAI21_X2 _46925_ (.A(_19595_),
    .B1(_18386_),
    .B2(_18387_),
    .ZN(_19843_));
 NAND2_X4 _46926_ (.A1(_19842_),
    .A2(_19843_),
    .ZN(_19844_));
 OAI21_X1 _46927_ (.A(_19841_),
    .B1(_19844_),
    .B2(_19820_),
    .ZN(_04896_));
 NAND2_X1 _46928_ (.A1(_19807_),
    .A2(\icache.lce.lce_cmd_inst.data_r [107]),
    .ZN(_19845_));
 NAND3_X1 _46929_ (.A1(_18392_),
    .A2(_18393_),
    .A3(_15409_),
    .ZN(_19846_));
 OAI21_X1 _46930_ (.A(_19183_),
    .B1(_18395_),
    .B2(_18396_),
    .ZN(_19847_));
 AND2_X2 _46931_ (.A1(_19846_),
    .A2(_19847_),
    .ZN(_19848_));
 OAI21_X1 _46932_ (.A(_19845_),
    .B1(_19848_),
    .B2(_19820_),
    .ZN(_04897_));
 BUF_X8 _46933_ (.A(_19635_),
    .Z(_19849_));
 NAND2_X1 _46934_ (.A1(_19849_),
    .A2(\icache.lce.lce_cmd_inst.data_r [108]),
    .ZN(_19850_));
 AND3_X1 _46935_ (.A1(_18400_),
    .A2(_18401_),
    .A3(_15686_),
    .ZN(_19851_));
 AOI21_X2 _46936_ (.A(_19696_),
    .B1(_18403_),
    .B2(_18404_),
    .ZN(_19852_));
 NOR2_X4 _46937_ (.A1(_19851_),
    .A2(_19852_),
    .ZN(_19853_));
 OAI21_X1 _46938_ (.A(_19850_),
    .B1(_19853_),
    .B2(_19820_),
    .ZN(_04898_));
 NAND2_X1 _46939_ (.A1(_19849_),
    .A2(\icache.lce.lce_cmd_inst.data_r [109]),
    .ZN(_19854_));
 AND3_X1 _46940_ (.A1(_18408_),
    .A2(_18805_),
    .A3(_18409_),
    .ZN(_19855_));
 AOI21_X2 _46941_ (.A(_19682_),
    .B1(_18411_),
    .B2(_18412_),
    .ZN(_19856_));
 NOR2_X4 _46942_ (.A1(_19855_),
    .A2(_19856_),
    .ZN(_19857_));
 OAI21_X1 _46943_ (.A(_19854_),
    .B1(_19857_),
    .B2(_19820_),
    .ZN(_04899_));
 NAND2_X1 _46944_ (.A1(_19849_),
    .A2(\icache.lce.lce_cmd_inst.data_r [110]),
    .ZN(_19858_));
 AND3_X1 _46945_ (.A1(_18420_),
    .A2(_18805_),
    .A3(_18421_),
    .ZN(_19859_));
 AOI21_X2 _46946_ (.A(_19682_),
    .B1(_18416_),
    .B2(_18417_),
    .ZN(_19860_));
 NOR2_X4 _46947_ (.A1(_19859_),
    .A2(_19860_),
    .ZN(_19861_));
 BUF_X16 _46948_ (.A(_19649_),
    .Z(_19862_));
 OAI21_X1 _46949_ (.A(_19858_),
    .B1(_19861_),
    .B2(_19862_),
    .ZN(_04901_));
 NAND2_X1 _46950_ (.A1(_19849_),
    .A2(\icache.lce.lce_cmd_inst.data_r [111]),
    .ZN(_19863_));
 NAND2_X1 _46951_ (.A1(_18431_),
    .A2(_19579_),
    .ZN(_19864_));
 NAND2_X1 _46952_ (.A1(_18427_),
    .A2(_15905_),
    .ZN(_19865_));
 NAND2_X2 _46953_ (.A1(_19864_),
    .A2(_19865_),
    .ZN(_19866_));
 OAI21_X1 _46954_ (.A(_19863_),
    .B1(_19866_),
    .B2(_19862_),
    .ZN(_04902_));
 NAND2_X1 _46955_ (.A1(_19849_),
    .A2(\icache.lce.lce_cmd_inst.data_r [112]),
    .ZN(_19867_));
 NAND2_X1 _46956_ (.A1(_18437_),
    .A2(_19593_),
    .ZN(_19868_));
 NAND3_X2 _46957_ (.A1(_18439_),
    .A2(_18747_),
    .A3(_18440_),
    .ZN(_19869_));
 NAND2_X4 _46958_ (.A1(_19868_),
    .A2(_19869_),
    .ZN(_19870_));
 OAI21_X1 _46959_ (.A(_19867_),
    .B1(_19870_),
    .B2(_19862_),
    .ZN(_04903_));
 NAND2_X1 _46960_ (.A1(_19849_),
    .A2(\icache.lce.lce_cmd_inst.data_r [113]),
    .ZN(_19871_));
 AOI21_X2 _46961_ (.A(_19505_),
    .B1(_18444_),
    .B2(_18445_),
    .ZN(_19872_));
 AOI21_X2 _46962_ (.A(_19682_),
    .B1(_18447_),
    .B2(_18448_),
    .ZN(_19873_));
 NOR2_X4 _46963_ (.A1(_19872_),
    .A2(_19873_),
    .ZN(_19874_));
 OAI21_X1 _46964_ (.A(_19871_),
    .B1(_19874_),
    .B2(_19862_),
    .ZN(_04904_));
 NAND2_X1 _46965_ (.A1(_19849_),
    .A2(\icache.lce.lce_cmd_inst.data_r [114]),
    .ZN(_19875_));
 AOI21_X2 _46966_ (.A(_15368_),
    .B1(_18453_),
    .B2(_18454_),
    .ZN(_19876_));
 AOI21_X2 _46967_ (.A(_19696_),
    .B1(_18457_),
    .B2(_18459_),
    .ZN(_19877_));
 NOR2_X4 _46968_ (.A1(_19876_),
    .A2(_19877_),
    .ZN(_19878_));
 OAI21_X1 _46969_ (.A(_19875_),
    .B1(_19878_),
    .B2(_19862_),
    .ZN(_04905_));
 NAND2_X1 _46970_ (.A1(_19849_),
    .A2(\icache.lce.lce_cmd_inst.data_r [115]),
    .ZN(_19879_));
 AOI21_X1 _46971_ (.A(_19505_),
    .B1(_18464_),
    .B2(_18465_),
    .ZN(_19880_));
 AOI21_X1 _46972_ (.A(_19682_),
    .B1(_18468_),
    .B2(_18469_),
    .ZN(_19881_));
 NOR2_X2 _46973_ (.A1(_19880_),
    .A2(_19881_),
    .ZN(_19882_));
 OAI21_X1 _46974_ (.A(_19879_),
    .B1(_19882_),
    .B2(_19862_),
    .ZN(_04906_));
 NAND2_X1 _46975_ (.A1(_19849_),
    .A2(\icache.lce.lce_cmd_inst.data_r [94]),
    .ZN(_19883_));
 OR3_X2 _46976_ (.A1(_18271_),
    .A2(_15734_),
    .A3(_18272_),
    .ZN(_19884_));
 NAND3_X2 _46977_ (.A1(_18274_),
    .A2(_18275_),
    .A3(_15354_),
    .ZN(_19885_));
 NAND2_X4 _46978_ (.A1(_19884_),
    .A2(_19885_),
    .ZN(_19886_));
 OAI21_X1 _46979_ (.A(_19883_),
    .B1(_19886_),
    .B2(_19862_),
    .ZN(_05394_));
 NAND2_X1 _46980_ (.A1(_19849_),
    .A2(\icache.lce.lce_cmd_inst.data_r [95]),
    .ZN(_19887_));
 AOI21_X2 _46981_ (.A(_19505_),
    .B1(_18279_),
    .B2(_18280_),
    .ZN(_19888_));
 AOI21_X2 _46982_ (.A(_19682_),
    .B1(_18282_),
    .B2(_18283_),
    .ZN(_19889_));
 NOR2_X4 _46983_ (.A1(_19888_),
    .A2(_19889_),
    .ZN(_19890_));
 OAI21_X1 _46984_ (.A(_19887_),
    .B1(_19890_),
    .B2(_19862_),
    .ZN(_05395_));
 BUF_X8 _46985_ (.A(_19635_),
    .Z(_19891_));
 NAND2_X1 _46986_ (.A1(_19891_),
    .A2(\icache.lce.lce_cmd_inst.data_r [96]),
    .ZN(_19892_));
 OAI21_X1 _46987_ (.A(_18922_),
    .B1(_18287_),
    .B2(_18288_),
    .ZN(_19893_));
 NAND3_X1 _46988_ (.A1(_18290_),
    .A2(_18291_),
    .A3(_15849_),
    .ZN(_19894_));
 AND2_X4 _46989_ (.A1(_19893_),
    .A2(_19894_),
    .ZN(_19895_));
 OAI21_X1 _46990_ (.A(_19892_),
    .B1(_19895_),
    .B2(_19862_),
    .ZN(_05396_));
 NAND2_X1 _46991_ (.A1(_19891_),
    .A2(\icache.lce.lce_cmd_inst.data_r [17]),
    .ZN(_19896_));
 NAND2_X1 _46992_ (.A1(_19209_),
    .A2(_19593_),
    .ZN(_19897_));
 NAND3_X2 _46993_ (.A1(_19211_),
    .A2(_18747_),
    .A3(_19212_),
    .ZN(_19898_));
 NAND2_X4 _46994_ (.A1(_19897_),
    .A2(_19898_),
    .ZN(_19899_));
 OAI21_X1 _46995_ (.A(_19896_),
    .B1(_19899_),
    .B2(_19862_),
    .ZN(_04977_));
 NAND2_X1 _46996_ (.A1(_19891_),
    .A2(\icache.lce.lce_cmd_inst.data_r [18]),
    .ZN(_19900_));
 NOR2_X1 _46997_ (.A1(_19218_),
    .A2(_16200_),
    .ZN(_19901_));
 AOI21_X2 _46998_ (.A(_19696_),
    .B1(_19220_),
    .B2(_19221_),
    .ZN(_19902_));
 NOR2_X4 _46999_ (.A1(_19901_),
    .A2(_19902_),
    .ZN(_19903_));
 BUF_X8 _47000_ (.A(_19649_),
    .Z(_19904_));
 OAI21_X1 _47001_ (.A(_19900_),
    .B1(_19903_),
    .B2(_19904_),
    .ZN(_04988_));
 NAND2_X1 _47002_ (.A1(_19891_),
    .A2(\icache.lce.lce_cmd_inst.data_r [19]),
    .ZN(_19905_));
 AND3_X2 _47003_ (.A1(_19226_),
    .A2(_15940_),
    .A3(_19227_),
    .ZN(_19906_));
 BUF_X16 _47004_ (.A(_15408_),
    .Z(_19907_));
 AOI21_X2 _47005_ (.A(_19907_),
    .B1(_19229_),
    .B2(_19230_),
    .ZN(_19908_));
 NOR2_X4 _47006_ (.A1(_19906_),
    .A2(_19908_),
    .ZN(_19909_));
 OAI21_X1 _47007_ (.A(_19905_),
    .B1(_19909_),
    .B2(_19904_),
    .ZN(_04999_));
 NAND2_X1 _47008_ (.A1(_19891_),
    .A2(\icache.lce.lce_cmd_inst.data_r [20]),
    .ZN(_19910_));
 OR3_X1 _47009_ (.A1(_19234_),
    .A2(_15734_),
    .A3(_19235_),
    .ZN(_19911_));
 NAND3_X2 _47010_ (.A1(_19237_),
    .A2(_19239_),
    .A3(_15354_),
    .ZN(_19912_));
 NAND2_X4 _47011_ (.A1(_19911_),
    .A2(_19912_),
    .ZN(_19913_));
 OAI21_X1 _47012_ (.A(_19910_),
    .B1(_19913_),
    .B2(_19904_),
    .ZN(_05011_));
 NAND2_X1 _47013_ (.A1(_19891_),
    .A2(\icache.lce.lce_cmd_inst.data_r [21]),
    .ZN(_19914_));
 AOI21_X2 _47014_ (.A(_15368_),
    .B1(_19243_),
    .B2(_19245_),
    .ZN(_19915_));
 AND3_X1 _47015_ (.A1(_19247_),
    .A2(_16265_),
    .A3(_19249_),
    .ZN(_19916_));
 NOR2_X4 _47016_ (.A1(_19915_),
    .A2(_19916_),
    .ZN(_19917_));
 OAI21_X1 _47017_ (.A(_19914_),
    .B1(_19917_),
    .B2(_19904_),
    .ZN(_05022_));
 NAND2_X1 _47018_ (.A1(_19891_),
    .A2(\icache.lce.lce_cmd_inst.data_r [22]),
    .ZN(_19918_));
 NAND3_X1 _47019_ (.A1(_19253_),
    .A2(_19254_),
    .A3(_15834_),
    .ZN(_19919_));
 OAI21_X1 _47020_ (.A(_18366_),
    .B1(_19256_),
    .B2(_19257_),
    .ZN(_19920_));
 AND2_X4 _47021_ (.A1(_19919_),
    .A2(_19920_),
    .ZN(_19921_));
 OAI21_X1 _47022_ (.A(_19918_),
    .B1(_19921_),
    .B2(_19904_),
    .ZN(_05033_));
 NAND2_X1 _47023_ (.A1(_19891_),
    .A2(\icache.lce.lce_cmd_inst.data_r [23]),
    .ZN(_19922_));
 OAI21_X1 _47024_ (.A(_19366_),
    .B1(_19261_),
    .B2(_19262_),
    .ZN(_19923_));
 OAI21_X2 _47025_ (.A(_19595_),
    .B1(_19264_),
    .B2(_19265_),
    .ZN(_19924_));
 NAND2_X4 _47026_ (.A1(_19923_),
    .A2(_19924_),
    .ZN(_19925_));
 OAI21_X1 _47027_ (.A(_19922_),
    .B1(_19925_),
    .B2(_19904_),
    .ZN(_05044_));
 NAND2_X1 _47028_ (.A1(_19891_),
    .A2(\icache.lce.lce_cmd_inst.data_r [24]),
    .ZN(_19926_));
 OAI21_X2 _47029_ (.A(_19366_),
    .B1(_19269_),
    .B2(_19270_),
    .ZN(_19927_));
 NAND3_X2 _47030_ (.A1(_19272_),
    .A2(_19273_),
    .A3(_15354_),
    .ZN(_19928_));
 NAND2_X4 _47031_ (.A1(_19927_),
    .A2(_19928_),
    .ZN(_19929_));
 OAI21_X1 _47032_ (.A(_19926_),
    .B1(_19929_),
    .B2(_19904_),
    .ZN(_05055_));
 NAND2_X1 _47033_ (.A1(_19891_),
    .A2(\icache.lce.lce_cmd_inst.data_r [25]),
    .ZN(_19930_));
 AOI21_X2 _47034_ (.A(_15329_),
    .B1(_19280_),
    .B2(_19281_),
    .ZN(_19931_));
 AOI21_X2 _47035_ (.A(_19907_),
    .B1(_19277_),
    .B2(_19278_),
    .ZN(_19932_));
 NOR2_X4 _47036_ (.A1(_19931_),
    .A2(_19932_),
    .ZN(_19933_));
 OAI21_X1 _47037_ (.A(_19930_),
    .B1(_19933_),
    .B2(_19904_),
    .ZN(_05066_));
 BUF_X4 _47038_ (.A(_19635_),
    .Z(_19934_));
 NAND2_X1 _47039_ (.A1(_19934_),
    .A2(\icache.lce.lce_cmd_inst.data_r [26]),
    .ZN(_19935_));
 NOR3_X2 _47040_ (.A1(_19286_),
    .A2(_19287_),
    .A3(_18085_),
    .ZN(_19936_));
 AOI21_X2 _47041_ (.A(_19696_),
    .B1(_19289_),
    .B2(_19290_),
    .ZN(_19937_));
 NOR2_X4 _47042_ (.A1(_19936_),
    .A2(_19937_),
    .ZN(_19938_));
 OAI21_X1 _47043_ (.A(_19935_),
    .B1(_19938_),
    .B2(_19904_),
    .ZN(_05077_));
 NAND2_X1 _47044_ (.A1(_19934_),
    .A2(\icache.lce.lce_cmd_inst.data_r [27]),
    .ZN(_19939_));
 OAI21_X2 _47045_ (.A(_19510_),
    .B1(_19294_),
    .B2(_19295_),
    .ZN(_19940_));
 BUF_X16 _47046_ (.A(_16012_),
    .Z(_19941_));
 NAND3_X2 _47047_ (.A1(_19297_),
    .A2(_19941_),
    .A3(_19298_),
    .ZN(_19942_));
 NAND2_X4 _47048_ (.A1(_19940_),
    .A2(_19942_),
    .ZN(_19943_));
 OAI21_X1 _47049_ (.A(_19939_),
    .B1(_19943_),
    .B2(_19904_),
    .ZN(_05088_));
 NAND2_X1 _47050_ (.A1(_19934_),
    .A2(\icache.lce.lce_cmd_inst.data_r [28]),
    .ZN(_19944_));
 NAND2_X1 _47051_ (.A1(_19304_),
    .A2(_19579_),
    .ZN(_19945_));
 NAND2_X1 _47052_ (.A1(_19308_),
    .A2(_15905_),
    .ZN(_19946_));
 NAND2_X4 _47053_ (.A1(_19945_),
    .A2(_19946_),
    .ZN(_19947_));
 BUF_X4 _47054_ (.A(_19649_),
    .Z(_19948_));
 OAI21_X1 _47055_ (.A(_19944_),
    .B1(_19947_),
    .B2(_19948_),
    .ZN(_05099_));
 NAND2_X1 _47056_ (.A1(_19934_),
    .A2(\icache.lce.lce_cmd_inst.data_r [29]),
    .ZN(_19949_));
 OAI21_X1 _47057_ (.A(_19510_),
    .B1(_19313_),
    .B2(_19314_),
    .ZN(_19950_));
 BUF_X16 _47058_ (.A(_15655_),
    .Z(_19951_));
 OAI21_X2 _47059_ (.A(_19951_),
    .B1(_19316_),
    .B2(_19317_),
    .ZN(_19952_));
 NAND2_X4 _47060_ (.A1(_19950_),
    .A2(_19952_),
    .ZN(_19953_));
 OAI21_X1 _47061_ (.A(_19949_),
    .B1(_19953_),
    .B2(_19948_),
    .ZN(_05110_));
 NAND2_X1 _47062_ (.A1(_19934_),
    .A2(\icache.lce.lce_cmd_inst.data_r [30]),
    .ZN(_19954_));
 NAND2_X1 _47063_ (.A1(_19323_),
    .A2(_19579_),
    .ZN(_19955_));
 OAI21_X2 _47064_ (.A(_19951_),
    .B1(_19325_),
    .B2(_19326_),
    .ZN(_19956_));
 NAND2_X4 _47065_ (.A1(_19955_),
    .A2(_19956_),
    .ZN(_19957_));
 OAI21_X1 _47066_ (.A(_19954_),
    .B1(_19957_),
    .B2(_19948_),
    .ZN(_05122_));
 NAND2_X1 _47067_ (.A1(_19934_),
    .A2(\icache.lce.lce_cmd_inst.data_r [31]),
    .ZN(_19958_));
 OAI21_X2 _47068_ (.A(_19510_),
    .B1(_19330_),
    .B2(_19331_),
    .ZN(_19959_));
 NAND3_X2 _47069_ (.A1(_19334_),
    .A2(_19336_),
    .A3(_18470_),
    .ZN(_19960_));
 NAND2_X4 _47070_ (.A1(_19959_),
    .A2(_19960_),
    .ZN(_19961_));
 OAI21_X1 _47071_ (.A(_19958_),
    .B1(_19961_),
    .B2(_19948_),
    .ZN(_05133_));
 NAND2_X1 _47072_ (.A1(_19934_),
    .A2(\icache.lce.lce_cmd_inst.data_r [32]),
    .ZN(_19962_));
 BUF_X16 _47073_ (.A(_15734_),
    .Z(_19963_));
 OAI21_X2 _47074_ (.A(_19963_),
    .B1(_19340_),
    .B2(_19341_),
    .ZN(_19964_));
 OAI21_X2 _47075_ (.A(_19951_),
    .B1(_19343_),
    .B2(_19344_),
    .ZN(_19965_));
 NAND2_X4 _47076_ (.A1(_19964_),
    .A2(_19965_),
    .ZN(_19966_));
 OAI21_X1 _47077_ (.A(_19962_),
    .B1(_19966_),
    .B2(_19948_),
    .ZN(_05144_));
 NAND2_X1 _47078_ (.A1(_19934_),
    .A2(\icache.lce.lce_cmd_inst.data_r [33]),
    .ZN(_19967_));
 AOI21_X2 _47079_ (.A(_15329_),
    .B1(_19349_),
    .B2(_19350_),
    .ZN(_19968_));
 AOI21_X2 _47080_ (.A(_19907_),
    .B1(_19352_),
    .B2(_19353_),
    .ZN(_19969_));
 NOR2_X4 _47081_ (.A1(_19968_),
    .A2(_19969_),
    .ZN(_19970_));
 OAI21_X1 _47082_ (.A(_19967_),
    .B1(_19970_),
    .B2(_19948_),
    .ZN(_05155_));
 NAND2_X1 _47083_ (.A1(_19934_),
    .A2(\icache.lce.lce_cmd_inst.data_r [34]),
    .ZN(_19971_));
 AOI21_X2 _47084_ (.A(_15329_),
    .B1(_19357_),
    .B2(_19358_),
    .ZN(_19972_));
 AOI21_X2 _47085_ (.A(_19907_),
    .B1(_19360_),
    .B2(_19362_),
    .ZN(_19973_));
 NOR2_X4 _47086_ (.A1(_19972_),
    .A2(_19973_),
    .ZN(_19974_));
 OAI21_X1 _47087_ (.A(_19971_),
    .B1(_19974_),
    .B2(_19948_),
    .ZN(_05166_));
 NAND2_X1 _47088_ (.A1(_19934_),
    .A2(\icache.lce.lce_cmd_inst.data_r [35]),
    .ZN(_19975_));
 NOR3_X2 _47089_ (.A1(_19367_),
    .A2(_19368_),
    .A3(_18085_),
    .ZN(_19976_));
 AOI21_X2 _47090_ (.A(_19696_),
    .B1(_19370_),
    .B2(_19372_),
    .ZN(_19977_));
 NOR2_X4 _47091_ (.A1(_19976_),
    .A2(_19977_),
    .ZN(_19978_));
 OAI21_X1 _47092_ (.A(_19975_),
    .B1(_19978_),
    .B2(_19948_),
    .ZN(_05177_));
 BUF_X4 _47093_ (.A(_19635_),
    .Z(_19979_));
 NAND2_X1 _47094_ (.A1(_19979_),
    .A2(\icache.lce.lce_cmd_inst.data_r [36]),
    .ZN(_19980_));
 OAI21_X2 _47095_ (.A(_19963_),
    .B1(_18856_),
    .B2(_18857_),
    .ZN(_19981_));
 NAND3_X2 _47096_ (.A1(_18859_),
    .A2(_18860_),
    .A3(_18470_),
    .ZN(_19982_));
 NAND2_X4 _47097_ (.A1(_19981_),
    .A2(_19982_),
    .ZN(_19983_));
 OAI21_X1 _47098_ (.A(_19980_),
    .B1(_19983_),
    .B2(_19948_),
    .ZN(_05188_));
 NAND2_X1 _47099_ (.A1(_19979_),
    .A2(\icache.lce.lce_cmd_inst.data_r [37]),
    .ZN(_19984_));
 NAND3_X1 _47100_ (.A1(_18864_),
    .A2(_18865_),
    .A3(_15645_),
    .ZN(_19985_));
 NAND3_X1 _47101_ (.A1(_18868_),
    .A2(_19941_),
    .A3(_18869_),
    .ZN(_19986_));
 NAND2_X2 _47102_ (.A1(_19985_),
    .A2(_19986_),
    .ZN(_19987_));
 OAI21_X1 _47103_ (.A(_19984_),
    .B1(_19987_),
    .B2(_19948_),
    .ZN(_05199_));
 NAND2_X1 _47104_ (.A1(_19979_),
    .A2(\icache.lce.lce_cmd_inst.data_r [38]),
    .ZN(_19988_));
 AND3_X1 _47105_ (.A1(_18873_),
    .A2(_18874_),
    .A3(_15503_),
    .ZN(_19989_));
 AOI21_X2 _47106_ (.A(_19907_),
    .B1(_18876_),
    .B2(_18878_),
    .ZN(_19990_));
 NOR2_X4 _47107_ (.A1(_19989_),
    .A2(_19990_),
    .ZN(_19991_));
 BUF_X4 _47108_ (.A(_19649_),
    .Z(_19992_));
 OAI21_X1 _47109_ (.A(_19988_),
    .B1(_19991_),
    .B2(_19992_),
    .ZN(_05210_));
 NAND2_X1 _47110_ (.A1(_19979_),
    .A2(\icache.lce.lce_cmd_inst.data_r [39]),
    .ZN(_19993_));
 AOI21_X2 _47111_ (.A(_15368_),
    .B1(_18691_),
    .B2(_18692_),
    .ZN(_19994_));
 AOI21_X2 _47112_ (.A(_17990_),
    .B1(_18694_),
    .B2(_18695_),
    .ZN(_19995_));
 NOR2_X4 _47113_ (.A1(_19994_),
    .A2(_19995_),
    .ZN(_19996_));
 OAI21_X1 _47114_ (.A(_19993_),
    .B1(_19996_),
    .B2(_19992_),
    .ZN(_05221_));
 NAND2_X1 _47115_ (.A1(_19979_),
    .A2(\icache.lce.lce_cmd_inst.data_r [40]),
    .ZN(_19997_));
 NOR3_X2 _47116_ (.A1(_18699_),
    .A2(_18700_),
    .A3(_18132_),
    .ZN(_19998_));
 AOI21_X2 _47117_ (.A(_19907_),
    .B1(_18702_),
    .B2(_18703_),
    .ZN(_19999_));
 NOR2_X4 _47118_ (.A1(_19998_),
    .A2(_19999_),
    .ZN(_20000_));
 OAI21_X1 _47119_ (.A(_19997_),
    .B1(_20000_),
    .B2(_19992_),
    .ZN(_05233_));
 NAND2_X1 _47120_ (.A1(_19979_),
    .A2(\icache.lce.lce_cmd_inst.data_r [41]),
    .ZN(_20001_));
 NAND2_X1 _47121_ (.A1(_18710_),
    .A2(_19593_),
    .ZN(_20002_));
 OAI21_X2 _47122_ (.A(_19595_),
    .B1(_18712_),
    .B2(_18713_),
    .ZN(_20003_));
 NAND2_X4 _47123_ (.A1(_20002_),
    .A2(_20003_),
    .ZN(_20004_));
 OAI21_X1 _47124_ (.A(_20001_),
    .B1(_20004_),
    .B2(_19992_),
    .ZN(_05244_));
 NAND2_X1 _47125_ (.A1(_19979_),
    .A2(\icache.lce.lce_cmd_inst.data_r [42]),
    .ZN(_20005_));
 NAND3_X2 _47126_ (.A1(_18717_),
    .A2(_18718_),
    .A3(_16143_),
    .ZN(_20006_));
 NAND3_X2 _47127_ (.A1(_18720_),
    .A2(_16237_),
    .A3(_18721_),
    .ZN(_20007_));
 NAND2_X4 _47128_ (.A1(_20006_),
    .A2(_20007_),
    .ZN(_20008_));
 OAI21_X1 _47129_ (.A(_20005_),
    .B1(_20008_),
    .B2(_19992_),
    .ZN(_05255_));
 NAND2_X1 _47130_ (.A1(_19979_),
    .A2(\icache.lce.lce_cmd_inst.data_r [43]),
    .ZN(_20009_));
 AOI21_X2 _47131_ (.A(_15368_),
    .B1(_18725_),
    .B2(_18726_),
    .ZN(_20010_));
 AOI21_X2 _47132_ (.A(_17990_),
    .B1(_18728_),
    .B2(_18729_),
    .ZN(_20011_));
 NOR2_X4 _47133_ (.A1(_20010_),
    .A2(_20011_),
    .ZN(_20012_));
 OAI21_X1 _47134_ (.A(_20009_),
    .B1(_20012_),
    .B2(_19992_),
    .ZN(_05266_));
 NAND2_X1 _47135_ (.A1(_19979_),
    .A2(\icache.lce.lce_cmd_inst.data_r [44]),
    .ZN(_20013_));
 NAND2_X1 _47136_ (.A1(_18735_),
    .A2(_19579_),
    .ZN(_20014_));
 NAND3_X2 _47137_ (.A1(_18737_),
    .A2(_18738_),
    .A3(_16200_),
    .ZN(_20015_));
 NAND2_X4 _47138_ (.A1(_20014_),
    .A2(_20015_),
    .ZN(_20016_));
 OAI21_X1 _47139_ (.A(_20013_),
    .B1(_20016_),
    .B2(_19992_),
    .ZN(_05277_));
 NAND2_X1 _47140_ (.A1(_19979_),
    .A2(\icache.lce.lce_cmd_inst.data_r [45]),
    .ZN(_20017_));
 NAND2_X2 _47141_ (.A1(_18744_),
    .A2(_19579_),
    .ZN(_20018_));
 NAND3_X2 _47142_ (.A1(_18746_),
    .A2(_19941_),
    .A3(_18748_),
    .ZN(_20019_));
 NAND2_X4 _47143_ (.A1(_20018_),
    .A2(_20019_),
    .ZN(_20020_));
 OAI21_X1 _47144_ (.A(_20017_),
    .B1(_20020_),
    .B2(_19992_),
    .ZN(_05288_));
 BUF_X4 _47145_ (.A(_19635_),
    .Z(_20021_));
 NAND2_X1 _47146_ (.A1(_20021_),
    .A2(\icache.lce.lce_cmd_inst.data_r [46]),
    .ZN(_20022_));
 NAND3_X1 _47147_ (.A1(_18752_),
    .A2(_18753_),
    .A3(_15409_),
    .ZN(_20023_));
 OAI21_X1 _47148_ (.A(_19183_),
    .B1(_18755_),
    .B2(_18756_),
    .ZN(_20024_));
 AND2_X4 _47149_ (.A1(_20023_),
    .A2(_20024_),
    .ZN(_20025_));
 OAI21_X1 _47150_ (.A(_20022_),
    .B1(_20025_),
    .B2(_19992_),
    .ZN(_05299_));
 NAND2_X1 _47151_ (.A1(_20021_),
    .A2(\icache.lce.lce_cmd_inst.data_r [47]),
    .ZN(_20026_));
 NAND3_X2 _47152_ (.A1(_18760_),
    .A2(_18762_),
    .A3(_15645_),
    .ZN(_20027_));
 NAND3_X2 _47153_ (.A1(_18764_),
    .A2(_19941_),
    .A3(_18765_),
    .ZN(_20028_));
 NAND2_X4 _47154_ (.A1(_20027_),
    .A2(_20028_),
    .ZN(_20029_));
 OAI21_X1 _47155_ (.A(_20026_),
    .B1(_20029_),
    .B2(_19992_),
    .ZN(_05310_));
 NAND2_X1 _47156_ (.A1(_20021_),
    .A2(\icache.lce.lce_cmd_inst.data_r [48]),
    .ZN(_20030_));
 NAND2_X1 _47157_ (.A1(_18772_),
    .A2(_17634_),
    .ZN(_20031_));
 NAND3_X2 _47158_ (.A1(_18774_),
    .A2(_19941_),
    .A3(_18775_),
    .ZN(_20032_));
 NAND2_X4 _47159_ (.A1(_20031_),
    .A2(_20032_),
    .ZN(_20033_));
 BUF_X4 _47160_ (.A(_19649_),
    .Z(_20034_));
 OAI21_X1 _47161_ (.A(_20030_),
    .B1(_20033_),
    .B2(_20034_),
    .ZN(_05321_));
 NAND2_X1 _47162_ (.A1(_20021_),
    .A2(\icache.lce.lce_cmd_inst.data_r [49]),
    .ZN(_20035_));
 OAI21_X1 _47163_ (.A(_18922_),
    .B1(_18779_),
    .B2(_18780_),
    .ZN(_20036_));
 NAND3_X1 _47164_ (.A1(_18782_),
    .A2(_17415_),
    .A3(_18783_),
    .ZN(_20037_));
 AND2_X4 _47165_ (.A1(_20036_),
    .A2(_20037_),
    .ZN(_20038_));
 OAI21_X1 _47166_ (.A(_20035_),
    .B1(_20038_),
    .B2(_20034_),
    .ZN(_05332_));
 NAND2_X1 _47167_ (.A1(_20021_),
    .A2(\icache.lce.lce_cmd_inst.data_r [50]),
    .ZN(_20039_));
 OAI21_X2 _47168_ (.A(_19366_),
    .B1(_18790_),
    .B2(_18791_),
    .ZN(_20040_));
 OAI21_X2 _47169_ (.A(_15996_),
    .B1(_18787_),
    .B2(_18788_),
    .ZN(_20041_));
 NAND2_X4 _47170_ (.A1(_20040_),
    .A2(_20041_),
    .ZN(_20042_));
 OAI21_X1 _47171_ (.A(_20039_),
    .B1(_20042_),
    .B2(_20034_),
    .ZN(_05344_));
 NAND2_X1 _47172_ (.A1(_20021_),
    .A2(\icache.lce.lce_cmd_inst.data_r [51]),
    .ZN(_20043_));
 OAI21_X1 _47173_ (.A(_19179_),
    .B1(_18796_),
    .B2(_18797_),
    .ZN(_20044_));
 NAND3_X1 _47174_ (.A1(_18799_),
    .A2(_16640_),
    .A3(_18800_),
    .ZN(_20045_));
 AND2_X4 _47175_ (.A1(_20044_),
    .A2(_20045_),
    .ZN(_20046_));
 OAI21_X1 _47176_ (.A(_20043_),
    .B1(_20046_),
    .B2(_20034_),
    .ZN(_05347_));
 NAND2_X1 _47177_ (.A1(_20021_),
    .A2(\icache.lce.lce_cmd_inst.data_r [52]),
    .ZN(_20047_));
 AND3_X1 _47178_ (.A1(_18804_),
    .A2(_15621_),
    .A3(_18806_),
    .ZN(_20048_));
 AOI21_X2 _47179_ (.A(_17990_),
    .B1(_18808_),
    .B2(_18810_),
    .ZN(_20049_));
 NOR2_X4 _47180_ (.A1(_20048_),
    .A2(_20049_),
    .ZN(_20050_));
 OAI21_X1 _47181_ (.A(_20047_),
    .B1(_20050_),
    .B2(_20034_),
    .ZN(_05348_));
 NAND2_X1 _47182_ (.A1(_20021_),
    .A2(\icache.lce.lce_cmd_inst.data_r [53]),
    .ZN(_20051_));
 OR3_X2 _47183_ (.A1(_18814_),
    .A2(_15644_),
    .A3(_18815_),
    .ZN(_20052_));
 NAND2_X1 _47184_ (.A1(_18819_),
    .A2(_17567_),
    .ZN(_20053_));
 NAND2_X4 _47185_ (.A1(_20052_),
    .A2(_20053_),
    .ZN(_20054_));
 OAI21_X1 _47186_ (.A(_20051_),
    .B1(_20054_),
    .B2(_20034_),
    .ZN(_05349_));
 NAND2_X1 _47187_ (.A1(_20021_),
    .A2(\icache.lce.lce_cmd_inst.data_r [54]),
    .ZN(_20055_));
 AOI21_X1 _47188_ (.A(_15724_),
    .B1(_18823_),
    .B2(_18824_),
    .ZN(_20056_));
 AND3_X1 _47189_ (.A1(_18826_),
    .A2(_15430_),
    .A3(_18827_),
    .ZN(_20057_));
 OR2_X4 _47190_ (.A1(_20056_),
    .A2(_20057_),
    .ZN(_20058_));
 OAI21_X1 _47191_ (.A(_20055_),
    .B1(_20058_),
    .B2(_20034_),
    .ZN(_05350_));
 NAND2_X1 _47192_ (.A1(_20021_),
    .A2(\icache.lce.lce_cmd_inst.data_r [55]),
    .ZN(_20059_));
 AOI21_X1 _47193_ (.A(_15329_),
    .B1(_18831_),
    .B2(_18832_),
    .ZN(_20060_));
 AOI21_X1 _47194_ (.A(_19907_),
    .B1(_18834_),
    .B2(_18835_),
    .ZN(_20061_));
 NOR2_X2 _47195_ (.A1(_20060_),
    .A2(_20061_),
    .ZN(_20062_));
 OAI21_X1 _47196_ (.A(_20059_),
    .B1(_20062_),
    .B2(_20034_),
    .ZN(_05351_));
 BUF_X16 _47197_ (.A(_15302_),
    .Z(_20063_));
 NAND2_X1 _47198_ (.A1(_20063_),
    .A2(\icache.lce.lce_cmd_inst.data_r [56]),
    .ZN(_20064_));
 AOI21_X1 _47199_ (.A(_16406_),
    .B1(_18839_),
    .B2(_18840_),
    .ZN(_20065_));
 AND3_X1 _47200_ (.A1(_18842_),
    .A2(_18843_),
    .A3(_15367_),
    .ZN(_20066_));
 OR2_X4 _47201_ (.A1(_20065_),
    .A2(_20066_),
    .ZN(_20067_));
 OAI21_X1 _47202_ (.A(_20064_),
    .B1(_20067_),
    .B2(_20034_),
    .ZN(_05352_));
 NAND2_X1 _47203_ (.A1(_20063_),
    .A2(\icache.lce.lce_cmd_inst.data_r [57]),
    .ZN(_20068_));
 OAI21_X1 _47204_ (.A(_18922_),
    .B1(_18847_),
    .B2(_18848_),
    .ZN(_20069_));
 NAND3_X1 _47205_ (.A1(_18850_),
    .A2(_18851_),
    .A3(_15849_),
    .ZN(_20070_));
 AND2_X4 _47206_ (.A1(_20069_),
    .A2(_20070_),
    .ZN(_20071_));
 OAI21_X1 _47207_ (.A(_20068_),
    .B1(_20071_),
    .B2(_20034_),
    .ZN(_05353_));
 NAND2_X1 _47208_ (.A1(_20063_),
    .A2(\icache.lce.lce_cmd_inst.data_r [58]),
    .ZN(_20072_));
 NAND3_X1 _47209_ (.A1(_17949_),
    .A2(_17950_),
    .A3(_15834_),
    .ZN(_20073_));
 OAI21_X1 _47210_ (.A(_18366_),
    .B1(_17952_),
    .B2(_17953_),
    .ZN(_20074_));
 AND2_X4 _47211_ (.A1(_20073_),
    .A2(_20074_),
    .ZN(_20075_));
 BUF_X16 _47212_ (.A(_15601_),
    .Z(_20076_));
 OAI21_X1 _47213_ (.A(_20072_),
    .B1(_20075_),
    .B2(_20076_),
    .ZN(_05354_));
 NAND2_X1 _47214_ (.A1(_20063_),
    .A2(\icache.lce.lce_cmd_inst.data_r [59]),
    .ZN(_20077_));
 NAND2_X1 _47215_ (.A1(_17959_),
    .A2(_17634_),
    .ZN(_20078_));
 NAND2_X1 _47216_ (.A1(_17964_),
    .A2(_15905_),
    .ZN(_20079_));
 NAND2_X2 _47217_ (.A1(_20078_),
    .A2(_20079_),
    .ZN(_20080_));
 OAI21_X1 _47218_ (.A(_20077_),
    .B1(_20080_),
    .B2(_20076_),
    .ZN(_05355_));
 NAND2_X1 _47219_ (.A1(_20063_),
    .A2(\icache.lce.lce_cmd_inst.data_r [60]),
    .ZN(_20081_));
 OAI21_X1 _47220_ (.A(_19963_),
    .B1(_17972_),
    .B2(_17973_),
    .ZN(_20082_));
 OAI21_X1 _47221_ (.A(_19951_),
    .B1(_17968_),
    .B2(_17969_),
    .ZN(_20083_));
 NAND2_X2 _47222_ (.A1(_20082_),
    .A2(_20083_),
    .ZN(_20084_));
 OAI21_X1 _47223_ (.A(_20081_),
    .B1(_20084_),
    .B2(_20076_),
    .ZN(_05357_));
 NAND2_X1 _47224_ (.A1(_20063_),
    .A2(\icache.lce.lce_cmd_inst.data_r [61]),
    .ZN(_20085_));
 NAND2_X1 _47225_ (.A1(_17979_),
    .A2(_17634_),
    .ZN(_20086_));
 OAI21_X1 _47226_ (.A(_19951_),
    .B1(_17982_),
    .B2(_17983_),
    .ZN(_20087_));
 NAND2_X2 _47227_ (.A1(_20086_),
    .A2(_20087_),
    .ZN(_20088_));
 OAI21_X1 _47228_ (.A(_20085_),
    .B1(_20088_),
    .B2(_20076_),
    .ZN(_05358_));
 NAND2_X1 _47229_ (.A1(_20063_),
    .A2(\icache.lce.lce_cmd_inst.data_r [62]),
    .ZN(_20089_));
 OAI21_X1 _47230_ (.A(_19963_),
    .B1(_17987_),
    .B2(_17989_),
    .ZN(_20090_));
 NAND3_X1 _47231_ (.A1(_17992_),
    .A2(_19941_),
    .A3(_17993_),
    .ZN(_20091_));
 NAND2_X2 _47232_ (.A1(_20090_),
    .A2(_20091_),
    .ZN(_20092_));
 OAI21_X1 _47233_ (.A(_20089_),
    .B1(_20092_),
    .B2(_20076_),
    .ZN(_05359_));
 NAND2_X1 _47234_ (.A1(_20063_),
    .A2(\icache.lce.lce_cmd_inst.data_r [63]),
    .ZN(_20093_));
 OR3_X2 _47235_ (.A1(_17997_),
    .A2(_16012_),
    .A3(_17998_),
    .ZN(_20094_));
 OAI21_X2 _47236_ (.A(_19951_),
    .B1(_18000_),
    .B2(_18001_),
    .ZN(_20095_));
 NAND2_X4 _47237_ (.A1(_20094_),
    .A2(_20095_),
    .ZN(_20096_));
 OAI21_X1 _47238_ (.A(_20093_),
    .B1(_20096_),
    .B2(_20076_),
    .ZN(_05360_));
 NAND2_X1 _47239_ (.A1(_20063_),
    .A2(\icache.lce.lce_cmd_inst.data_r [64]),
    .ZN(_20097_));
 OAI21_X2 _47240_ (.A(_15834_),
    .B1(_18007_),
    .B2(_18008_),
    .ZN(_20098_));
 OR3_X1 _47241_ (.A1(_18010_),
    .A2(_18011_),
    .A3(_15314_),
    .ZN(_20099_));
 AND2_X4 _47242_ (.A1(_20098_),
    .A2(_20099_),
    .ZN(_20100_));
 OAI21_X1 _47243_ (.A(_20097_),
    .B1(_20100_),
    .B2(_20076_),
    .ZN(_05361_));
 NAND2_X1 _47244_ (.A1(_20063_),
    .A2(\icache.lce.lce_cmd_inst.data_r [65]),
    .ZN(_20101_));
 AND3_X1 _47245_ (.A1(_18015_),
    .A2(_18016_),
    .A3(_15503_),
    .ZN(_20102_));
 AOI21_X2 _47246_ (.A(_19907_),
    .B1(_18018_),
    .B2(_18021_),
    .ZN(_20103_));
 NOR2_X4 _47247_ (.A1(_20102_),
    .A2(_20103_),
    .ZN(_20104_));
 OAI21_X1 _47248_ (.A(_20101_),
    .B1(_20104_),
    .B2(_20076_),
    .ZN(_05362_));
 BUF_X4 _47249_ (.A(_15302_),
    .Z(_20105_));
 NAND2_X1 _47250_ (.A1(_20105_),
    .A2(\icache.lce.lce_cmd_inst.data_r [66]),
    .ZN(_20106_));
 NOR3_X1 _47251_ (.A1(_18025_),
    .A2(_18026_),
    .A3(_18085_),
    .ZN(_20107_));
 AOI21_X1 _47252_ (.A(_17990_),
    .B1(_18028_),
    .B2(_18030_),
    .ZN(_20108_));
 NOR2_X2 _47253_ (.A1(_20107_),
    .A2(_20108_),
    .ZN(_20109_));
 OAI21_X1 _47254_ (.A(_20106_),
    .B1(_20109_),
    .B2(_20076_),
    .ZN(_05363_));
 NAND2_X1 _47255_ (.A1(_20105_),
    .A2(\icache.lce.lce_cmd_inst.data_r [67]),
    .ZN(_20110_));
 AOI21_X2 _47256_ (.A(_16406_),
    .B1(_18035_),
    .B2(_18036_),
    .ZN(_20111_));
 AND3_X1 _47257_ (.A1(_18038_),
    .A2(_15819_),
    .A3(_18039_),
    .ZN(_20112_));
 OR2_X2 _47258_ (.A1(_20111_),
    .A2(_20112_),
    .ZN(_20113_));
 OAI21_X1 _47259_ (.A(_20110_),
    .B1(_20113_),
    .B2(_20076_),
    .ZN(_05364_));
 NAND2_X1 _47260_ (.A1(_20105_),
    .A2(\icache.lce.lce_cmd_inst.data_r [68]),
    .ZN(_20114_));
 OAI21_X1 _47261_ (.A(_19963_),
    .B1(_18043_),
    .B2(_18044_),
    .ZN(_20115_));
 OAI21_X1 _47262_ (.A(_19951_),
    .B1(_18046_),
    .B2(_18047_),
    .ZN(_20116_));
 NAND2_X2 _47263_ (.A1(_20115_),
    .A2(_20116_),
    .ZN(_20117_));
 BUF_X8 _47264_ (.A(_15601_),
    .Z(_20118_));
 OAI21_X1 _47265_ (.A(_20114_),
    .B1(_20117_),
    .B2(_20118_),
    .ZN(_05365_));
 NAND2_X1 _47266_ (.A1(_20105_),
    .A2(\icache.lce.lce_cmd_inst.data_r [69]),
    .ZN(_20119_));
 AND3_X1 _47267_ (.A1(_18051_),
    .A2(_15621_),
    .A3(_18052_),
    .ZN(_20120_));
 AOI21_X1 _47268_ (.A(_17990_),
    .B1(_18054_),
    .B2(_18055_),
    .ZN(_20121_));
 NOR2_X2 _47269_ (.A1(_20120_),
    .A2(_20121_),
    .ZN(_20122_));
 OAI21_X1 _47270_ (.A(_20119_),
    .B1(_20122_),
    .B2(_20118_),
    .ZN(_05366_));
 NAND2_X1 _47271_ (.A1(_20105_),
    .A2(\icache.lce.lce_cmd_inst.data_r [70]),
    .ZN(_20123_));
 AOI21_X4 _47272_ (.A(_15368_),
    .B1(_18059_),
    .B2(_18060_),
    .ZN(_20124_));
 AOI21_X1 _47273_ (.A(_17990_),
    .B1(_18062_),
    .B2(_18063_),
    .ZN(_20125_));
 NOR2_X2 _47274_ (.A1(_20124_),
    .A2(_20125_),
    .ZN(_20126_));
 OAI21_X1 _47275_ (.A(_20123_),
    .B1(_20126_),
    .B2(_20118_),
    .ZN(_05368_));
 NAND2_X1 _47276_ (.A1(_20105_),
    .A2(\icache.lce.lce_cmd_inst.data_r [71]),
    .ZN(_20127_));
 OAI21_X1 _47277_ (.A(_19963_),
    .B1(_18067_),
    .B2(_18068_),
    .ZN(_20128_));
 OAI21_X1 _47278_ (.A(_19951_),
    .B1(_18070_),
    .B2(_18071_),
    .ZN(_20129_));
 NAND2_X2 _47279_ (.A1(_20128_),
    .A2(_20129_),
    .ZN(_20130_));
 OAI21_X1 _47280_ (.A(_20127_),
    .B1(_20130_),
    .B2(_20118_),
    .ZN(_05369_));
 NAND2_X1 _47281_ (.A1(_20105_),
    .A2(\icache.lce.lce_cmd_inst.data_r [72]),
    .ZN(_20131_));
 OAI21_X2 _47282_ (.A(_19963_),
    .B1(_18075_),
    .B2(_18076_),
    .ZN(_20132_));
 NAND3_X2 _47283_ (.A1(_18078_),
    .A2(_19941_),
    .A3(_18079_),
    .ZN(_20133_));
 NAND2_X4 _47284_ (.A1(_20132_),
    .A2(_20133_),
    .ZN(_20134_));
 OAI21_X1 _47285_ (.A(_20131_),
    .B1(_20134_),
    .B2(_20118_),
    .ZN(_05370_));
 NAND2_X1 _47286_ (.A1(_20105_),
    .A2(\icache.lce.lce_cmd_inst.data_r [73]),
    .ZN(_20135_));
 OAI21_X1 _47287_ (.A(_19366_),
    .B1(_18083_),
    .B2(_18084_),
    .ZN(_20136_));
 NAND3_X1 _47288_ (.A1(_18087_),
    .A2(_18088_),
    .A3(_15354_),
    .ZN(_20137_));
 NAND2_X2 _47289_ (.A1(_20136_),
    .A2(_20137_),
    .ZN(_20138_));
 OAI21_X1 _47290_ (.A(_20135_),
    .B1(_20138_),
    .B2(_20118_),
    .ZN(_05371_));
 NAND2_X1 _47291_ (.A1(_20105_),
    .A2(\icache.lce.lce_cmd_inst.data_r [74]),
    .ZN(_20139_));
 NAND2_X1 _47292_ (.A1(_18095_),
    .A2(_19593_),
    .ZN(_20140_));
 OAI21_X2 _47293_ (.A(_15996_),
    .B1(_18097_),
    .B2(_18098_),
    .ZN(_20141_));
 NAND2_X4 _47294_ (.A1(_20140_),
    .A2(_20141_),
    .ZN(_20142_));
 OAI21_X1 _47295_ (.A(_20139_),
    .B1(_20142_),
    .B2(_20118_),
    .ZN(_05372_));
 NAND2_X1 _47296_ (.A1(_20105_),
    .A2(\icache.lce.lce_cmd_inst.data_r [75]),
    .ZN(_20143_));
 NOR3_X1 _47297_ (.A1(_18102_),
    .A2(_18103_),
    .A3(_18132_),
    .ZN(_20144_));
 AOI21_X4 _47298_ (.A(_19907_),
    .B1(_18105_),
    .B2(_18107_),
    .ZN(_20145_));
 NOR2_X2 _47299_ (.A1(_20144_),
    .A2(_20145_),
    .ZN(_20146_));
 OAI21_X1 _47300_ (.A(_20143_),
    .B1(_20146_),
    .B2(_20118_),
    .ZN(_05373_));
 BUF_X4 _47301_ (.A(_15302_),
    .Z(_20147_));
 NAND2_X1 _47302_ (.A1(_20147_),
    .A2(\icache.lce.lce_cmd_inst.data_r [76]),
    .ZN(_20148_));
 OAI21_X1 _47303_ (.A(_16143_),
    .B1(_18111_),
    .B2(_18112_),
    .ZN(_20149_));
 NAND3_X1 _47304_ (.A1(_18114_),
    .A2(_16237_),
    .A3(_18117_),
    .ZN(_20150_));
 NAND2_X2 _47305_ (.A1(_20149_),
    .A2(_20150_),
    .ZN(_20151_));
 OAI21_X1 _47306_ (.A(_20148_),
    .B1(_20151_),
    .B2(_20118_),
    .ZN(_05374_));
 NAND2_X1 _47307_ (.A1(_20147_),
    .A2(\icache.lce.lce_cmd_inst.data_r [77]),
    .ZN(_20152_));
 OAI21_X1 _47308_ (.A(_16143_),
    .B1(_18122_),
    .B2(_18123_),
    .ZN(_20153_));
 NAND3_X1 _47309_ (.A1(_18125_),
    .A2(_16237_),
    .A3(_18126_),
    .ZN(_20154_));
 NAND2_X2 _47310_ (.A1(_20153_),
    .A2(_20154_),
    .ZN(_20155_));
 OAI21_X1 _47311_ (.A(_20152_),
    .B1(_20155_),
    .B2(_20118_),
    .ZN(_05375_));
 NAND2_X1 _47312_ (.A1(_20147_),
    .A2(\icache.lce.lce_cmd_inst.data_r [78]),
    .ZN(_20156_));
 NOR3_X2 _47313_ (.A1(_18130_),
    .A2(_18131_),
    .A3(_18085_),
    .ZN(_20157_));
 AOI21_X2 _47314_ (.A(_17990_),
    .B1(_18134_),
    .B2(_18135_),
    .ZN(_20158_));
 NOR2_X4 _47315_ (.A1(_20157_),
    .A2(_20158_),
    .ZN(_20159_));
 BUF_X4 _47316_ (.A(_15601_),
    .Z(_20160_));
 OAI21_X1 _47317_ (.A(_20156_),
    .B1(_20159_),
    .B2(_20160_),
    .ZN(_05376_));
 NAND2_X1 _47318_ (.A1(_20147_),
    .A2(\icache.lce.lce_cmd_inst.data_r [79]),
    .ZN(_20161_));
 AND3_X1 _47319_ (.A1(_18139_),
    .A2(_18140_),
    .A3(_15503_),
    .ZN(_20162_));
 AOI21_X1 _47320_ (.A(_19907_),
    .B1(_18142_),
    .B2(_18143_),
    .ZN(_20163_));
 NOR2_X2 _47321_ (.A1(_20162_),
    .A2(_20163_),
    .ZN(_20164_));
 OAI21_X1 _47322_ (.A(_20161_),
    .B1(_20164_),
    .B2(_20160_),
    .ZN(_05377_));
 NAND2_X1 _47323_ (.A1(_20147_),
    .A2(\icache.lce.lce_cmd_inst.data_r [80]),
    .ZN(_20165_));
 OAI21_X2 _47324_ (.A(_19963_),
    .B1(_18147_),
    .B2(_18148_),
    .ZN(_20166_));
 OAI21_X2 _47325_ (.A(_19951_),
    .B1(_18150_),
    .B2(_18151_),
    .ZN(_20167_));
 NAND2_X4 _47326_ (.A1(_20166_),
    .A2(_20167_),
    .ZN(_20168_));
 OAI21_X1 _47327_ (.A(_20165_),
    .B1(_20168_),
    .B2(_20160_),
    .ZN(_05379_));
 NAND2_X1 _47328_ (.A1(_20147_),
    .A2(\icache.lce.lce_cmd_inst.data_r [81]),
    .ZN(_20169_));
 AOI21_X2 _47329_ (.A(_15724_),
    .B1(_18155_),
    .B2(_18156_),
    .ZN(_20170_));
 AND3_X1 _47330_ (.A1(_18158_),
    .A2(_15430_),
    .A3(_18159_),
    .ZN(_20171_));
 OR2_X4 _47331_ (.A1(_20170_),
    .A2(_20171_),
    .ZN(_20172_));
 OAI21_X1 _47332_ (.A(_20169_),
    .B1(_20172_),
    .B2(_20160_),
    .ZN(_05380_));
 NAND2_X1 _47333_ (.A1(_20147_),
    .A2(\icache.lce.lce_cmd_inst.data_r [82]),
    .ZN(_20173_));
 OAI21_X2 _47334_ (.A(_19963_),
    .B1(_18163_),
    .B2(_18165_),
    .ZN(_20174_));
 NAND3_X2 _47335_ (.A1(_18167_),
    .A2(_19941_),
    .A3(_18168_),
    .ZN(_20175_));
 NAND2_X4 _47336_ (.A1(_20174_),
    .A2(_20175_),
    .ZN(_20176_));
 OAI21_X1 _47337_ (.A(_20173_),
    .B1(_20176_),
    .B2(_20160_),
    .ZN(_05381_));
 NAND2_X1 _47338_ (.A1(_20147_),
    .A2(\icache.lce.lce_cmd_inst.data_r [83]),
    .ZN(_20177_));
 OAI21_X1 _47339_ (.A(_16143_),
    .B1(_18172_),
    .B2(_18173_),
    .ZN(_20178_));
 OAI21_X1 _47340_ (.A(_15996_),
    .B1(_18175_),
    .B2(_18176_),
    .ZN(_20179_));
 NAND2_X2 _47341_ (.A1(_20178_),
    .A2(_20179_),
    .ZN(_20180_));
 OAI21_X1 _47342_ (.A(_20177_),
    .B1(_20180_),
    .B2(_20160_),
    .ZN(_05382_));
 NAND2_X1 _47343_ (.A1(_20147_),
    .A2(\icache.lce.lce_cmd_inst.data_r [84]),
    .ZN(_20181_));
 AND3_X1 _47344_ (.A1(_18184_),
    .A2(_15522_),
    .A3(_18186_),
    .ZN(_20182_));
 AOI21_X1 _47345_ (.A(_18419_),
    .B1(_18181_),
    .B2(_18182_),
    .ZN(_20183_));
 OR2_X4 _47346_ (.A1(_20182_),
    .A2(_20183_),
    .ZN(_20184_));
 OAI21_X1 _47347_ (.A(_20181_),
    .B1(_20184_),
    .B2(_20160_),
    .ZN(_05383_));
 NAND2_X1 _47348_ (.A1(_20147_),
    .A2(\icache.lce.lce_cmd_inst.data_r [85]),
    .ZN(_20185_));
 NAND2_X1 _47349_ (.A1(_18192_),
    .A2(_17634_),
    .ZN(_20186_));
 NAND3_X1 _47350_ (.A1(_18194_),
    .A2(_19941_),
    .A3(_18195_),
    .ZN(_20187_));
 NAND2_X2 _47351_ (.A1(_20186_),
    .A2(_20187_),
    .ZN(_20188_));
 OAI21_X1 _47352_ (.A(_20185_),
    .B1(_20188_),
    .B2(_20160_),
    .ZN(_05384_));
 BUF_X4 _47353_ (.A(_15302_),
    .Z(_20189_));
 NAND2_X1 _47354_ (.A1(_20189_),
    .A2(\icache.lce.lce_cmd_inst.data_r [86]),
    .ZN(_20190_));
 NAND3_X1 _47355_ (.A1(_18199_),
    .A2(_18200_),
    .A3(_16143_),
    .ZN(_20191_));
 NAND3_X1 _47356_ (.A1(_18202_),
    .A2(_18203_),
    .A3(_15354_),
    .ZN(_20192_));
 NAND2_X2 _47357_ (.A1(_20191_),
    .A2(_20192_),
    .ZN(_20193_));
 OAI21_X1 _47358_ (.A(_20190_),
    .B1(_20193_),
    .B2(_20160_),
    .ZN(_05385_));
 NAND2_X1 _47359_ (.A1(_20189_),
    .A2(\icache.lce.lce_cmd_inst.data_r [87]),
    .ZN(_20194_));
 NAND2_X1 _47360_ (.A1(_18211_),
    .A2(_17634_),
    .ZN(_20195_));
 OAI21_X1 _47361_ (.A(_19951_),
    .B1(_18213_),
    .B2(_18214_),
    .ZN(_20196_));
 NAND2_X2 _47362_ (.A1(_20195_),
    .A2(_20196_),
    .ZN(_20197_));
 OAI21_X1 _47363_ (.A(_20194_),
    .B1(_20197_),
    .B2(_20160_),
    .ZN(_05386_));
 NAND2_X1 _47364_ (.A1(_20189_),
    .A2(\icache.lce.lce_cmd_inst.data_r [88]),
    .ZN(_20198_));
 OAI21_X1 _47365_ (.A(_19963_),
    .B1(_18218_),
    .B2(_18219_),
    .ZN(_20199_));
 NAND3_X1 _47366_ (.A1(_18221_),
    .A2(_18222_),
    .A3(_16200_),
    .ZN(_20200_));
 NAND2_X2 _47367_ (.A1(_20199_),
    .A2(_20200_),
    .ZN(_20201_));
 BUF_X8 _47368_ (.A(_15601_),
    .Z(_20202_));
 OAI21_X1 _47369_ (.A(_20198_),
    .B1(_20201_),
    .B2(_20202_),
    .ZN(_05387_));
 NAND2_X1 _47370_ (.A1(_20189_),
    .A2(\icache.lce.lce_cmd_inst.data_r [89]),
    .ZN(_20203_));
 NAND2_X1 _47371_ (.A1(_18228_),
    .A2(_17634_),
    .ZN(_20204_));
 NAND3_X2 _47372_ (.A1(_18230_),
    .A2(_19941_),
    .A3(_18231_),
    .ZN(_20205_));
 NAND2_X4 _47373_ (.A1(_20204_),
    .A2(_20205_),
    .ZN(_20206_));
 OAI21_X1 _47374_ (.A(_20203_),
    .B1(_20206_),
    .B2(_20202_),
    .ZN(_05388_));
 NAND2_X1 _47375_ (.A1(_20189_),
    .A2(\icache.lce.lce_cmd_inst.data_r [90]),
    .ZN(_20207_));
 NAND2_X1 _47376_ (.A1(_18237_),
    .A2(_15598_),
    .ZN(_20208_));
 NAND3_X1 _47377_ (.A1(_18239_),
    .A2(_16237_),
    .A3(_18241_),
    .ZN(_20209_));
 NAND2_X2 _47378_ (.A1(_20208_),
    .A2(_20209_),
    .ZN(_20210_));
 OAI21_X1 _47379_ (.A(_20207_),
    .B1(_20210_),
    .B2(_20202_),
    .ZN(_05390_));
 NAND2_X1 _47380_ (.A1(_20189_),
    .A2(\icache.lce.lce_cmd_inst.data_r [91]),
    .ZN(_20211_));
 OAI21_X1 _47381_ (.A(_15645_),
    .B1(_18245_),
    .B2(_18246_),
    .ZN(_20212_));
 NAND3_X1 _47382_ (.A1(_18248_),
    .A2(_16013_),
    .A3(_18249_),
    .ZN(_20213_));
 NAND2_X2 _47383_ (.A1(_20212_),
    .A2(_20213_),
    .ZN(_20214_));
 OAI21_X1 _47384_ (.A(_20211_),
    .B1(_20214_),
    .B2(_20202_),
    .ZN(_05391_));
 NAND2_X1 _47385_ (.A1(_20189_),
    .A2(\icache.lce.lce_cmd_inst.data_r [92]),
    .ZN(_20215_));
 AOI21_X1 _47386_ (.A(_15329_),
    .B1(_18253_),
    .B2(_18254_),
    .ZN(_20216_));
 AOI21_X1 _47387_ (.A(_18085_),
    .B1(_18256_),
    .B2(_18257_),
    .ZN(_20217_));
 NOR2_X2 _47388_ (.A1(_20216_),
    .A2(_20217_),
    .ZN(_20218_));
 OAI21_X1 _47389_ (.A(_20215_),
    .B1(_20218_),
    .B2(_20202_),
    .ZN(_05392_));
 NAND2_X1 _47390_ (.A1(_20189_),
    .A2(\icache.lce.lce_cmd_inst.data_r [93]),
    .ZN(_20219_));
 OAI21_X1 _47391_ (.A(_15834_),
    .B1(_18261_),
    .B2(_18262_),
    .ZN(_20220_));
 NAND3_X1 _47392_ (.A1(_18264_),
    .A2(_18265_),
    .A3(_15849_),
    .ZN(_20221_));
 AND2_X4 _47393_ (.A1(_20220_),
    .A2(_20221_),
    .ZN(_20222_));
 OAI21_X1 _47394_ (.A(_20219_),
    .B1(_20222_),
    .B2(_20202_),
    .ZN(_05393_));
 NAND2_X1 _47395_ (.A1(_20189_),
    .A2(\icache.lce.lce_cmd_inst.data_r [4]),
    .ZN(_20223_));
 NOR3_X2 _47396_ (.A1(_19094_),
    .A2(_19095_),
    .A3(_18132_),
    .ZN(_20224_));
 AOI21_X2 _47397_ (.A(_18085_),
    .B1(_19097_),
    .B2(_19099_),
    .ZN(_20225_));
 NOR2_X4 _47398_ (.A1(_20224_),
    .A2(_20225_),
    .ZN(_20226_));
 OAI21_X1 _47399_ (.A(_20223_),
    .B1(_20226_),
    .B2(_20202_),
    .ZN(_05333_));
 NAND2_X1 _47400_ (.A1(_20189_),
    .A2(\icache.lce.lce_cmd_inst.data_r [5]),
    .ZN(_20227_));
 NAND3_X1 _47401_ (.A1(_19103_),
    .A2(_16360_),
    .A3(_19104_),
    .ZN(_20228_));
 OAI21_X1 _47402_ (.A(_19183_),
    .B1(_19106_),
    .B2(_19107_),
    .ZN(_20229_));
 AND2_X4 _47403_ (.A1(_20228_),
    .A2(_20229_),
    .ZN(_20230_));
 OAI21_X1 _47404_ (.A(_20227_),
    .B1(_20230_),
    .B2(_20202_),
    .ZN(_05356_));
 BUF_X8 _47405_ (.A(_15302_),
    .Z(_20231_));
 NAND2_X1 _47406_ (.A1(_20231_),
    .A2(\icache.lce.lce_cmd_inst.data_r [6]),
    .ZN(_20232_));
 OAI21_X1 _47407_ (.A(_19179_),
    .B1(_19112_),
    .B2(_19113_),
    .ZN(_20233_));
 OAI21_X1 _47408_ (.A(_15315_),
    .B1(_19115_),
    .B2(_19116_),
    .ZN(_20234_));
 AND2_X4 _47409_ (.A1(_20233_),
    .A2(_20234_),
    .ZN(_20235_));
 OAI21_X1 _47410_ (.A(_20232_),
    .B1(_20235_),
    .B2(_20202_),
    .ZN(_05367_));
 NAND2_X1 _47411_ (.A1(_20231_),
    .A2(\icache.lce.lce_cmd_inst.data_r [7]),
    .ZN(_20236_));
 NAND2_X1 _47412_ (.A1(_19122_),
    .A2(_17634_),
    .ZN(_20237_));
 OAI21_X1 _47413_ (.A(_15656_),
    .B1(_19124_),
    .B2(_19125_),
    .ZN(_20238_));
 NAND2_X2 _47414_ (.A1(_20237_),
    .A2(_20238_),
    .ZN(_20239_));
 OAI21_X1 _47415_ (.A(_20236_),
    .B1(_20239_),
    .B2(_20202_),
    .ZN(_05378_));
 NAND2_X1 _47416_ (.A1(_20231_),
    .A2(\icache.lce.lce_cmd_inst.data_r [8]),
    .ZN(_20240_));
 OAI21_X1 _47417_ (.A(_15834_),
    .B1(_19129_),
    .B2(_19130_),
    .ZN(_20241_));
 OAI21_X1 _47418_ (.A(_18366_),
    .B1(_19132_),
    .B2(_19133_),
    .ZN(_20242_));
 AND2_X4 _47419_ (.A1(_20241_),
    .A2(_20242_),
    .ZN(_20243_));
 BUF_X8 _47420_ (.A(_15601_),
    .Z(_20244_));
 OAI21_X1 _47421_ (.A(_20240_),
    .B1(_20243_),
    .B2(_20244_),
    .ZN(_05389_));
 NAND2_X1 _47422_ (.A1(_20231_),
    .A2(\icache.lce.lce_cmd_inst.data_r [9]),
    .ZN(_20245_));
 AOI21_X2 _47423_ (.A(_15368_),
    .B1(_19138_),
    .B2(_19139_),
    .ZN(_20246_));
 AOI21_X1 _47424_ (.A(_17990_),
    .B1(_19141_),
    .B2(_19142_),
    .ZN(_20247_));
 NOR2_X2 _47425_ (.A1(_20246_),
    .A2(_20247_),
    .ZN(_20248_));
 OAI21_X1 _47426_ (.A(_20245_),
    .B1(_20248_),
    .B2(_20244_),
    .ZN(_05400_));
 NAND2_X1 _47427_ (.A1(_20231_),
    .A2(\icache.lce.lce_cmd_inst.data_r [10]),
    .ZN(_20249_));
 OAI21_X2 _47428_ (.A(_15645_),
    .B1(_19146_),
    .B2(_19147_),
    .ZN(_20250_));
 OAI21_X2 _47429_ (.A(_15656_),
    .B1(_19149_),
    .B2(_19150_),
    .ZN(_20251_));
 NAND2_X4 _47430_ (.A1(_20250_),
    .A2(_20251_),
    .ZN(_20252_));
 OAI21_X1 _47431_ (.A(_20249_),
    .B1(_20252_),
    .B2(_20244_),
    .ZN(_04900_));
 NAND2_X1 _47432_ (.A1(_20231_),
    .A2(\icache.lce.lce_cmd_inst.data_r [11]),
    .ZN(_20253_));
 NOR2_X1 _47433_ (.A1(_19156_),
    .A2(_15354_),
    .ZN(_20254_));
 AOI21_X2 _47434_ (.A(_18085_),
    .B1(_19158_),
    .B2(_19159_),
    .ZN(_20255_));
 NOR2_X4 _47435_ (.A1(_20254_),
    .A2(_20255_),
    .ZN(_20256_));
 OAI21_X1 _47436_ (.A(_20253_),
    .B1(_20256_),
    .B2(_20244_),
    .ZN(_04911_));
 NAND2_X1 _47437_ (.A1(_20231_),
    .A2(\icache.lce.lce_cmd_inst.data_r [12]),
    .ZN(_20257_));
 NAND3_X1 _47438_ (.A1(_19163_),
    .A2(_16438_),
    .A3(_19164_),
    .ZN(_20258_));
 OAI21_X1 _47439_ (.A(_18366_),
    .B1(_19166_),
    .B2(_19167_),
    .ZN(_20259_));
 AND2_X4 _47440_ (.A1(_20258_),
    .A2(_20259_),
    .ZN(_20260_));
 OAI21_X1 _47441_ (.A(_20257_),
    .B1(_20260_),
    .B2(_20244_),
    .ZN(_04922_));
 NAND2_X1 _47442_ (.A1(_20231_),
    .A2(\icache.lce.lce_cmd_inst.data_r [13]),
    .ZN(_20261_));
 NAND3_X1 _47443_ (.A1(_19171_),
    .A2(_19172_),
    .A3(_16372_),
    .ZN(_20262_));
 NAND3_X1 _47444_ (.A1(_19174_),
    .A2(_17415_),
    .A3(_19175_),
    .ZN(_20263_));
 AND2_X4 _47445_ (.A1(_20262_),
    .A2(_20263_),
    .ZN(_20264_));
 OAI21_X1 _47446_ (.A(_20261_),
    .B1(_20264_),
    .B2(_20244_),
    .ZN(_04933_));
 NAND2_X1 _47447_ (.A1(_20231_),
    .A2(\icache.lce.lce_cmd_inst.data_r [14]),
    .ZN(_20265_));
 OAI21_X1 _47448_ (.A(_15834_),
    .B1(_19180_),
    .B2(_19181_),
    .ZN(_20266_));
 OAI21_X1 _47449_ (.A(_15849_),
    .B1(_19185_),
    .B2(_19186_),
    .ZN(_20267_));
 AND2_X4 _47450_ (.A1(_20266_),
    .A2(_20267_),
    .ZN(_20268_));
 OAI21_X1 _47451_ (.A(_20265_),
    .B1(_20268_),
    .B2(_20244_),
    .ZN(_04944_));
 NAND2_X1 _47452_ (.A1(_20231_),
    .A2(\icache.lce.lce_cmd_inst.data_r [15]),
    .ZN(_20269_));
 OAI21_X2 _47453_ (.A(_15645_),
    .B1(_19190_),
    .B2(_19191_),
    .ZN(_20270_));
 NAND3_X2 _47454_ (.A1(_19193_),
    .A2(_19194_),
    .A3(_16200_),
    .ZN(_20271_));
 NAND2_X4 _47455_ (.A1(_20270_),
    .A2(_20271_),
    .ZN(_20272_));
 OAI21_X1 _47456_ (.A(_20269_),
    .B1(_20272_),
    .B2(_20244_),
    .ZN(_04955_));
 NAND2_X1 _47457_ (.A1(_15351_),
    .A2(\icache.lce.lce_cmd_inst.data_r [16]),
    .ZN(_20273_));
 NAND3_X1 _47458_ (.A1(_19199_),
    .A2(_16360_),
    .A3(_19200_),
    .ZN(_20274_));
 OAI21_X1 _47459_ (.A(_15315_),
    .B1(_19202_),
    .B2(_19203_),
    .ZN(_20275_));
 AND2_X4 _47460_ (.A1(_20274_),
    .A2(_20275_),
    .ZN(_20276_));
 OAI21_X1 _47461_ (.A(_20273_),
    .B1(_20276_),
    .B2(_20244_),
    .ZN(_04966_));
 NAND2_X1 _47462_ (.A1(_15351_),
    .A2(\icache.lce.lce_cmd_inst.data_r [3]),
    .ZN(_20277_));
 OR3_X1 _47463_ (.A1(_19089_),
    .A2(_19090_),
    .A3(_15408_),
    .ZN(_20278_));
 OAI21_X1 _47464_ (.A(_15849_),
    .B1(_19085_),
    .B2(_19086_),
    .ZN(_20279_));
 AND2_X4 _47465_ (.A1(_20278_),
    .A2(_20279_),
    .ZN(_20280_));
 OAI21_X1 _47466_ (.A(_20277_),
    .B1(_20280_),
    .B2(_20244_),
    .ZN(_05222_));
 NAND2_X1 _47467_ (.A1(_15351_),
    .A2(\icache.lce.lce_cmd_inst.data_r [1]),
    .ZN(_20281_));
 NAND2_X1 _47468_ (.A1(_19069_),
    .A2(_17634_),
    .ZN(_20282_));
 OAI21_X2 _47469_ (.A(_15656_),
    .B1(_19071_),
    .B2(_19072_),
    .ZN(_20283_));
 NAND2_X4 _47470_ (.A1(_20282_),
    .A2(_20283_),
    .ZN(_20284_));
 OAI21_X1 _47471_ (.A(_20281_),
    .B1(_20284_),
    .B2(_15303_),
    .ZN(_05000_));
 NAND2_X1 _47472_ (.A1(_15351_),
    .A2(\icache.lce.lce_cmd_inst.data_r [2]),
    .ZN(_20285_));
 NOR3_X2 _47473_ (.A1(_19076_),
    .A2(_19077_),
    .A3(_16360_),
    .ZN(_20286_));
 AOI21_X2 _47474_ (.A(_17990_),
    .B1(_19079_),
    .B2(_19080_),
    .ZN(_20287_));
 NOR2_X4 _47475_ (.A1(_20286_),
    .A2(_20287_),
    .ZN(_20288_));
 OAI21_X1 _47476_ (.A(_20285_),
    .B1(_20288_),
    .B2(_15303_),
    .ZN(_05111_));
 MUX2_X2 _47477_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [0]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [53]),
    .S(_07973_),
    .Z(_20289_));
 AND2_X4 _47478_ (.A1(_20289_),
    .A2(lce_data_cmd_v_o),
    .ZN(lce_data_cmd_o[0]));
 MUX2_X1 _47479_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [1]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [54]),
    .S(_07973_),
    .Z(_20290_));
 AND2_X4 _47480_ (.A1(_20290_),
    .A2(lce_data_cmd_v_o),
    .ZN(lce_data_cmd_o[1]));
 MUX2_X1 _47481_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [2]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [55]),
    .S(_07973_),
    .Z(_20291_));
 AND2_X4 _47482_ (.A1(_20291_),
    .A2(lce_data_cmd_v_o),
    .ZN(lce_data_cmd_o[2]));
 MUX2_X2 _47483_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [3]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [56]),
    .S(_07973_),
    .Z(_20292_));
 AND2_X4 _47484_ (.A1(_20292_),
    .A2(lce_data_cmd_v_o),
    .ZN(lce_data_cmd_o[5]));
 OAI21_X1 _47485_ (.A(lce_data_cmd_v_o),
    .B1(_15297_),
    .B2(\icache.lce.lce_cmd_inst.data_r [0]),
    .ZN(_20293_));
 BUF_X32 _47486_ (.A(_15295_),
    .Z(_20294_));
 BUF_X32 _47487_ (.A(_20294_),
    .Z(_20295_));
 AOI21_X4 _47488_ (.A(_20293_),
    .B1(_15350_),
    .B2(_20295_),
    .ZN(lce_data_cmd_o[6]));
 OAI21_X2 _47489_ (.A(lce_data_cmd_v_o),
    .B1(_15297_),
    .B2(\icache.lce.lce_cmd_inst.data_r [1]),
    .ZN(_20296_));
 AOI21_X4 _47490_ (.A(_20296_),
    .B1(_20284_),
    .B2(_20295_),
    .ZN(lce_data_cmd_o[7]));
 OAI21_X1 _47491_ (.A(lce_data_cmd_v_o),
    .B1(_15297_),
    .B2(\icache.lce.lce_cmd_inst.data_r [2]),
    .ZN(_20297_));
 AOI21_X4 _47492_ (.A(_20297_),
    .B1(_20288_),
    .B2(_20295_),
    .ZN(lce_data_cmd_o[8]));
 OAI21_X2 _47493_ (.A(lce_data_cmd_v_o),
    .B1(_15297_),
    .B2(\icache.lce.lce_cmd_inst.data_r [3]),
    .ZN(_20298_));
 AOI21_X4 _47494_ (.A(_20298_),
    .B1(_20280_),
    .B2(_20295_),
    .ZN(lce_data_cmd_o[9]));
 OAI21_X2 _47495_ (.A(lce_data_cmd_v_o),
    .B1(_15297_),
    .B2(\icache.lce.lce_cmd_inst.data_r [4]),
    .ZN(_20299_));
 AOI21_X4 _47496_ (.A(_20299_),
    .B1(_20226_),
    .B2(_20295_),
    .ZN(lce_data_cmd_o[10]));
 BUF_X16 _47497_ (.A(_07607_),
    .Z(_20300_));
 BUF_X8 _47498_ (.A(_20300_),
    .Z(_20301_));
 OAI21_X2 _47499_ (.A(_20301_),
    .B1(_15297_),
    .B2(\icache.lce.lce_cmd_inst.data_r [5]),
    .ZN(_20302_));
 AOI21_X4 _47500_ (.A(_20302_),
    .B1(_20230_),
    .B2(_20295_),
    .ZN(lce_data_cmd_o[11]));
 OAI21_X2 _47501_ (.A(_20301_),
    .B1(_15297_),
    .B2(\icache.lce.lce_cmd_inst.data_r [6]),
    .ZN(_20303_));
 AOI21_X4 _47502_ (.A(_20303_),
    .B1(_20235_),
    .B2(_20295_),
    .ZN(lce_data_cmd_o[12]));
 BUF_X8 _47503_ (.A(_15296_),
    .Z(_20304_));
 OAI21_X2 _47504_ (.A(_20301_),
    .B1(_20304_),
    .B2(\icache.lce.lce_cmd_inst.data_r [7]),
    .ZN(_20305_));
 AOI21_X4 _47505_ (.A(_20305_),
    .B1(_20239_),
    .B2(_20295_),
    .ZN(lce_data_cmd_o[13]));
 OAI21_X2 _47506_ (.A(_20301_),
    .B1(_20304_),
    .B2(\icache.lce.lce_cmd_inst.data_r [8]),
    .ZN(_20306_));
 AOI21_X4 _47507_ (.A(_20306_),
    .B1(_20243_),
    .B2(_20295_),
    .ZN(lce_data_cmd_o[14]));
 OAI21_X2 _47508_ (.A(_20301_),
    .B1(_20304_),
    .B2(\icache.lce.lce_cmd_inst.data_r [9]),
    .ZN(_20307_));
 AOI21_X4 _47509_ (.A(_20307_),
    .B1(_20248_),
    .B2(_20295_),
    .ZN(lce_data_cmd_o[15]));
 OAI21_X2 _47510_ (.A(_20301_),
    .B1(_20304_),
    .B2(\icache.lce.lce_cmd_inst.data_r [10]),
    .ZN(_20308_));
 BUF_X16 _47511_ (.A(_20294_),
    .Z(_20309_));
 AOI21_X4 _47512_ (.A(_20308_),
    .B1(_20252_),
    .B2(_20309_),
    .ZN(lce_data_cmd_o[16]));
 OAI21_X2 _47513_ (.A(_20301_),
    .B1(_20304_),
    .B2(\icache.lce.lce_cmd_inst.data_r [11]),
    .ZN(_20310_));
 AOI21_X4 _47514_ (.A(_20310_),
    .B1(_20256_),
    .B2(_20309_),
    .ZN(lce_data_cmd_o[17]));
 OAI21_X1 _47515_ (.A(_20301_),
    .B1(_20304_),
    .B2(\icache.lce.lce_cmd_inst.data_r [12]),
    .ZN(_20311_));
 AOI21_X4 _47516_ (.A(_20311_),
    .B1(_20260_),
    .B2(_20309_),
    .ZN(lce_data_cmd_o[18]));
 OAI21_X1 _47517_ (.A(_20301_),
    .B1(_20304_),
    .B2(\icache.lce.lce_cmd_inst.data_r [13]),
    .ZN(_20312_));
 AOI21_X4 _47518_ (.A(_20312_),
    .B1(_20264_),
    .B2(_20309_),
    .ZN(lce_data_cmd_o[19]));
 OAI21_X1 _47519_ (.A(_20301_),
    .B1(_20304_),
    .B2(\icache.lce.lce_cmd_inst.data_r [14]),
    .ZN(_20313_));
 AOI21_X4 _47520_ (.A(_20313_),
    .B1(_20268_),
    .B2(_20309_),
    .ZN(lce_data_cmd_o[20]));
 BUF_X8 _47521_ (.A(_20300_),
    .Z(_20314_));
 OAI21_X2 _47522_ (.A(_20314_),
    .B1(_20304_),
    .B2(\icache.lce.lce_cmd_inst.data_r [15]),
    .ZN(_20315_));
 AOI21_X4 _47523_ (.A(_20315_),
    .B1(_20272_),
    .B2(_20309_),
    .ZN(lce_data_cmd_o[21]));
 OAI21_X2 _47524_ (.A(_20314_),
    .B1(_20304_),
    .B2(\icache.lce.lce_cmd_inst.data_r [16]),
    .ZN(_20316_));
 AOI21_X4 _47525_ (.A(_20316_),
    .B1(_20276_),
    .B2(_20309_),
    .ZN(lce_data_cmd_o[22]));
 BUF_X8 _47526_ (.A(_15296_),
    .Z(_20317_));
 OAI21_X2 _47527_ (.A(_20314_),
    .B1(_20317_),
    .B2(\icache.lce.lce_cmd_inst.data_r [17]),
    .ZN(_20318_));
 AOI21_X4 _47528_ (.A(_20318_),
    .B1(_19899_),
    .B2(_20309_),
    .ZN(lce_data_cmd_o[23]));
 OAI21_X2 _47529_ (.A(_20314_),
    .B1(_20317_),
    .B2(\icache.lce.lce_cmd_inst.data_r [18]),
    .ZN(_20319_));
 AOI21_X4 _47530_ (.A(_20319_),
    .B1(_19903_),
    .B2(_20309_),
    .ZN(lce_data_cmd_o[24]));
 OAI21_X2 _47531_ (.A(_20314_),
    .B1(_20317_),
    .B2(\icache.lce.lce_cmd_inst.data_r [19]),
    .ZN(_20320_));
 AOI21_X4 _47532_ (.A(_20320_),
    .B1(_19909_),
    .B2(_20309_),
    .ZN(lce_data_cmd_o[25]));
 OAI21_X2 _47533_ (.A(_20314_),
    .B1(_20317_),
    .B2(\icache.lce.lce_cmd_inst.data_r [20]),
    .ZN(_20321_));
 BUF_X16 _47534_ (.A(_20294_),
    .Z(_20322_));
 AOI21_X4 _47535_ (.A(_20321_),
    .B1(_19913_),
    .B2(_20322_),
    .ZN(lce_data_cmd_o[26]));
 OAI21_X2 _47536_ (.A(_20314_),
    .B1(_20317_),
    .B2(\icache.lce.lce_cmd_inst.data_r [21]),
    .ZN(_20323_));
 AOI21_X4 _47537_ (.A(_20323_),
    .B1(_19917_),
    .B2(_20322_),
    .ZN(lce_data_cmd_o[27]));
 OAI21_X2 _47538_ (.A(_20314_),
    .B1(_20317_),
    .B2(\icache.lce.lce_cmd_inst.data_r [22]),
    .ZN(_20324_));
 AOI21_X4 _47539_ (.A(_20324_),
    .B1(_19921_),
    .B2(_20322_),
    .ZN(lce_data_cmd_o[28]));
 OAI21_X2 _47540_ (.A(_20314_),
    .B1(_20317_),
    .B2(\icache.lce.lce_cmd_inst.data_r [23]),
    .ZN(_20325_));
 AOI21_X4 _47541_ (.A(_20325_),
    .B1(_19925_),
    .B2(_20322_),
    .ZN(lce_data_cmd_o[29]));
 OAI21_X2 _47542_ (.A(_20314_),
    .B1(_20317_),
    .B2(\icache.lce.lce_cmd_inst.data_r [24]),
    .ZN(_20326_));
 AOI21_X4 _47543_ (.A(_20326_),
    .B1(_19929_),
    .B2(_20322_),
    .ZN(lce_data_cmd_o[30]));
 BUF_X8 _47544_ (.A(_20300_),
    .Z(_20327_));
 OAI21_X2 _47545_ (.A(_20327_),
    .B1(_20317_),
    .B2(\icache.lce.lce_cmd_inst.data_r [25]),
    .ZN(_20328_));
 AOI21_X4 _47546_ (.A(_20328_),
    .B1(_19933_),
    .B2(_20322_),
    .ZN(lce_data_cmd_o[31]));
 OAI21_X2 _47547_ (.A(_20327_),
    .B1(_20317_),
    .B2(\icache.lce.lce_cmd_inst.data_r [26]),
    .ZN(_20329_));
 AOI21_X4 _47548_ (.A(_20329_),
    .B1(_19938_),
    .B2(_20322_),
    .ZN(lce_data_cmd_o[32]));
 BUF_X8 _47549_ (.A(_15296_),
    .Z(_20330_));
 OAI21_X2 _47550_ (.A(_20327_),
    .B1(_20330_),
    .B2(\icache.lce.lce_cmd_inst.data_r [27]),
    .ZN(_20331_));
 AOI21_X4 _47551_ (.A(_20331_),
    .B1(_19943_),
    .B2(_20322_),
    .ZN(lce_data_cmd_o[33]));
 OAI21_X2 _47552_ (.A(_20327_),
    .B1(_20330_),
    .B2(\icache.lce.lce_cmd_inst.data_r [28]),
    .ZN(_20332_));
 AOI21_X4 _47553_ (.A(_20332_),
    .B1(_19947_),
    .B2(_20322_),
    .ZN(lce_data_cmd_o[34]));
 OAI21_X2 _47554_ (.A(_20327_),
    .B1(_20330_),
    .B2(\icache.lce.lce_cmd_inst.data_r [29]),
    .ZN(_20333_));
 AOI21_X4 _47555_ (.A(_20333_),
    .B1(_19953_),
    .B2(_20322_),
    .ZN(lce_data_cmd_o[35]));
 OAI21_X2 _47556_ (.A(_20327_),
    .B1(_20330_),
    .B2(\icache.lce.lce_cmd_inst.data_r [30]),
    .ZN(_20334_));
 BUF_X8 _47557_ (.A(_20294_),
    .Z(_20335_));
 AOI21_X4 _47558_ (.A(_20334_),
    .B1(_19957_),
    .B2(_20335_),
    .ZN(lce_data_cmd_o[36]));
 OAI21_X2 _47559_ (.A(_20327_),
    .B1(_20330_),
    .B2(\icache.lce.lce_cmd_inst.data_r [31]),
    .ZN(_20336_));
 AOI21_X4 _47560_ (.A(_20336_),
    .B1(_19961_),
    .B2(_20335_),
    .ZN(lce_data_cmd_o[37]));
 OAI21_X2 _47561_ (.A(_20327_),
    .B1(_20330_),
    .B2(\icache.lce.lce_cmd_inst.data_r [32]),
    .ZN(_20337_));
 AOI21_X4 _47562_ (.A(_20337_),
    .B1(_19966_),
    .B2(_20335_),
    .ZN(lce_data_cmd_o[38]));
 OAI21_X2 _47563_ (.A(_20327_),
    .B1(_20330_),
    .B2(\icache.lce.lce_cmd_inst.data_r [33]),
    .ZN(_20338_));
 AOI21_X4 _47564_ (.A(_20338_),
    .B1(_19970_),
    .B2(_20335_),
    .ZN(lce_data_cmd_o[39]));
 OAI21_X2 _47565_ (.A(_20327_),
    .B1(_20330_),
    .B2(\icache.lce.lce_cmd_inst.data_r [34]),
    .ZN(_20339_));
 AOI21_X4 _47566_ (.A(_20339_),
    .B1(_19974_),
    .B2(_20335_),
    .ZN(lce_data_cmd_o[40]));
 BUF_X32 _47567_ (.A(_07608_),
    .Z(_20340_));
 BUF_X4 _47568_ (.A(_20340_),
    .Z(_20341_));
 OAI21_X2 _47569_ (.A(_20341_),
    .B1(_20330_),
    .B2(\icache.lce.lce_cmd_inst.data_r [35]),
    .ZN(_20342_));
 AOI21_X4 _47570_ (.A(_20342_),
    .B1(_19978_),
    .B2(_20335_),
    .ZN(lce_data_cmd_o[41]));
 OAI21_X2 _47571_ (.A(_20341_),
    .B1(_20330_),
    .B2(\icache.lce.lce_cmd_inst.data_r [36]),
    .ZN(_20343_));
 AOI21_X4 _47572_ (.A(_20343_),
    .B1(_19983_),
    .B2(_20335_),
    .ZN(lce_data_cmd_o[42]));
 BUF_X32 _47573_ (.A(_15295_),
    .Z(_20344_));
 BUF_X4 _47574_ (.A(_20344_),
    .Z(_20345_));
 OAI21_X2 _47575_ (.A(_20341_),
    .B1(_20345_),
    .B2(\icache.lce.lce_cmd_inst.data_r [37]),
    .ZN(_20346_));
 AOI21_X4 _47576_ (.A(_20346_),
    .B1(_19987_),
    .B2(_20335_),
    .ZN(lce_data_cmd_o[43]));
 OAI21_X2 _47577_ (.A(_20341_),
    .B1(_20345_),
    .B2(\icache.lce.lce_cmd_inst.data_r [38]),
    .ZN(_20347_));
 AOI21_X4 _47578_ (.A(_20347_),
    .B1(_19991_),
    .B2(_20335_),
    .ZN(lce_data_cmd_o[44]));
 OAI21_X2 _47579_ (.A(_20341_),
    .B1(_20345_),
    .B2(\icache.lce.lce_cmd_inst.data_r [39]),
    .ZN(_20348_));
 AOI21_X4 _47580_ (.A(_20348_),
    .B1(_19996_),
    .B2(_20335_),
    .ZN(lce_data_cmd_o[45]));
 OAI21_X2 _47581_ (.A(_20341_),
    .B1(_20345_),
    .B2(\icache.lce.lce_cmd_inst.data_r [40]),
    .ZN(_20349_));
 BUF_X8 _47582_ (.A(_20294_),
    .Z(_20350_));
 AOI21_X4 _47583_ (.A(_20349_),
    .B1(_20000_),
    .B2(_20350_),
    .ZN(lce_data_cmd_o[46]));
 OAI21_X2 _47584_ (.A(_20341_),
    .B1(_20345_),
    .B2(\icache.lce.lce_cmd_inst.data_r [41]),
    .ZN(_20351_));
 AOI21_X4 _47585_ (.A(_20351_),
    .B1(_20004_),
    .B2(_20350_),
    .ZN(lce_data_cmd_o[47]));
 OAI21_X2 _47586_ (.A(_20341_),
    .B1(_20345_),
    .B2(\icache.lce.lce_cmd_inst.data_r [42]),
    .ZN(_20352_));
 AOI21_X4 _47587_ (.A(_20352_),
    .B1(_20008_),
    .B2(_20350_),
    .ZN(lce_data_cmd_o[48]));
 OAI21_X2 _47588_ (.A(_20341_),
    .B1(_20345_),
    .B2(\icache.lce.lce_cmd_inst.data_r [43]),
    .ZN(_20353_));
 AOI21_X4 _47589_ (.A(_20353_),
    .B1(_20012_),
    .B2(_20350_),
    .ZN(lce_data_cmd_o[49]));
 OAI21_X2 _47590_ (.A(_20341_),
    .B1(_20345_),
    .B2(\icache.lce.lce_cmd_inst.data_r [44]),
    .ZN(_20354_));
 AOI21_X4 _47591_ (.A(_20354_),
    .B1(_20016_),
    .B2(_20350_),
    .ZN(lce_data_cmd_o[50]));
 BUF_X8 _47592_ (.A(_20340_),
    .Z(_20355_));
 OAI21_X2 _47593_ (.A(_20355_),
    .B1(_20345_),
    .B2(\icache.lce.lce_cmd_inst.data_r [45]),
    .ZN(_20356_));
 AOI21_X4 _47594_ (.A(_20356_),
    .B1(_20020_),
    .B2(_20350_),
    .ZN(lce_data_cmd_o[51]));
 OAI21_X2 _47595_ (.A(_20355_),
    .B1(_20345_),
    .B2(\icache.lce.lce_cmd_inst.data_r [46]),
    .ZN(_20357_));
 AOI21_X4 _47596_ (.A(_20357_),
    .B1(_20025_),
    .B2(_20350_),
    .ZN(lce_data_cmd_o[52]));
 BUF_X8 _47597_ (.A(_20344_),
    .Z(_20358_));
 OAI21_X2 _47598_ (.A(_20355_),
    .B1(_20358_),
    .B2(\icache.lce.lce_cmd_inst.data_r [47]),
    .ZN(_20359_));
 AOI21_X4 _47599_ (.A(_20359_),
    .B1(_20029_),
    .B2(_20350_),
    .ZN(lce_data_cmd_o[53]));
 OAI21_X2 _47600_ (.A(_20355_),
    .B1(_20358_),
    .B2(\icache.lce.lce_cmd_inst.data_r [48]),
    .ZN(_20360_));
 AOI21_X4 _47601_ (.A(_20360_),
    .B1(_20033_),
    .B2(_20350_),
    .ZN(lce_data_cmd_o[54]));
 OAI21_X2 _47602_ (.A(_20355_),
    .B1(_20358_),
    .B2(\icache.lce.lce_cmd_inst.data_r [49]),
    .ZN(_20361_));
 AOI21_X4 _47603_ (.A(_20361_),
    .B1(_20038_),
    .B2(_20350_),
    .ZN(lce_data_cmd_o[55]));
 OAI21_X2 _47604_ (.A(_20355_),
    .B1(_20358_),
    .B2(\icache.lce.lce_cmd_inst.data_r [50]),
    .ZN(_20362_));
 BUF_X32 _47605_ (.A(_15295_),
    .Z(_20363_));
 BUF_X32 _47606_ (.A(_20363_),
    .Z(_20364_));
 BUF_X8 _47607_ (.A(_20364_),
    .Z(_20365_));
 AOI21_X4 _47608_ (.A(_20362_),
    .B1(_20042_),
    .B2(_20365_),
    .ZN(lce_data_cmd_o[56]));
 OAI21_X2 _47609_ (.A(_20355_),
    .B1(_20358_),
    .B2(\icache.lce.lce_cmd_inst.data_r [51]),
    .ZN(_20366_));
 AOI21_X4 _47610_ (.A(_20366_),
    .B1(_20046_),
    .B2(_20365_),
    .ZN(lce_data_cmd_o[57]));
 OAI21_X2 _47611_ (.A(_20355_),
    .B1(_20358_),
    .B2(\icache.lce.lce_cmd_inst.data_r [52]),
    .ZN(_20367_));
 AOI21_X4 _47612_ (.A(_20367_),
    .B1(_20050_),
    .B2(_20365_),
    .ZN(lce_data_cmd_o[58]));
 OAI21_X2 _47613_ (.A(_20355_),
    .B1(_20358_),
    .B2(\icache.lce.lce_cmd_inst.data_r [53]),
    .ZN(_20368_));
 AOI21_X4 _47614_ (.A(_20368_),
    .B1(_20054_),
    .B2(_20365_),
    .ZN(lce_data_cmd_o[59]));
 OAI21_X2 _47615_ (.A(_20355_),
    .B1(_20358_),
    .B2(\icache.lce.lce_cmd_inst.data_r [54]),
    .ZN(_20369_));
 AOI21_X4 _47616_ (.A(_20369_),
    .B1(_20058_),
    .B2(_20365_),
    .ZN(lce_data_cmd_o[60]));
 BUF_X16 _47617_ (.A(_20340_),
    .Z(_20370_));
 OAI21_X2 _47618_ (.A(_20370_),
    .B1(_20358_),
    .B2(\icache.lce.lce_cmd_inst.data_r [55]),
    .ZN(_20371_));
 AOI21_X4 _47619_ (.A(_20371_),
    .B1(_20062_),
    .B2(_20365_),
    .ZN(lce_data_cmd_o[61]));
 OAI21_X2 _47620_ (.A(_20370_),
    .B1(_20358_),
    .B2(\icache.lce.lce_cmd_inst.data_r [56]),
    .ZN(_20372_));
 AOI21_X4 _47621_ (.A(_20372_),
    .B1(_20067_),
    .B2(_20365_),
    .ZN(lce_data_cmd_o[62]));
 BUF_X16 _47622_ (.A(_20344_),
    .Z(_20373_));
 OAI21_X2 _47623_ (.A(_20370_),
    .B1(_20373_),
    .B2(\icache.lce.lce_cmd_inst.data_r [57]),
    .ZN(_20374_));
 AOI21_X4 _47624_ (.A(_20374_),
    .B1(_20071_),
    .B2(_20365_),
    .ZN(lce_data_cmd_o[63]));
 OAI21_X2 _47625_ (.A(_20370_),
    .B1(_20373_),
    .B2(\icache.lce.lce_cmd_inst.data_r [58]),
    .ZN(_20375_));
 AOI21_X4 _47626_ (.A(_20375_),
    .B1(_20075_),
    .B2(_20365_),
    .ZN(lce_data_cmd_o[64]));
 OAI21_X2 _47627_ (.A(_20370_),
    .B1(_20373_),
    .B2(\icache.lce.lce_cmd_inst.data_r [59]),
    .ZN(_20376_));
 AOI21_X4 _47628_ (.A(_20376_),
    .B1(_20080_),
    .B2(_20365_),
    .ZN(lce_data_cmd_o[65]));
 OAI21_X2 _47629_ (.A(_20370_),
    .B1(_20373_),
    .B2(\icache.lce.lce_cmd_inst.data_r [60]),
    .ZN(_20377_));
 BUF_X16 _47630_ (.A(_20364_),
    .Z(_20378_));
 AOI21_X4 _47631_ (.A(_20377_),
    .B1(_20084_),
    .B2(_20378_),
    .ZN(lce_data_cmd_o[66]));
 OAI21_X2 _47632_ (.A(_20370_),
    .B1(_20373_),
    .B2(\icache.lce.lce_cmd_inst.data_r [61]),
    .ZN(_20379_));
 AOI21_X4 _47633_ (.A(_20379_),
    .B1(_20088_),
    .B2(_20378_),
    .ZN(lce_data_cmd_o[67]));
 OAI21_X2 _47634_ (.A(_20370_),
    .B1(_20373_),
    .B2(\icache.lce.lce_cmd_inst.data_r [62]),
    .ZN(_20380_));
 AOI21_X4 _47635_ (.A(_20380_),
    .B1(_20092_),
    .B2(_20378_),
    .ZN(lce_data_cmd_o[68]));
 OAI21_X2 _47636_ (.A(_20370_),
    .B1(_20373_),
    .B2(\icache.lce.lce_cmd_inst.data_r [63]),
    .ZN(_20381_));
 AOI21_X4 _47637_ (.A(_20381_),
    .B1(_20096_),
    .B2(_20378_),
    .ZN(lce_data_cmd_o[69]));
 OAI21_X2 _47638_ (.A(_20370_),
    .B1(_20373_),
    .B2(\icache.lce.lce_cmd_inst.data_r [64]),
    .ZN(_20382_));
 AOI21_X4 _47639_ (.A(_20382_),
    .B1(_20100_),
    .B2(_20378_),
    .ZN(lce_data_cmd_o[70]));
 BUF_X8 _47640_ (.A(_20340_),
    .Z(_20383_));
 OAI21_X2 _47641_ (.A(_20383_),
    .B1(_20373_),
    .B2(\icache.lce.lce_cmd_inst.data_r [65]),
    .ZN(_20384_));
 AOI21_X4 _47642_ (.A(_20384_),
    .B1(_20104_),
    .B2(_20378_),
    .ZN(lce_data_cmd_o[71]));
 OAI21_X1 _47643_ (.A(_20383_),
    .B1(_20373_),
    .B2(\icache.lce.lce_cmd_inst.data_r [66]),
    .ZN(_20385_));
 AOI21_X4 _47644_ (.A(_20385_),
    .B1(_20109_),
    .B2(_20378_),
    .ZN(lce_data_cmd_o[72]));
 BUF_X8 _47645_ (.A(_20344_),
    .Z(_20386_));
 OAI21_X2 _47646_ (.A(_20383_),
    .B1(_20386_),
    .B2(\icache.lce.lce_cmd_inst.data_r [67]),
    .ZN(_20387_));
 AOI21_X4 _47647_ (.A(_20387_),
    .B1(_20113_),
    .B2(_20378_),
    .ZN(lce_data_cmd_o[73]));
 OAI21_X2 _47648_ (.A(_20383_),
    .B1(_20386_),
    .B2(\icache.lce.lce_cmd_inst.data_r [68]),
    .ZN(_20388_));
 AOI21_X4 _47649_ (.A(_20388_),
    .B1(_20117_),
    .B2(_20378_),
    .ZN(lce_data_cmd_o[74]));
 OAI21_X2 _47650_ (.A(_20383_),
    .B1(_20386_),
    .B2(\icache.lce.lce_cmd_inst.data_r [69]),
    .ZN(_20389_));
 AOI21_X4 _47651_ (.A(_20389_),
    .B1(_20122_),
    .B2(_20378_),
    .ZN(lce_data_cmd_o[75]));
 OAI21_X2 _47652_ (.A(_20383_),
    .B1(_20386_),
    .B2(\icache.lce.lce_cmd_inst.data_r [70]),
    .ZN(_20390_));
 BUF_X16 _47653_ (.A(_20364_),
    .Z(_20391_));
 AOI21_X4 _47654_ (.A(_20390_),
    .B1(_20126_),
    .B2(_20391_),
    .ZN(lce_data_cmd_o[76]));
 OAI21_X1 _47655_ (.A(_20383_),
    .B1(_20386_),
    .B2(\icache.lce.lce_cmd_inst.data_r [71]),
    .ZN(_20392_));
 AOI21_X4 _47656_ (.A(_20392_),
    .B1(_20130_),
    .B2(_20391_),
    .ZN(lce_data_cmd_o[77]));
 OAI21_X1 _47657_ (.A(_20383_),
    .B1(_20386_),
    .B2(\icache.lce.lce_cmd_inst.data_r [72]),
    .ZN(_20393_));
 AOI21_X4 _47658_ (.A(_20393_),
    .B1(_20134_),
    .B2(_20391_),
    .ZN(lce_data_cmd_o[78]));
 OAI21_X2 _47659_ (.A(_20383_),
    .B1(_20386_),
    .B2(\icache.lce.lce_cmd_inst.data_r [73]),
    .ZN(_20394_));
 AOI21_X4 _47660_ (.A(_20394_),
    .B1(_20138_),
    .B2(_20391_),
    .ZN(lce_data_cmd_o[79]));
 OAI21_X2 _47661_ (.A(_20383_),
    .B1(_20386_),
    .B2(\icache.lce.lce_cmd_inst.data_r [74]),
    .ZN(_20395_));
 AOI21_X4 _47662_ (.A(_20395_),
    .B1(_20142_),
    .B2(_20391_),
    .ZN(lce_data_cmd_o[80]));
 BUF_X8 _47663_ (.A(_20340_),
    .Z(_20396_));
 OAI21_X2 _47664_ (.A(_20396_),
    .B1(_20386_),
    .B2(\icache.lce.lce_cmd_inst.data_r [75]),
    .ZN(_20397_));
 AOI21_X4 _47665_ (.A(_20397_),
    .B1(_20146_),
    .B2(_20391_),
    .ZN(lce_data_cmd_o[81]));
 OAI21_X2 _47666_ (.A(_20396_),
    .B1(_20386_),
    .B2(\icache.lce.lce_cmd_inst.data_r [76]),
    .ZN(_20398_));
 AOI21_X4 _47667_ (.A(_20398_),
    .B1(_20151_),
    .B2(_20391_),
    .ZN(lce_data_cmd_o[82]));
 BUF_X8 _47668_ (.A(_20344_),
    .Z(_20399_));
 OAI21_X2 _47669_ (.A(_20396_),
    .B1(_20399_),
    .B2(\icache.lce.lce_cmd_inst.data_r [77]),
    .ZN(_20400_));
 AOI21_X4 _47670_ (.A(_20400_),
    .B1(_20155_),
    .B2(_20391_),
    .ZN(lce_data_cmd_o[83]));
 OAI21_X1 _47671_ (.A(_20396_),
    .B1(_20399_),
    .B2(\icache.lce.lce_cmd_inst.data_r [78]),
    .ZN(_20401_));
 AOI21_X4 _47672_ (.A(_20401_),
    .B1(_20159_),
    .B2(_20391_),
    .ZN(lce_data_cmd_o[84]));
 OAI21_X2 _47673_ (.A(_20396_),
    .B1(_20399_),
    .B2(\icache.lce.lce_cmd_inst.data_r [79]),
    .ZN(_20402_));
 AOI21_X4 _47674_ (.A(_20402_),
    .B1(_20164_),
    .B2(_20391_),
    .ZN(lce_data_cmd_o[85]));
 OAI21_X2 _47675_ (.A(_20396_),
    .B1(_20399_),
    .B2(\icache.lce.lce_cmd_inst.data_r [80]),
    .ZN(_20403_));
 BUF_X16 _47676_ (.A(_20364_),
    .Z(_20404_));
 AOI21_X4 _47677_ (.A(_20403_),
    .B1(_20168_),
    .B2(_20404_),
    .ZN(lce_data_cmd_o[86]));
 OAI21_X2 _47678_ (.A(_20396_),
    .B1(_20399_),
    .B2(\icache.lce.lce_cmd_inst.data_r [81]),
    .ZN(_20405_));
 AOI21_X4 _47679_ (.A(_20405_),
    .B1(_20172_),
    .B2(_20404_),
    .ZN(lce_data_cmd_o[87]));
 OAI21_X1 _47680_ (.A(_20396_),
    .B1(_20399_),
    .B2(\icache.lce.lce_cmd_inst.data_r [82]),
    .ZN(_20406_));
 AOI21_X4 _47681_ (.A(_20406_),
    .B1(_20176_),
    .B2(_20404_),
    .ZN(lce_data_cmd_o[88]));
 OAI21_X2 _47682_ (.A(_20396_),
    .B1(_20399_),
    .B2(\icache.lce.lce_cmd_inst.data_r [83]),
    .ZN(_20407_));
 AOI21_X4 _47683_ (.A(_20407_),
    .B1(_20180_),
    .B2(_20404_),
    .ZN(lce_data_cmd_o[89]));
 OAI21_X2 _47684_ (.A(_20396_),
    .B1(_20399_),
    .B2(\icache.lce.lce_cmd_inst.data_r [84]),
    .ZN(_20408_));
 AOI21_X4 _47685_ (.A(_20408_),
    .B1(_20184_),
    .B2(_20404_),
    .ZN(lce_data_cmd_o[90]));
 BUF_X8 _47686_ (.A(_20340_),
    .Z(_20409_));
 OAI21_X2 _47687_ (.A(_20409_),
    .B1(_20399_),
    .B2(\icache.lce.lce_cmd_inst.data_r [85]),
    .ZN(_20410_));
 AOI21_X4 _47688_ (.A(_20410_),
    .B1(_20188_),
    .B2(_20404_),
    .ZN(lce_data_cmd_o[91]));
 OAI21_X2 _47689_ (.A(_20409_),
    .B1(_20399_),
    .B2(\icache.lce.lce_cmd_inst.data_r [86]),
    .ZN(_20411_));
 AOI21_X4 _47690_ (.A(_20411_),
    .B1(_20193_),
    .B2(_20404_),
    .ZN(lce_data_cmd_o[92]));
 BUF_X8 _47691_ (.A(_20344_),
    .Z(_20412_));
 OAI21_X2 _47692_ (.A(_20409_),
    .B1(_20412_),
    .B2(\icache.lce.lce_cmd_inst.data_r [87]),
    .ZN(_20413_));
 AOI21_X4 _47693_ (.A(_20413_),
    .B1(_20197_),
    .B2(_20404_),
    .ZN(lce_data_cmd_o[93]));
 OAI21_X2 _47694_ (.A(_20409_),
    .B1(_20412_),
    .B2(\icache.lce.lce_cmd_inst.data_r [88]),
    .ZN(_20414_));
 AOI21_X4 _47695_ (.A(_20414_),
    .B1(_20201_),
    .B2(_20404_),
    .ZN(lce_data_cmd_o[94]));
 OAI21_X1 _47696_ (.A(_20409_),
    .B1(_20412_),
    .B2(\icache.lce.lce_cmd_inst.data_r [89]),
    .ZN(_20415_));
 AOI21_X4 _47697_ (.A(_20415_),
    .B1(_20206_),
    .B2(_20404_),
    .ZN(lce_data_cmd_o[95]));
 OAI21_X2 _47698_ (.A(_20409_),
    .B1(_20412_),
    .B2(\icache.lce.lce_cmd_inst.data_r [90]),
    .ZN(_20416_));
 BUF_X16 _47699_ (.A(_20364_),
    .Z(_20417_));
 AOI21_X4 _47700_ (.A(_20416_),
    .B1(_20210_),
    .B2(_20417_),
    .ZN(lce_data_cmd_o[96]));
 OAI21_X2 _47701_ (.A(_20409_),
    .B1(_20412_),
    .B2(\icache.lce.lce_cmd_inst.data_r [91]),
    .ZN(_20418_));
 AOI21_X4 _47702_ (.A(_20418_),
    .B1(_20214_),
    .B2(_20417_),
    .ZN(lce_data_cmd_o[97]));
 OAI21_X2 _47703_ (.A(_20409_),
    .B1(_20412_),
    .B2(\icache.lce.lce_cmd_inst.data_r [92]),
    .ZN(_20419_));
 AOI21_X4 _47704_ (.A(_20419_),
    .B1(_20218_),
    .B2(_20417_),
    .ZN(lce_data_cmd_o[98]));
 OAI21_X2 _47705_ (.A(_20409_),
    .B1(_20412_),
    .B2(\icache.lce.lce_cmd_inst.data_r [93]),
    .ZN(_20420_));
 AOI21_X4 _47706_ (.A(_20420_),
    .B1(_20222_),
    .B2(_20417_),
    .ZN(lce_data_cmd_o[99]));
 OAI21_X2 _47707_ (.A(_20409_),
    .B1(_20412_),
    .B2(\icache.lce.lce_cmd_inst.data_r [94]),
    .ZN(_20421_));
 AOI21_X4 _47708_ (.A(_20421_),
    .B1(_19886_),
    .B2(_20417_),
    .ZN(lce_data_cmd_o[100]));
 BUF_X4 _47709_ (.A(_20340_),
    .Z(_20422_));
 OAI21_X2 _47710_ (.A(_20422_),
    .B1(_20412_),
    .B2(\icache.lce.lce_cmd_inst.data_r [95]),
    .ZN(_20423_));
 AOI21_X4 _47711_ (.A(_20423_),
    .B1(_19890_),
    .B2(_20417_),
    .ZN(lce_data_cmd_o[101]));
 OAI21_X2 _47712_ (.A(_20422_),
    .B1(_20412_),
    .B2(\icache.lce.lce_cmd_inst.data_r [96]),
    .ZN(_20424_));
 AOI21_X4 _47713_ (.A(_20424_),
    .B1(_19895_),
    .B2(_20417_),
    .ZN(lce_data_cmd_o[102]));
 BUF_X8 _47714_ (.A(_20344_),
    .Z(_20425_));
 OAI21_X2 _47715_ (.A(_20422_),
    .B1(_20425_),
    .B2(\icache.lce.lce_cmd_inst.data_r [97]),
    .ZN(_20426_));
 AOI21_X4 _47716_ (.A(_20426_),
    .B1(_19806_),
    .B2(_20417_),
    .ZN(lce_data_cmd_o[103]));
 OAI21_X2 _47717_ (.A(_20422_),
    .B1(_20425_),
    .B2(\icache.lce.lce_cmd_inst.data_r [98]),
    .ZN(_20427_));
 AOI21_X4 _47718_ (.A(_20427_),
    .B1(_19811_),
    .B2(_20417_),
    .ZN(lce_data_cmd_o[104]));
 OAI21_X2 _47719_ (.A(_20422_),
    .B1(_20425_),
    .B2(\icache.lce.lce_cmd_inst.data_r [99]),
    .ZN(_20428_));
 AOI21_X4 _47720_ (.A(_20428_),
    .B1(_19815_),
    .B2(_20417_),
    .ZN(lce_data_cmd_o[105]));
 OAI21_X2 _47721_ (.A(_20422_),
    .B1(_20425_),
    .B2(\icache.lce.lce_cmd_inst.data_r [100]),
    .ZN(_20429_));
 BUF_X16 _47722_ (.A(_20364_),
    .Z(_20430_));
 AOI21_X4 _47723_ (.A(_20429_),
    .B1(_19819_),
    .B2(_20430_),
    .ZN(lce_data_cmd_o[106]));
 OAI21_X2 _47724_ (.A(_20422_),
    .B1(_20425_),
    .B2(\icache.lce.lce_cmd_inst.data_r [101]),
    .ZN(_20431_));
 AOI21_X4 _47725_ (.A(_20431_),
    .B1(_19824_),
    .B2(_20430_),
    .ZN(lce_data_cmd_o[107]));
 OAI21_X2 _47726_ (.A(_20422_),
    .B1(_20425_),
    .B2(\icache.lce.lce_cmd_inst.data_r [102]),
    .ZN(_20432_));
 AOI21_X4 _47727_ (.A(_20432_),
    .B1(_19828_),
    .B2(_20430_),
    .ZN(lce_data_cmd_o[108]));
 OAI21_X2 _47728_ (.A(_20422_),
    .B1(_20425_),
    .B2(\icache.lce.lce_cmd_inst.data_r [103]),
    .ZN(_20433_));
 AOI21_X4 _47729_ (.A(_20433_),
    .B1(_19832_),
    .B2(_20430_),
    .ZN(lce_data_cmd_o[109]));
 OAI21_X1 _47730_ (.A(_20422_),
    .B1(_20425_),
    .B2(\icache.lce.lce_cmd_inst.data_r [104]),
    .ZN(_20434_));
 AOI21_X4 _47731_ (.A(_20434_),
    .B1(_19836_),
    .B2(_20430_),
    .ZN(lce_data_cmd_o[110]));
 BUF_X4 _47732_ (.A(_20340_),
    .Z(_20435_));
 OAI21_X2 _47733_ (.A(_20435_),
    .B1(_20425_),
    .B2(\icache.lce.lce_cmd_inst.data_r [105]),
    .ZN(_20436_));
 AOI21_X4 _47734_ (.A(_20436_),
    .B1(_19840_),
    .B2(_20430_),
    .ZN(lce_data_cmd_o[111]));
 OAI21_X2 _47735_ (.A(_20435_),
    .B1(_20425_),
    .B2(\icache.lce.lce_cmd_inst.data_r [106]),
    .ZN(_20437_));
 AOI21_X4 _47736_ (.A(_20437_),
    .B1(_19844_),
    .B2(_20430_),
    .ZN(lce_data_cmd_o[112]));
 BUF_X8 _47737_ (.A(_20344_),
    .Z(_20438_));
 OAI21_X2 _47738_ (.A(_20435_),
    .B1(_20438_),
    .B2(\icache.lce.lce_cmd_inst.data_r [107]),
    .ZN(_20439_));
 AOI21_X4 _47739_ (.A(_20439_),
    .B1(_19848_),
    .B2(_20430_),
    .ZN(lce_data_cmd_o[113]));
 OAI21_X2 _47740_ (.A(_20435_),
    .B1(_20438_),
    .B2(\icache.lce.lce_cmd_inst.data_r [108]),
    .ZN(_20440_));
 AOI21_X4 _47741_ (.A(_20440_),
    .B1(_19853_),
    .B2(_20430_),
    .ZN(lce_data_cmd_o[114]));
 OAI21_X2 _47742_ (.A(_20435_),
    .B1(_20438_),
    .B2(\icache.lce.lce_cmd_inst.data_r [109]),
    .ZN(_20441_));
 AOI21_X4 _47743_ (.A(_20441_),
    .B1(_19857_),
    .B2(_20430_),
    .ZN(lce_data_cmd_o[115]));
 OAI21_X2 _47744_ (.A(_20435_),
    .B1(_20438_),
    .B2(\icache.lce.lce_cmd_inst.data_r [110]),
    .ZN(_20442_));
 BUF_X16 _47745_ (.A(_20364_),
    .Z(_20443_));
 AOI21_X4 _47746_ (.A(_20442_),
    .B1(_19861_),
    .B2(_20443_),
    .ZN(lce_data_cmd_o[116]));
 OAI21_X2 _47747_ (.A(_20435_),
    .B1(_20438_),
    .B2(\icache.lce.lce_cmd_inst.data_r [111]),
    .ZN(_20444_));
 AOI21_X4 _47748_ (.A(_20444_),
    .B1(_19866_),
    .B2(_20443_),
    .ZN(lce_data_cmd_o[117]));
 OAI21_X1 _47749_ (.A(_20435_),
    .B1(_20438_),
    .B2(\icache.lce.lce_cmd_inst.data_r [112]),
    .ZN(_20445_));
 AOI21_X4 _47750_ (.A(_20445_),
    .B1(_19870_),
    .B2(_20443_),
    .ZN(lce_data_cmd_o[118]));
 OAI21_X2 _47751_ (.A(_20435_),
    .B1(_20438_),
    .B2(\icache.lce.lce_cmd_inst.data_r [113]),
    .ZN(_20446_));
 AOI21_X4 _47752_ (.A(_20446_),
    .B1(_19874_),
    .B2(_20443_),
    .ZN(lce_data_cmd_o[119]));
 OAI21_X1 _47753_ (.A(_20435_),
    .B1(_20438_),
    .B2(\icache.lce.lce_cmd_inst.data_r [114]),
    .ZN(_20447_));
 AOI21_X4 _47754_ (.A(_20447_),
    .B1(_19878_),
    .B2(_20443_),
    .ZN(lce_data_cmd_o[120]));
 BUF_X16 _47755_ (.A(_20340_),
    .Z(_20448_));
 OAI21_X2 _47756_ (.A(_20448_),
    .B1(_20438_),
    .B2(\icache.lce.lce_cmd_inst.data_r [115]),
    .ZN(_20449_));
 AOI21_X4 _47757_ (.A(_20449_),
    .B1(_19882_),
    .B2(_20443_),
    .ZN(lce_data_cmd_o[121]));
 OAI21_X2 _47758_ (.A(_20448_),
    .B1(_20438_),
    .B2(\icache.lce.lce_cmd_inst.data_r [116]),
    .ZN(_20450_));
 AOI21_X4 _47759_ (.A(_20450_),
    .B1(_19473_),
    .B2(_20443_),
    .ZN(lce_data_cmd_o[122]));
 BUF_X16 _47760_ (.A(_20344_),
    .Z(_20451_));
 OAI21_X1 _47761_ (.A(_20448_),
    .B1(_20451_),
    .B2(\icache.lce.lce_cmd_inst.data_r [117]),
    .ZN(_20452_));
 AOI21_X4 _47762_ (.A(_20452_),
    .B1(_19478_),
    .B2(_20443_),
    .ZN(lce_data_cmd_o[123]));
 OAI21_X2 _47763_ (.A(_20448_),
    .B1(_20451_),
    .B2(\icache.lce.lce_cmd_inst.data_r [118]),
    .ZN(_20453_));
 AOI21_X4 _47764_ (.A(_20453_),
    .B1(_19482_),
    .B2(_20443_),
    .ZN(lce_data_cmd_o[124]));
 OAI21_X2 _47765_ (.A(_20448_),
    .B1(_20451_),
    .B2(\icache.lce.lce_cmd_inst.data_r [119]),
    .ZN(_20454_));
 AOI21_X4 _47766_ (.A(_20454_),
    .B1(_19486_),
    .B2(_20443_),
    .ZN(lce_data_cmd_o[125]));
 OAI21_X1 _47767_ (.A(_20448_),
    .B1(_20451_),
    .B2(\icache.lce.lce_cmd_inst.data_r [120]),
    .ZN(_20455_));
 BUF_X16 _47768_ (.A(_20364_),
    .Z(_20456_));
 AOI21_X4 _47769_ (.A(_20455_),
    .B1(_19490_),
    .B2(_20456_),
    .ZN(lce_data_cmd_o[126]));
 OAI21_X2 _47770_ (.A(_20448_),
    .B1(_20451_),
    .B2(\icache.lce.lce_cmd_inst.data_r [121]),
    .ZN(_20457_));
 AOI21_X4 _47771_ (.A(_20457_),
    .B1(_19494_),
    .B2(_20456_),
    .ZN(lce_data_cmd_o[127]));
 OAI21_X1 _47772_ (.A(_20448_),
    .B1(_20451_),
    .B2(\icache.lce.lce_cmd_inst.data_r [122]),
    .ZN(_20458_));
 AOI21_X4 _47773_ (.A(_20458_),
    .B1(_19498_),
    .B2(_20456_),
    .ZN(lce_data_cmd_o[128]));
 OAI21_X2 _47774_ (.A(_20448_),
    .B1(_20451_),
    .B2(\icache.lce.lce_cmd_inst.data_r [123]),
    .ZN(_20459_));
 AOI21_X4 _47775_ (.A(_20459_),
    .B1(_19502_),
    .B2(_20456_),
    .ZN(lce_data_cmd_o[129]));
 OAI21_X2 _47776_ (.A(_20448_),
    .B1(_20451_),
    .B2(\icache.lce.lce_cmd_inst.data_r [124]),
    .ZN(_20460_));
 AOI21_X4 _47777_ (.A(_20460_),
    .B1(_19508_),
    .B2(_20456_),
    .ZN(lce_data_cmd_o[130]));
 BUF_X16 _47778_ (.A(_20340_),
    .Z(_20461_));
 OAI21_X2 _47779_ (.A(_20461_),
    .B1(_20451_),
    .B2(\icache.lce.lce_cmd_inst.data_r [125]),
    .ZN(_20462_));
 AOI21_X4 _47780_ (.A(_20462_),
    .B1(_19513_),
    .B2(_20456_),
    .ZN(lce_data_cmd_o[131]));
 OAI21_X2 _47781_ (.A(_20461_),
    .B1(_20451_),
    .B2(\icache.lce.lce_cmd_inst.data_r [126]),
    .ZN(_20463_));
 AOI21_X4 _47782_ (.A(_20463_),
    .B1(_19517_),
    .B2(_20456_),
    .ZN(lce_data_cmd_o[132]));
 BUF_X8 _47783_ (.A(_20344_),
    .Z(_20464_));
 OAI21_X2 _47784_ (.A(_20461_),
    .B1(_20464_),
    .B2(\icache.lce.lce_cmd_inst.data_r [127]),
    .ZN(_20465_));
 AOI21_X4 _47785_ (.A(_20465_),
    .B1(_19522_),
    .B2(_20456_),
    .ZN(lce_data_cmd_o[133]));
 OAI21_X1 _47786_ (.A(_20461_),
    .B1(_20464_),
    .B2(\icache.lce.lce_cmd_inst.data_r [128]),
    .ZN(_20466_));
 AOI21_X4 _47787_ (.A(_20466_),
    .B1(_19527_),
    .B2(_20456_),
    .ZN(lce_data_cmd_o[134]));
 OAI21_X2 _47788_ (.A(_20461_),
    .B1(_20464_),
    .B2(\icache.lce.lce_cmd_inst.data_r [129]),
    .ZN(_20467_));
 AOI21_X4 _47789_ (.A(_20467_),
    .B1(_19531_),
    .B2(_20456_),
    .ZN(lce_data_cmd_o[135]));
 OAI21_X2 _47790_ (.A(_20461_),
    .B1(_20464_),
    .B2(\icache.lce.lce_cmd_inst.data_r [130]),
    .ZN(_20468_));
 BUF_X16 _47791_ (.A(_20364_),
    .Z(_20469_));
 AOI21_X4 _47792_ (.A(_20468_),
    .B1(_19535_),
    .B2(_20469_),
    .ZN(lce_data_cmd_o[136]));
 OAI21_X1 _47793_ (.A(_20461_),
    .B1(_20464_),
    .B2(\icache.lce.lce_cmd_inst.data_r [131]),
    .ZN(_20470_));
 AOI21_X4 _47794_ (.A(_20470_),
    .B1(_19539_),
    .B2(_20469_),
    .ZN(lce_data_cmd_o[137]));
 OAI21_X2 _47795_ (.A(_20461_),
    .B1(_20464_),
    .B2(\icache.lce.lce_cmd_inst.data_r [132]),
    .ZN(_20471_));
 AOI21_X4 _47796_ (.A(_20471_),
    .B1(_19543_),
    .B2(_20469_),
    .ZN(lce_data_cmd_o[138]));
 OAI21_X2 _47797_ (.A(_20461_),
    .B1(_20464_),
    .B2(\icache.lce.lce_cmd_inst.data_r [133]),
    .ZN(_20472_));
 AOI21_X4 _47798_ (.A(_20472_),
    .B1(_19547_),
    .B2(_20469_),
    .ZN(lce_data_cmd_o[139]));
 OAI21_X2 _47799_ (.A(_20461_),
    .B1(_20464_),
    .B2(\icache.lce.lce_cmd_inst.data_r [134]),
    .ZN(_20473_));
 AOI21_X4 _47800_ (.A(_20473_),
    .B1(_19552_),
    .B2(_20469_),
    .ZN(lce_data_cmd_o[140]));
 BUF_X16 _47801_ (.A(_07607_),
    .Z(_20474_));
 BUF_X8 _47802_ (.A(_20474_),
    .Z(_20475_));
 OAI21_X2 _47803_ (.A(_20475_),
    .B1(_20464_),
    .B2(\icache.lce.lce_cmd_inst.data_r [135]),
    .ZN(_20476_));
 AOI21_X4 _47804_ (.A(_20476_),
    .B1(_19556_),
    .B2(_20469_),
    .ZN(lce_data_cmd_o[141]));
 OAI21_X2 _47805_ (.A(_20475_),
    .B1(_20464_),
    .B2(\icache.lce.lce_cmd_inst.data_r [136]),
    .ZN(_20477_));
 AOI21_X4 _47806_ (.A(_20477_),
    .B1(_19560_),
    .B2(_20469_),
    .ZN(lce_data_cmd_o[142]));
 BUF_X16 _47807_ (.A(_15295_),
    .Z(_20478_));
 BUF_X8 _47808_ (.A(_20478_),
    .Z(_20479_));
 OAI21_X1 _47809_ (.A(_20475_),
    .B1(_20479_),
    .B2(\icache.lce.lce_cmd_inst.data_r [137]),
    .ZN(_20480_));
 AOI21_X4 _47810_ (.A(_20480_),
    .B1(_19565_),
    .B2(_20469_),
    .ZN(lce_data_cmd_o[143]));
 OAI21_X2 _47811_ (.A(_20475_),
    .B1(_20479_),
    .B2(\icache.lce.lce_cmd_inst.data_r [138]),
    .ZN(_20481_));
 AOI21_X4 _47812_ (.A(_20481_),
    .B1(_19569_),
    .B2(_20469_),
    .ZN(lce_data_cmd_o[144]));
 OAI21_X2 _47813_ (.A(_20475_),
    .B1(_20479_),
    .B2(\icache.lce.lce_cmd_inst.data_r [139]),
    .ZN(_20482_));
 AOI21_X4 _47814_ (.A(_20482_),
    .B1(_19573_),
    .B2(_20469_),
    .ZN(lce_data_cmd_o[145]));
 OAI21_X2 _47815_ (.A(_20475_),
    .B1(_20479_),
    .B2(\icache.lce.lce_cmd_inst.data_r [140]),
    .ZN(_20483_));
 BUF_X16 _47816_ (.A(_20364_),
    .Z(_20484_));
 AOI21_X4 _47817_ (.A(_20483_),
    .B1(_19577_),
    .B2(_20484_),
    .ZN(lce_data_cmd_o[146]));
 OAI21_X2 _47818_ (.A(_20475_),
    .B1(_20479_),
    .B2(\icache.lce.lce_cmd_inst.data_r [141]),
    .ZN(_20485_));
 AOI21_X4 _47819_ (.A(_20485_),
    .B1(_19582_),
    .B2(_20484_),
    .ZN(lce_data_cmd_o[147]));
 OAI21_X2 _47820_ (.A(_20475_),
    .B1(_20479_),
    .B2(\icache.lce.lce_cmd_inst.data_r [142]),
    .ZN(_20486_));
 AOI21_X4 _47821_ (.A(_20486_),
    .B1(_19586_),
    .B2(_20484_),
    .ZN(lce_data_cmd_o[148]));
 OAI21_X2 _47822_ (.A(_20475_),
    .B1(_20479_),
    .B2(\icache.lce.lce_cmd_inst.data_r [143]),
    .ZN(_20487_));
 AOI21_X4 _47823_ (.A(_20487_),
    .B1(_19590_),
    .B2(_20484_),
    .ZN(lce_data_cmd_o[149]));
 OAI21_X2 _47824_ (.A(_20475_),
    .B1(_20479_),
    .B2(\icache.lce.lce_cmd_inst.data_r [144]),
    .ZN(_20488_));
 AOI21_X4 _47825_ (.A(_20488_),
    .B1(_19597_),
    .B2(_20484_),
    .ZN(lce_data_cmd_o[150]));
 BUF_X4 _47826_ (.A(_20474_),
    .Z(_20489_));
 OAI21_X2 _47827_ (.A(_20489_),
    .B1(_20479_),
    .B2(\icache.lce.lce_cmd_inst.data_r [145]),
    .ZN(_20490_));
 AOI21_X4 _47828_ (.A(_20490_),
    .B1(_19601_),
    .B2(_20484_),
    .ZN(lce_data_cmd_o[151]));
 OAI21_X1 _47829_ (.A(_20489_),
    .B1(_20479_),
    .B2(\icache.lce.lce_cmd_inst.data_r [146]),
    .ZN(_20491_));
 AOI21_X4 _47830_ (.A(_20491_),
    .B1(_19605_),
    .B2(_20484_),
    .ZN(lce_data_cmd_o[152]));
 BUF_X4 _47831_ (.A(_20478_),
    .Z(_20492_));
 OAI21_X2 _47832_ (.A(_20489_),
    .B1(_20492_),
    .B2(\icache.lce.lce_cmd_inst.data_r [147]),
    .ZN(_20493_));
 AOI21_X4 _47833_ (.A(_20493_),
    .B1(_19610_),
    .B2(_20484_),
    .ZN(lce_data_cmd_o[153]));
 OAI21_X2 _47834_ (.A(_20489_),
    .B1(_20492_),
    .B2(\icache.lce.lce_cmd_inst.data_r [148]),
    .ZN(_20494_));
 AOI21_X4 _47835_ (.A(_20494_),
    .B1(_19614_),
    .B2(_20484_),
    .ZN(lce_data_cmd_o[154]));
 OAI21_X2 _47836_ (.A(_20489_),
    .B1(_20492_),
    .B2(\icache.lce.lce_cmd_inst.data_r [149]),
    .ZN(_20495_));
 AOI21_X4 _47837_ (.A(_20495_),
    .B1(_19618_),
    .B2(_20484_),
    .ZN(lce_data_cmd_o[155]));
 OAI21_X2 _47838_ (.A(_20489_),
    .B1(_20492_),
    .B2(\icache.lce.lce_cmd_inst.data_r [150]),
    .ZN(_20496_));
 BUF_X32 _47839_ (.A(_20363_),
    .Z(_20497_));
 BUF_X8 _47840_ (.A(_20497_),
    .Z(_20498_));
 AOI21_X4 _47841_ (.A(_20496_),
    .B1(_19622_),
    .B2(_20498_),
    .ZN(lce_data_cmd_o[156]));
 OAI21_X1 _47842_ (.A(_20489_),
    .B1(_20492_),
    .B2(\icache.lce.lce_cmd_inst.data_r [151]),
    .ZN(_20499_));
 AOI21_X4 _47843_ (.A(_20499_),
    .B1(_19626_),
    .B2(_20498_),
    .ZN(lce_data_cmd_o[157]));
 OAI21_X2 _47844_ (.A(_20489_),
    .B1(_20492_),
    .B2(\icache.lce.lce_cmd_inst.data_r [152]),
    .ZN(_20500_));
 AOI21_X4 _47845_ (.A(_20500_),
    .B1(_19630_),
    .B2(_20498_),
    .ZN(lce_data_cmd_o[158]));
 OAI21_X2 _47846_ (.A(_20489_),
    .B1(_20492_),
    .B2(\icache.lce.lce_cmd_inst.data_r [153]),
    .ZN(_20501_));
 AOI21_X4 _47847_ (.A(_20501_),
    .B1(_19634_),
    .B2(_20498_),
    .ZN(lce_data_cmd_o[159]));
 OAI21_X2 _47848_ (.A(_20489_),
    .B1(_20492_),
    .B2(\icache.lce.lce_cmd_inst.data_r [154]),
    .ZN(_20502_));
 AOI21_X4 _47849_ (.A(_20502_),
    .B1(_19640_),
    .B2(_20498_),
    .ZN(lce_data_cmd_o[160]));
 BUF_X8 _47850_ (.A(_20474_),
    .Z(_20503_));
 OAI21_X2 _47851_ (.A(_20503_),
    .B1(_20492_),
    .B2(\icache.lce.lce_cmd_inst.data_r [155]),
    .ZN(_20504_));
 AOI21_X4 _47852_ (.A(_20504_),
    .B1(_19644_),
    .B2(_20498_),
    .ZN(lce_data_cmd_o[161]));
 OAI21_X2 _47853_ (.A(_20503_),
    .B1(_20492_),
    .B2(\icache.lce.lce_cmd_inst.data_r [156]),
    .ZN(_20505_));
 AOI21_X4 _47854_ (.A(_20505_),
    .B1(_19648_),
    .B2(_20498_),
    .ZN(lce_data_cmd_o[162]));
 BUF_X8 _47855_ (.A(_20478_),
    .Z(_20506_));
 OAI21_X2 _47856_ (.A(_20503_),
    .B1(_20506_),
    .B2(\icache.lce.lce_cmd_inst.data_r [157]),
    .ZN(_20507_));
 AOI21_X4 _47857_ (.A(_20507_),
    .B1(_19654_),
    .B2(_20498_),
    .ZN(lce_data_cmd_o[163]));
 OAI21_X2 _47858_ (.A(_20503_),
    .B1(_20506_),
    .B2(\icache.lce.lce_cmd_inst.data_r [158]),
    .ZN(_20508_));
 AOI21_X4 _47859_ (.A(_20508_),
    .B1(_19658_),
    .B2(_20498_),
    .ZN(lce_data_cmd_o[164]));
 OAI21_X2 _47860_ (.A(_20503_),
    .B1(_20506_),
    .B2(\icache.lce.lce_cmd_inst.data_r [159]),
    .ZN(_20509_));
 AOI21_X4 _47861_ (.A(_20509_),
    .B1(_19662_),
    .B2(_20498_),
    .ZN(lce_data_cmd_o[165]));
 OAI21_X2 _47862_ (.A(_20503_),
    .B1(_20506_),
    .B2(\icache.lce.lce_cmd_inst.data_r [160]),
    .ZN(_20510_));
 BUF_X16 _47863_ (.A(_20497_),
    .Z(_20511_));
 AOI21_X4 _47864_ (.A(_20510_),
    .B1(_19666_),
    .B2(_20511_),
    .ZN(lce_data_cmd_o[166]));
 OAI21_X2 _47865_ (.A(_20503_),
    .B1(_20506_),
    .B2(\icache.lce.lce_cmd_inst.data_r [161]),
    .ZN(_20512_));
 AOI21_X4 _47866_ (.A(_20512_),
    .B1(_19670_),
    .B2(_20511_),
    .ZN(lce_data_cmd_o[167]));
 OAI21_X2 _47867_ (.A(_20503_),
    .B1(_20506_),
    .B2(\icache.lce.lce_cmd_inst.data_r [162]),
    .ZN(_20513_));
 AOI21_X4 _47868_ (.A(_20513_),
    .B1(_19674_),
    .B2(_20511_),
    .ZN(lce_data_cmd_o[168]));
 OAI21_X2 _47869_ (.A(_20503_),
    .B1(_20506_),
    .B2(\icache.lce.lce_cmd_inst.data_r [163]),
    .ZN(_20514_));
 AOI21_X4 _47870_ (.A(_20514_),
    .B1(_19678_),
    .B2(_20511_),
    .ZN(lce_data_cmd_o[169]));
 OAI21_X2 _47871_ (.A(_20503_),
    .B1(_20506_),
    .B2(\icache.lce.lce_cmd_inst.data_r [164]),
    .ZN(_20515_));
 AOI21_X4 _47872_ (.A(_20515_),
    .B1(_19684_),
    .B2(_20511_),
    .ZN(lce_data_cmd_o[170]));
 BUF_X8 _47873_ (.A(_20474_),
    .Z(_20516_));
 OAI21_X2 _47874_ (.A(_20516_),
    .B1(_20506_),
    .B2(\icache.lce.lce_cmd_inst.data_r [165]),
    .ZN(_20517_));
 AOI21_X4 _47875_ (.A(_20517_),
    .B1(_19688_),
    .B2(_20511_),
    .ZN(lce_data_cmd_o[171]));
 OAI21_X2 _47876_ (.A(_20516_),
    .B1(_20506_),
    .B2(\icache.lce.lce_cmd_inst.data_r [166]),
    .ZN(_20518_));
 AOI21_X4 _47877_ (.A(_20518_),
    .B1(_19692_),
    .B2(_20511_),
    .ZN(lce_data_cmd_o[172]));
 BUF_X8 _47878_ (.A(_20478_),
    .Z(_20519_));
 OAI21_X1 _47879_ (.A(_20516_),
    .B1(_20519_),
    .B2(\icache.lce.lce_cmd_inst.data_r [167]),
    .ZN(_20520_));
 AOI21_X4 _47880_ (.A(_20520_),
    .B1(_19698_),
    .B2(_20511_),
    .ZN(lce_data_cmd_o[173]));
 OAI21_X2 _47881_ (.A(_20516_),
    .B1(_20519_),
    .B2(\icache.lce.lce_cmd_inst.data_r [168]),
    .ZN(_20521_));
 AOI21_X4 _47882_ (.A(_20521_),
    .B1(_19702_),
    .B2(_20511_),
    .ZN(lce_data_cmd_o[174]));
 OAI21_X2 _47883_ (.A(_20516_),
    .B1(_20519_),
    .B2(\icache.lce.lce_cmd_inst.data_r [169]),
    .ZN(_20522_));
 AOI21_X4 _47884_ (.A(_20522_),
    .B1(_19706_),
    .B2(_20511_),
    .ZN(lce_data_cmd_o[175]));
 OAI21_X2 _47885_ (.A(_20516_),
    .B1(_20519_),
    .B2(\icache.lce.lce_cmd_inst.data_r [170]),
    .ZN(_20523_));
 BUF_X8 _47886_ (.A(_20497_),
    .Z(_20524_));
 AOI21_X4 _47887_ (.A(_20523_),
    .B1(_19710_),
    .B2(_20524_),
    .ZN(lce_data_cmd_o[176]));
 OAI21_X2 _47888_ (.A(_20516_),
    .B1(_20519_),
    .B2(\icache.lce.lce_cmd_inst.data_r [171]),
    .ZN(_20525_));
 AOI21_X4 _47889_ (.A(_20525_),
    .B1(_19714_),
    .B2(_20524_),
    .ZN(lce_data_cmd_o[177]));
 OAI21_X2 _47890_ (.A(_20516_),
    .B1(_20519_),
    .B2(\icache.lce.lce_cmd_inst.data_r [172]),
    .ZN(_20526_));
 AOI21_X4 _47891_ (.A(_20526_),
    .B1(_19718_),
    .B2(_20524_),
    .ZN(lce_data_cmd_o[178]));
 OAI21_X2 _47892_ (.A(_20516_),
    .B1(_20519_),
    .B2(\icache.lce.lce_cmd_inst.data_r [173]),
    .ZN(_20527_));
 AOI21_X4 _47893_ (.A(_20527_),
    .B1(_19722_),
    .B2(_20524_),
    .ZN(lce_data_cmd_o[179]));
 OAI21_X2 _47894_ (.A(_20516_),
    .B1(_20519_),
    .B2(\icache.lce.lce_cmd_inst.data_r [174]),
    .ZN(_20528_));
 AOI21_X4 _47895_ (.A(_20528_),
    .B1(_19727_),
    .B2(_20524_),
    .ZN(lce_data_cmd_o[180]));
 BUF_X8 _47896_ (.A(_20474_),
    .Z(_20529_));
 OAI21_X2 _47897_ (.A(_20529_),
    .B1(_20519_),
    .B2(\icache.lce.lce_cmd_inst.data_r [175]),
    .ZN(_20530_));
 AOI21_X4 _47898_ (.A(_20530_),
    .B1(_19731_),
    .B2(_20524_),
    .ZN(lce_data_cmd_o[181]));
 OAI21_X2 _47899_ (.A(_20529_),
    .B1(_20519_),
    .B2(\icache.lce.lce_cmd_inst.data_r [176]),
    .ZN(_20531_));
 AOI21_X4 _47900_ (.A(_20531_),
    .B1(_19735_),
    .B2(_20524_),
    .ZN(lce_data_cmd_o[182]));
 BUF_X4 _47901_ (.A(_20478_),
    .Z(_20532_));
 OAI21_X2 _47902_ (.A(_20529_),
    .B1(_20532_),
    .B2(\icache.lce.lce_cmd_inst.data_r [177]),
    .ZN(_20533_));
 AOI21_X4 _47903_ (.A(_20533_),
    .B1(_19740_),
    .B2(_20524_),
    .ZN(lce_data_cmd_o[183]));
 OAI21_X2 _47904_ (.A(_20529_),
    .B1(_20532_),
    .B2(\icache.lce.lce_cmd_inst.data_r [178]),
    .ZN(_20534_));
 AOI21_X4 _47905_ (.A(_20534_),
    .B1(_19744_),
    .B2(_20524_),
    .ZN(lce_data_cmd_o[184]));
 OAI21_X2 _47906_ (.A(_20529_),
    .B1(_20532_),
    .B2(\icache.lce.lce_cmd_inst.data_r [179]),
    .ZN(_20535_));
 AOI21_X4 _47907_ (.A(_20535_),
    .B1(_19748_),
    .B2(_20524_),
    .ZN(lce_data_cmd_o[185]));
 OAI21_X2 _47908_ (.A(_20529_),
    .B1(_20532_),
    .B2(\icache.lce.lce_cmd_inst.data_r [180]),
    .ZN(_20536_));
 BUF_X16 _47909_ (.A(_20497_),
    .Z(_20537_));
 AOI21_X4 _47910_ (.A(_20536_),
    .B1(_19752_),
    .B2(_20537_),
    .ZN(lce_data_cmd_o[186]));
 OAI21_X2 _47911_ (.A(_20529_),
    .B1(_20532_),
    .B2(\icache.lce.lce_cmd_inst.data_r [181]),
    .ZN(_20538_));
 AOI21_X4 _47912_ (.A(_20538_),
    .B1(_19756_),
    .B2(_20537_),
    .ZN(lce_data_cmd_o[187]));
 OAI21_X2 _47913_ (.A(_20529_),
    .B1(_20532_),
    .B2(\icache.lce.lce_cmd_inst.data_r [182]),
    .ZN(_20539_));
 AOI21_X4 _47914_ (.A(_20539_),
    .B1(_19760_),
    .B2(_20537_),
    .ZN(lce_data_cmd_o[188]));
 OAI21_X2 _47915_ (.A(_20529_),
    .B1(_20532_),
    .B2(\icache.lce.lce_cmd_inst.data_r [183]),
    .ZN(_20540_));
 AOI21_X4 _47916_ (.A(_20540_),
    .B1(_19764_),
    .B2(_20537_),
    .ZN(lce_data_cmd_o[189]));
 OAI21_X1 _47917_ (.A(_20529_),
    .B1(_20532_),
    .B2(\icache.lce.lce_cmd_inst.data_r [184]),
    .ZN(_20541_));
 AOI21_X4 _47918_ (.A(_20541_),
    .B1(_19769_),
    .B2(_20537_),
    .ZN(lce_data_cmd_o[190]));
 BUF_X16 _47919_ (.A(_20474_),
    .Z(_20542_));
 OAI21_X2 _47920_ (.A(_20542_),
    .B1(_20532_),
    .B2(\icache.lce.lce_cmd_inst.data_r [185]),
    .ZN(_20543_));
 AOI21_X4 _47921_ (.A(_20543_),
    .B1(_19773_),
    .B2(_20537_),
    .ZN(lce_data_cmd_o[191]));
 OAI21_X2 _47922_ (.A(_20542_),
    .B1(_20532_),
    .B2(\icache.lce.lce_cmd_inst.data_r [186]),
    .ZN(_20544_));
 AOI21_X4 _47923_ (.A(_20544_),
    .B1(_19777_),
    .B2(_20537_),
    .ZN(lce_data_cmd_o[192]));
 BUF_X8 _47924_ (.A(_20478_),
    .Z(_20545_));
 OAI21_X2 _47925_ (.A(_20542_),
    .B1(_20545_),
    .B2(\icache.lce.lce_cmd_inst.data_r [187]),
    .ZN(_20546_));
 AOI21_X4 _47926_ (.A(_20546_),
    .B1(_19782_),
    .B2(_20537_),
    .ZN(lce_data_cmd_o[193]));
 OAI21_X2 _47927_ (.A(_20542_),
    .B1(_20545_),
    .B2(\icache.lce.lce_cmd_inst.data_r [188]),
    .ZN(_20547_));
 AOI21_X4 _47928_ (.A(_20547_),
    .B1(_19786_),
    .B2(_20537_),
    .ZN(lce_data_cmd_o[194]));
 OAI21_X2 _47929_ (.A(_20542_),
    .B1(_20545_),
    .B2(\icache.lce.lce_cmd_inst.data_r [189]),
    .ZN(_20548_));
 AOI21_X4 _47930_ (.A(_20548_),
    .B1(_19790_),
    .B2(_20537_),
    .ZN(lce_data_cmd_o[195]));
 OAI21_X2 _47931_ (.A(_20542_),
    .B1(_20545_),
    .B2(\icache.lce.lce_cmd_inst.data_r [190]),
    .ZN(_20549_));
 BUF_X16 _47932_ (.A(_20497_),
    .Z(_20550_));
 AOI21_X4 _47933_ (.A(_20549_),
    .B1(_19794_),
    .B2(_20550_),
    .ZN(lce_data_cmd_o[196]));
 OAI21_X2 _47934_ (.A(_20542_),
    .B1(_20545_),
    .B2(\icache.lce.lce_cmd_inst.data_r [191]),
    .ZN(_20551_));
 AOI21_X4 _47935_ (.A(_20551_),
    .B1(_19798_),
    .B2(_20550_),
    .ZN(lce_data_cmd_o[197]));
 OAI21_X2 _47936_ (.A(_20542_),
    .B1(_20545_),
    .B2(\icache.lce.lce_cmd_inst.data_r [192]),
    .ZN(_20552_));
 AOI21_X4 _47937_ (.A(_20552_),
    .B1(_19802_),
    .B2(_20550_),
    .ZN(lce_data_cmd_o[198]));
 OAI21_X2 _47938_ (.A(_20542_),
    .B1(_20545_),
    .B2(\icache.lce.lce_cmd_inst.data_r [193]),
    .ZN(_20553_));
 AOI21_X4 _47939_ (.A(_20553_),
    .B1(_19460_),
    .B2(_20550_),
    .ZN(lce_data_cmd_o[199]));
 OAI21_X1 _47940_ (.A(_20542_),
    .B1(_20545_),
    .B2(\icache.lce.lce_cmd_inst.data_r [194]),
    .ZN(_20554_));
 AOI21_X4 _47941_ (.A(_20554_),
    .B1(_19465_),
    .B2(_20550_),
    .ZN(lce_data_cmd_o[200]));
 BUF_X8 _47942_ (.A(_20474_),
    .Z(_20555_));
 OAI21_X2 _47943_ (.A(_20555_),
    .B1(_20545_),
    .B2(\icache.lce.lce_cmd_inst.data_r [195]),
    .ZN(_20556_));
 AOI21_X4 _47944_ (.A(_20556_),
    .B1(_19469_),
    .B2(_20550_),
    .ZN(lce_data_cmd_o[201]));
 OAI21_X2 _47945_ (.A(_20555_),
    .B1(_20545_),
    .B2(\icache.lce.lce_cmd_inst.data_r [196]),
    .ZN(_20557_));
 AOI21_X4 _47946_ (.A(_20557_),
    .B1(_19379_),
    .B2(_20550_),
    .ZN(lce_data_cmd_o[202]));
 BUF_X8 _47947_ (.A(_20478_),
    .Z(_20558_));
 OAI21_X2 _47948_ (.A(_20555_),
    .B1(_20558_),
    .B2(\icache.lce.lce_cmd_inst.data_r [197]),
    .ZN(_20559_));
 AOI21_X4 _47949_ (.A(_20559_),
    .B1(_19383_),
    .B2(_20550_),
    .ZN(lce_data_cmd_o[203]));
 OAI21_X2 _47950_ (.A(_20555_),
    .B1(_20558_),
    .B2(\icache.lce.lce_cmd_inst.data_r [198]),
    .ZN(_20560_));
 AOI21_X4 _47951_ (.A(_20560_),
    .B1(_19387_),
    .B2(_20550_),
    .ZN(lce_data_cmd_o[204]));
 OAI21_X1 _47952_ (.A(_20555_),
    .B1(_20558_),
    .B2(\icache.lce.lce_cmd_inst.data_r [199]),
    .ZN(_20561_));
 AOI21_X4 _47953_ (.A(_20561_),
    .B1(_19392_),
    .B2(_20550_),
    .ZN(lce_data_cmd_o[205]));
 OAI21_X1 _47954_ (.A(_20555_),
    .B1(_20558_),
    .B2(\icache.lce.lce_cmd_inst.data_r [200]),
    .ZN(_20562_));
 BUF_X8 _47955_ (.A(_20497_),
    .Z(_20563_));
 AOI21_X4 _47956_ (.A(_20562_),
    .B1(_19396_),
    .B2(_20563_),
    .ZN(lce_data_cmd_o[206]));
 OAI21_X2 _47957_ (.A(_20555_),
    .B1(_20558_),
    .B2(\icache.lce.lce_cmd_inst.data_r [201]),
    .ZN(_20564_));
 AOI21_X4 _47958_ (.A(_20564_),
    .B1(_19401_),
    .B2(_20563_),
    .ZN(lce_data_cmd_o[207]));
 OAI21_X1 _47959_ (.A(_20555_),
    .B1(_20558_),
    .B2(\icache.lce.lce_cmd_inst.data_r [202]),
    .ZN(_20565_));
 AOI21_X4 _47960_ (.A(_20565_),
    .B1(_19405_),
    .B2(_20563_),
    .ZN(lce_data_cmd_o[208]));
 OAI21_X1 _47961_ (.A(_20555_),
    .B1(_20558_),
    .B2(\icache.lce.lce_cmd_inst.data_r [203]),
    .ZN(_20566_));
 AOI21_X4 _47962_ (.A(_20566_),
    .B1(_19409_),
    .B2(_20563_),
    .ZN(lce_data_cmd_o[209]));
 OAI21_X2 _47963_ (.A(_20555_),
    .B1(_20558_),
    .B2(\icache.lce.lce_cmd_inst.data_r [204]),
    .ZN(_20567_));
 AOI21_X4 _47964_ (.A(_20567_),
    .B1(_19413_),
    .B2(_20563_),
    .ZN(lce_data_cmd_o[210]));
 BUF_X8 _47965_ (.A(_20474_),
    .Z(_20568_));
 OAI21_X2 _47966_ (.A(_20568_),
    .B1(_20558_),
    .B2(\icache.lce.lce_cmd_inst.data_r [205]),
    .ZN(_20569_));
 AOI21_X4 _47967_ (.A(_20569_),
    .B1(_19417_),
    .B2(_20563_),
    .ZN(lce_data_cmd_o[211]));
 OAI21_X2 _47968_ (.A(_20568_),
    .B1(_20558_),
    .B2(\icache.lce.lce_cmd_inst.data_r [206]),
    .ZN(_20570_));
 AOI21_X4 _47969_ (.A(_20570_),
    .B1(_19422_),
    .B2(_20563_),
    .ZN(lce_data_cmd_o[212]));
 BUF_X8 _47970_ (.A(_20478_),
    .Z(_20571_));
 OAI21_X2 _47971_ (.A(_20568_),
    .B1(_20571_),
    .B2(\icache.lce.lce_cmd_inst.data_r [207]),
    .ZN(_20572_));
 AOI21_X4 _47972_ (.A(_20572_),
    .B1(_19427_),
    .B2(_20563_),
    .ZN(lce_data_cmd_o[213]));
 OAI21_X2 _47973_ (.A(_20568_),
    .B1(_20571_),
    .B2(\icache.lce.lce_cmd_inst.data_r [208]),
    .ZN(_20573_));
 AOI21_X4 _47974_ (.A(_20573_),
    .B1(_19431_),
    .B2(_20563_),
    .ZN(lce_data_cmd_o[214]));
 OAI21_X2 _47975_ (.A(_20568_),
    .B1(_20571_),
    .B2(\icache.lce.lce_cmd_inst.data_r [209]),
    .ZN(_20574_));
 AOI21_X4 _47976_ (.A(_20574_),
    .B1(_19436_),
    .B2(_20563_),
    .ZN(lce_data_cmd_o[215]));
 OAI21_X2 _47977_ (.A(_20568_),
    .B1(_20571_),
    .B2(\icache.lce.lce_cmd_inst.data_r [210]),
    .ZN(_20575_));
 BUF_X16 _47978_ (.A(_20497_),
    .Z(_20576_));
 AOI21_X4 _47979_ (.A(_20575_),
    .B1(_19440_),
    .B2(_20576_),
    .ZN(lce_data_cmd_o[216]));
 OAI21_X2 _47980_ (.A(_20568_),
    .B1(_20571_),
    .B2(\icache.lce.lce_cmd_inst.data_r [211]),
    .ZN(_20577_));
 AOI21_X4 _47981_ (.A(_20577_),
    .B1(_19444_),
    .B2(_20576_),
    .ZN(lce_data_cmd_o[217]));
 OAI21_X1 _47982_ (.A(_20568_),
    .B1(_20571_),
    .B2(\icache.lce.lce_cmd_inst.data_r [212]),
    .ZN(_20578_));
 AOI21_X4 _47983_ (.A(_20578_),
    .B1(_19448_),
    .B2(_20576_),
    .ZN(lce_data_cmd_o[218]));
 OAI21_X2 _47984_ (.A(_20568_),
    .B1(_20571_),
    .B2(\icache.lce.lce_cmd_inst.data_r [213]),
    .ZN(_20579_));
 AOI21_X4 _47985_ (.A(_20579_),
    .B1(_19452_),
    .B2(_20576_),
    .ZN(lce_data_cmd_o[219]));
 OAI21_X2 _47986_ (.A(_20568_),
    .B1(_20571_),
    .B2(\icache.lce.lce_cmd_inst.data_r [214]),
    .ZN(_20580_));
 AOI21_X4 _47987_ (.A(_20580_),
    .B1(_19456_),
    .B2(_20576_),
    .ZN(lce_data_cmd_o[220]));
 BUF_X8 _47988_ (.A(_20474_),
    .Z(_20581_));
 OAI21_X2 _47989_ (.A(_20581_),
    .B1(_20571_),
    .B2(\icache.lce.lce_cmd_inst.data_r [215]),
    .ZN(_20582_));
 AOI21_X4 _47990_ (.A(_20582_),
    .B1(_18885_),
    .B2(_20576_),
    .ZN(lce_data_cmd_o[221]));
 OAI21_X2 _47991_ (.A(_20581_),
    .B1(_20571_),
    .B2(\icache.lce.lce_cmd_inst.data_r [216]),
    .ZN(_20583_));
 AOI21_X4 _47992_ (.A(_20583_),
    .B1(_18889_),
    .B2(_20576_),
    .ZN(lce_data_cmd_o[222]));
 BUF_X8 _47993_ (.A(_20478_),
    .Z(_20584_));
 OAI21_X2 _47994_ (.A(_20581_),
    .B1(_20584_),
    .B2(\icache.lce.lce_cmd_inst.data_r [217]),
    .ZN(_20585_));
 AOI21_X4 _47995_ (.A(_20585_),
    .B1(_18893_),
    .B2(_20576_),
    .ZN(lce_data_cmd_o[223]));
 OAI21_X1 _47996_ (.A(_20581_),
    .B1(_20584_),
    .B2(\icache.lce.lce_cmd_inst.data_r [218]),
    .ZN(_20586_));
 AOI21_X4 _47997_ (.A(_20586_),
    .B1(_18897_),
    .B2(_20576_),
    .ZN(lce_data_cmd_o[224]));
 OAI21_X2 _47998_ (.A(_20581_),
    .B1(_20584_),
    .B2(\icache.lce.lce_cmd_inst.data_r [219]),
    .ZN(_20587_));
 AOI21_X4 _47999_ (.A(_20587_),
    .B1(_18901_),
    .B2(_20576_),
    .ZN(lce_data_cmd_o[225]));
 OAI21_X2 _48000_ (.A(_20581_),
    .B1(_20584_),
    .B2(\icache.lce.lce_cmd_inst.data_r [220]),
    .ZN(_20588_));
 BUF_X8 _48001_ (.A(_20497_),
    .Z(_20589_));
 AOI21_X4 _48002_ (.A(_20588_),
    .B1(_18906_),
    .B2(_20589_),
    .ZN(lce_data_cmd_o[226]));
 OAI21_X2 _48003_ (.A(_20581_),
    .B1(_20584_),
    .B2(\icache.lce.lce_cmd_inst.data_r [221]),
    .ZN(_20590_));
 AOI21_X4 _48004_ (.A(_20590_),
    .B1(_18910_),
    .B2(_20589_),
    .ZN(lce_data_cmd_o[227]));
 OAI21_X2 _48005_ (.A(_20581_),
    .B1(_20584_),
    .B2(\icache.lce.lce_cmd_inst.data_r [222]),
    .ZN(_20591_));
 AOI21_X4 _48006_ (.A(_20591_),
    .B1(_18915_),
    .B2(_20589_),
    .ZN(lce_data_cmd_o[228]));
 OAI21_X2 _48007_ (.A(_20581_),
    .B1(_20584_),
    .B2(\icache.lce.lce_cmd_inst.data_r [223]),
    .ZN(_20592_));
 AOI21_X4 _48008_ (.A(_20592_),
    .B1(_18920_),
    .B2(_20589_),
    .ZN(lce_data_cmd_o[229]));
 OAI21_X2 _48009_ (.A(_20581_),
    .B1(_20584_),
    .B2(\icache.lce.lce_cmd_inst.data_r [224]),
    .ZN(_20593_));
 AOI21_X4 _48010_ (.A(_20593_),
    .B1(_18925_),
    .B2(_20589_),
    .ZN(lce_data_cmd_o[230]));
 BUF_X8 _48011_ (.A(_20474_),
    .Z(_20594_));
 OAI21_X2 _48012_ (.A(_20594_),
    .B1(_20584_),
    .B2(\icache.lce.lce_cmd_inst.data_r [225]),
    .ZN(_20595_));
 AOI21_X4 _48013_ (.A(_20595_),
    .B1(_18930_),
    .B2(_20589_),
    .ZN(lce_data_cmd_o[231]));
 OAI21_X2 _48014_ (.A(_20594_),
    .B1(_20584_),
    .B2(\icache.lce.lce_cmd_inst.data_r [226]),
    .ZN(_20596_));
 AOI21_X4 _48015_ (.A(_20596_),
    .B1(_18934_),
    .B2(_20589_),
    .ZN(lce_data_cmd_o[232]));
 BUF_X16 _48016_ (.A(_20478_),
    .Z(_20597_));
 OAI21_X2 _48017_ (.A(_20594_),
    .B1(_20597_),
    .B2(\icache.lce.lce_cmd_inst.data_r [227]),
    .ZN(_20598_));
 AOI21_X4 _48018_ (.A(_20598_),
    .B1(_18938_),
    .B2(_20589_),
    .ZN(lce_data_cmd_o[233]));
 OAI21_X2 _48019_ (.A(_20594_),
    .B1(_20597_),
    .B2(\icache.lce.lce_cmd_inst.data_r [228]),
    .ZN(_20599_));
 AOI21_X4 _48020_ (.A(_20599_),
    .B1(_18942_),
    .B2(_20589_),
    .ZN(lce_data_cmd_o[234]));
 OAI21_X2 _48021_ (.A(_20594_),
    .B1(_20597_),
    .B2(\icache.lce.lce_cmd_inst.data_r [229]),
    .ZN(_20600_));
 AOI21_X4 _48022_ (.A(_20600_),
    .B1(_18946_),
    .B2(_20589_),
    .ZN(lce_data_cmd_o[235]));
 OAI21_X2 _48023_ (.A(_20594_),
    .B1(_20597_),
    .B2(\icache.lce.lce_cmd_inst.data_r [230]),
    .ZN(_20601_));
 BUF_X16 _48024_ (.A(_20497_),
    .Z(_20602_));
 AOI21_X4 _48025_ (.A(_20601_),
    .B1(_18950_),
    .B2(_20602_),
    .ZN(lce_data_cmd_o[236]));
 OAI21_X2 _48026_ (.A(_20594_),
    .B1(_20597_),
    .B2(\icache.lce.lce_cmd_inst.data_r [231]),
    .ZN(_20603_));
 AOI21_X4 _48027_ (.A(_20603_),
    .B1(_18954_),
    .B2(_20602_),
    .ZN(lce_data_cmd_o[237]));
 OAI21_X2 _48028_ (.A(_20594_),
    .B1(_20597_),
    .B2(\icache.lce.lce_cmd_inst.data_r [232]),
    .ZN(_20604_));
 AOI21_X4 _48029_ (.A(_20604_),
    .B1(_18959_),
    .B2(_20602_),
    .ZN(lce_data_cmd_o[238]));
 OAI21_X2 _48030_ (.A(_20594_),
    .B1(_20597_),
    .B2(\icache.lce.lce_cmd_inst.data_r [233]),
    .ZN(_20605_));
 AOI21_X4 _48031_ (.A(_20605_),
    .B1(_18963_),
    .B2(_20602_),
    .ZN(lce_data_cmd_o[239]));
 OAI21_X2 _48032_ (.A(_20594_),
    .B1(_20597_),
    .B2(\icache.lce.lce_cmd_inst.data_r [234]),
    .ZN(_20606_));
 AOI21_X4 _48033_ (.A(_20606_),
    .B1(_18967_),
    .B2(_20602_),
    .ZN(lce_data_cmd_o[240]));
 BUF_X32 _48034_ (.A(_07607_),
    .Z(_20607_));
 BUF_X8 _48035_ (.A(_20607_),
    .Z(_20608_));
 OAI21_X2 _48036_ (.A(_20608_),
    .B1(_20597_),
    .B2(\icache.lce.lce_cmd_inst.data_r [235]),
    .ZN(_20609_));
 AOI21_X4 _48037_ (.A(_20609_),
    .B1(_18972_),
    .B2(_20602_),
    .ZN(lce_data_cmd_o[241]));
 OAI21_X2 _48038_ (.A(_20608_),
    .B1(_20597_),
    .B2(\icache.lce.lce_cmd_inst.data_r [236]),
    .ZN(_20610_));
 AOI21_X4 _48039_ (.A(_20610_),
    .B1(_18976_),
    .B2(_20602_),
    .ZN(lce_data_cmd_o[242]));
 BUF_X32 _48040_ (.A(_15295_),
    .Z(_20611_));
 BUF_X8 _48041_ (.A(_20611_),
    .Z(_20612_));
 OAI21_X2 _48042_ (.A(_20608_),
    .B1(_20612_),
    .B2(\icache.lce.lce_cmd_inst.data_r [237]),
    .ZN(_20613_));
 AOI21_X4 _48043_ (.A(_20613_),
    .B1(_18980_),
    .B2(_20602_),
    .ZN(lce_data_cmd_o[243]));
 OAI21_X2 _48044_ (.A(_20608_),
    .B1(_20612_),
    .B2(\icache.lce.lce_cmd_inst.data_r [238]),
    .ZN(_20614_));
 AOI21_X4 _48045_ (.A(_20614_),
    .B1(_18984_),
    .B2(_20602_),
    .ZN(lce_data_cmd_o[244]));
 OAI21_X2 _48046_ (.A(_20608_),
    .B1(_20612_),
    .B2(\icache.lce.lce_cmd_inst.data_r [239]),
    .ZN(_20615_));
 AOI21_X4 _48047_ (.A(_20615_),
    .B1(_18988_),
    .B2(_20602_),
    .ZN(lce_data_cmd_o[245]));
 OAI21_X1 _48048_ (.A(_20608_),
    .B1(_20612_),
    .B2(\icache.lce.lce_cmd_inst.data_r [240]),
    .ZN(_20616_));
 BUF_X16 _48049_ (.A(_20497_),
    .Z(_20617_));
 AOI21_X4 _48050_ (.A(_20616_),
    .B1(_18992_),
    .B2(_20617_),
    .ZN(lce_data_cmd_o[246]));
 OAI21_X1 _48051_ (.A(_20608_),
    .B1(_20612_),
    .B2(\icache.lce.lce_cmd_inst.data_r [241]),
    .ZN(_20618_));
 AOI21_X4 _48052_ (.A(_20618_),
    .B1(_18996_),
    .B2(_20617_),
    .ZN(lce_data_cmd_o[247]));
 OAI21_X2 _48053_ (.A(_20608_),
    .B1(_20612_),
    .B2(\icache.lce.lce_cmd_inst.data_r [242]),
    .ZN(_20619_));
 AOI21_X4 _48054_ (.A(_20619_),
    .B1(_19002_),
    .B2(_20617_),
    .ZN(lce_data_cmd_o[248]));
 OAI21_X2 _48055_ (.A(_20608_),
    .B1(_20612_),
    .B2(\icache.lce.lce_cmd_inst.data_r [243]),
    .ZN(_20620_));
 AOI21_X4 _48056_ (.A(_20620_),
    .B1(_19007_),
    .B2(_20617_),
    .ZN(lce_data_cmd_o[249]));
 OAI21_X2 _48057_ (.A(_20608_),
    .B1(_20612_),
    .B2(\icache.lce.lce_cmd_inst.data_r [244]),
    .ZN(_20621_));
 AOI21_X4 _48058_ (.A(_20621_),
    .B1(_19011_),
    .B2(_20617_),
    .ZN(lce_data_cmd_o[250]));
 BUF_X16 _48059_ (.A(_20607_),
    .Z(_20622_));
 OAI21_X2 _48060_ (.A(_20622_),
    .B1(_20612_),
    .B2(\icache.lce.lce_cmd_inst.data_r [245]),
    .ZN(_20623_));
 AOI21_X4 _48061_ (.A(_20623_),
    .B1(_19016_),
    .B2(_20617_),
    .ZN(lce_data_cmd_o[251]));
 OAI21_X2 _48062_ (.A(_20622_),
    .B1(_20612_),
    .B2(\icache.lce.lce_cmd_inst.data_r [246]),
    .ZN(_20624_));
 AOI21_X4 _48063_ (.A(_20624_),
    .B1(_19020_),
    .B2(_20617_),
    .ZN(lce_data_cmd_o[252]));
 BUF_X8 _48064_ (.A(_20611_),
    .Z(_20625_));
 OAI21_X2 _48065_ (.A(_20622_),
    .B1(_20625_),
    .B2(\icache.lce.lce_cmd_inst.data_r [247]),
    .ZN(_20626_));
 AOI21_X4 _48066_ (.A(_20626_),
    .B1(_19024_),
    .B2(_20617_),
    .ZN(lce_data_cmd_o[253]));
 OAI21_X1 _48067_ (.A(_20622_),
    .B1(_20625_),
    .B2(\icache.lce.lce_cmd_inst.data_r [248]),
    .ZN(_20627_));
 AOI21_X4 _48068_ (.A(_20627_),
    .B1(_19028_),
    .B2(_20617_),
    .ZN(lce_data_cmd_o[254]));
 OAI21_X2 _48069_ (.A(_20622_),
    .B1(_20625_),
    .B2(\icache.lce.lce_cmd_inst.data_r [249]),
    .ZN(_20628_));
 AOI21_X4 _48070_ (.A(_20628_),
    .B1(_19032_),
    .B2(_20617_),
    .ZN(lce_data_cmd_o[255]));
 OAI21_X2 _48071_ (.A(_20622_),
    .B1(_20625_),
    .B2(\icache.lce.lce_cmd_inst.data_r [250]),
    .ZN(_20629_));
 BUF_X32 _48072_ (.A(_20363_),
    .Z(_20630_));
 BUF_X8 _48073_ (.A(_20630_),
    .Z(_20631_));
 AOI21_X4 _48074_ (.A(_20629_),
    .B1(_19037_),
    .B2(_20631_),
    .ZN(lce_data_cmd_o[256]));
 OAI21_X2 _48075_ (.A(_20622_),
    .B1(_20625_),
    .B2(\icache.lce.lce_cmd_inst.data_r [251]),
    .ZN(_20632_));
 AOI21_X4 _48076_ (.A(_20632_),
    .B1(_19041_),
    .B2(_20631_),
    .ZN(lce_data_cmd_o[257]));
 OAI21_X2 _48077_ (.A(_20622_),
    .B1(_20625_),
    .B2(\icache.lce.lce_cmd_inst.data_r [252]),
    .ZN(_20633_));
 AOI21_X4 _48078_ (.A(_20633_),
    .B1(_19047_),
    .B2(_20631_),
    .ZN(lce_data_cmd_o[258]));
 OAI21_X1 _48079_ (.A(_20622_),
    .B1(_20625_),
    .B2(\icache.lce.lce_cmd_inst.data_r [253]),
    .ZN(_20634_));
 AOI21_X4 _48080_ (.A(_20634_),
    .B1(_19051_),
    .B2(_20631_),
    .ZN(lce_data_cmd_o[259]));
 OAI21_X2 _48081_ (.A(_20622_),
    .B1(_20625_),
    .B2(\icache.lce.lce_cmd_inst.data_r [254]),
    .ZN(_20635_));
 AOI21_X4 _48082_ (.A(_20635_),
    .B1(_19055_),
    .B2(_20631_),
    .ZN(lce_data_cmd_o[260]));
 BUF_X8 _48083_ (.A(_20607_),
    .Z(_20636_));
 OAI21_X2 _48084_ (.A(_20636_),
    .B1(_20625_),
    .B2(\icache.lce.lce_cmd_inst.data_r [255]),
    .ZN(_20637_));
 AOI21_X4 _48085_ (.A(_20637_),
    .B1(_19061_),
    .B2(_20631_),
    .ZN(lce_data_cmd_o[261]));
 OAI21_X2 _48086_ (.A(_20636_),
    .B1(_20625_),
    .B2(\icache.lce.lce_cmd_inst.data_r [256]),
    .ZN(_20638_));
 AOI21_X4 _48087_ (.A(_20638_),
    .B1(_19065_),
    .B2(_20631_),
    .ZN(lce_data_cmd_o[262]));
 BUF_X8 _48088_ (.A(_20611_),
    .Z(_20639_));
 OAI21_X2 _48089_ (.A(_20636_),
    .B1(_20639_),
    .B2(\icache.lce.lce_cmd_inst.data_r [257]),
    .ZN(_20640_));
 AOI21_X4 _48090_ (.A(_20640_),
    .B1(_19074_),
    .B2(_20631_),
    .ZN(lce_data_cmd_o[263]));
 OAI21_X2 _48091_ (.A(_20636_),
    .B1(_20639_),
    .B2(\icache.lce.lce_cmd_inst.data_r [258]),
    .ZN(_20641_));
 AOI21_X4 _48092_ (.A(_20641_),
    .B1(_19082_),
    .B2(_20631_),
    .ZN(lce_data_cmd_o[264]));
 OAI21_X2 _48093_ (.A(_20636_),
    .B1(_20639_),
    .B2(\icache.lce.lce_cmd_inst.data_r [259]),
    .ZN(_20642_));
 AOI21_X4 _48094_ (.A(_20642_),
    .B1(_19092_),
    .B2(_20631_),
    .ZN(lce_data_cmd_o[265]));
 OAI21_X2 _48095_ (.A(_20636_),
    .B1(_20639_),
    .B2(\icache.lce.lce_cmd_inst.data_r [260]),
    .ZN(_20643_));
 BUF_X8 _48096_ (.A(_20630_),
    .Z(_20644_));
 AOI21_X4 _48097_ (.A(_20643_),
    .B1(_19101_),
    .B2(_20644_),
    .ZN(lce_data_cmd_o[266]));
 OAI21_X1 _48098_ (.A(_20636_),
    .B1(_20639_),
    .B2(\icache.lce.lce_cmd_inst.data_r [261]),
    .ZN(_20645_));
 AOI21_X4 _48099_ (.A(_20645_),
    .B1(_19109_),
    .B2(_20644_),
    .ZN(lce_data_cmd_o[267]));
 OAI21_X2 _48100_ (.A(_20636_),
    .B1(_20639_),
    .B2(\icache.lce.lce_cmd_inst.data_r [262]),
    .ZN(_20646_));
 AOI21_X4 _48101_ (.A(_20646_),
    .B1(_19118_),
    .B2(_20644_),
    .ZN(lce_data_cmd_o[268]));
 OAI21_X2 _48102_ (.A(_20636_),
    .B1(_20639_),
    .B2(\icache.lce.lce_cmd_inst.data_r [263]),
    .ZN(_20647_));
 AOI21_X4 _48103_ (.A(_20647_),
    .B1(_19127_),
    .B2(_20644_),
    .ZN(lce_data_cmd_o[269]));
 OAI21_X2 _48104_ (.A(_20636_),
    .B1(_20639_),
    .B2(\icache.lce.lce_cmd_inst.data_r [264]),
    .ZN(_20648_));
 AOI21_X4 _48105_ (.A(_20648_),
    .B1(_19135_),
    .B2(_20644_),
    .ZN(lce_data_cmd_o[270]));
 BUF_X4 _48106_ (.A(_20607_),
    .Z(_20649_));
 OAI21_X2 _48107_ (.A(_20649_),
    .B1(_20639_),
    .B2(\icache.lce.lce_cmd_inst.data_r [265]),
    .ZN(_20650_));
 AOI21_X4 _48108_ (.A(_20650_),
    .B1(_19144_),
    .B2(_20644_),
    .ZN(lce_data_cmd_o[271]));
 OAI21_X2 _48109_ (.A(_20649_),
    .B1(_20639_),
    .B2(\icache.lce.lce_cmd_inst.data_r [266]),
    .ZN(_20651_));
 AOI21_X4 _48110_ (.A(_20651_),
    .B1(_19152_),
    .B2(_20644_),
    .ZN(lce_data_cmd_o[272]));
 BUF_X4 _48111_ (.A(_20611_),
    .Z(_20652_));
 OAI21_X2 _48112_ (.A(_20649_),
    .B1(_20652_),
    .B2(\icache.lce.lce_cmd_inst.data_r [267]),
    .ZN(_20653_));
 AOI21_X4 _48113_ (.A(_20653_),
    .B1(_19161_),
    .B2(_20644_),
    .ZN(lce_data_cmd_o[273]));
 OAI21_X2 _48114_ (.A(_20649_),
    .B1(_20652_),
    .B2(\icache.lce.lce_cmd_inst.data_r [268]),
    .ZN(_20654_));
 AOI21_X4 _48115_ (.A(_20654_),
    .B1(_19169_),
    .B2(_20644_),
    .ZN(lce_data_cmd_o[274]));
 OAI21_X1 _48116_ (.A(_20649_),
    .B1(_20652_),
    .B2(\icache.lce.lce_cmd_inst.data_r [269]),
    .ZN(_20655_));
 AOI21_X4 _48117_ (.A(_20655_),
    .B1(_19177_),
    .B2(_20644_),
    .ZN(lce_data_cmd_o[275]));
 OAI21_X1 _48118_ (.A(_20649_),
    .B1(_20652_),
    .B2(\icache.lce.lce_cmd_inst.data_r [270]),
    .ZN(_20656_));
 BUF_X8 _48119_ (.A(_20630_),
    .Z(_20657_));
 AOI21_X4 _48120_ (.A(_20656_),
    .B1(_19188_),
    .B2(_20657_),
    .ZN(lce_data_cmd_o[276]));
 OAI21_X2 _48121_ (.A(_20649_),
    .B1(_20652_),
    .B2(\icache.lce.lce_cmd_inst.data_r [271]),
    .ZN(_20658_));
 AOI21_X4 _48122_ (.A(_20658_),
    .B1(_19196_),
    .B2(_20657_),
    .ZN(lce_data_cmd_o[277]));
 OAI21_X2 _48123_ (.A(_20649_),
    .B1(_20652_),
    .B2(\icache.lce.lce_cmd_inst.data_r [272]),
    .ZN(_20659_));
 AOI21_X4 _48124_ (.A(_20659_),
    .B1(_19205_),
    .B2(_20657_),
    .ZN(lce_data_cmd_o[278]));
 OAI21_X2 _48125_ (.A(_20649_),
    .B1(_20652_),
    .B2(\icache.lce.lce_cmd_inst.data_r [273]),
    .ZN(_20660_));
 AOI21_X4 _48126_ (.A(_20660_),
    .B1(_19214_),
    .B2(_20657_),
    .ZN(lce_data_cmd_o[279]));
 OAI21_X2 _48127_ (.A(_20649_),
    .B1(_20652_),
    .B2(\icache.lce.lce_cmd_inst.data_r [274]),
    .ZN(_20661_));
 AOI21_X4 _48128_ (.A(_20661_),
    .B1(_19223_),
    .B2(_20657_),
    .ZN(lce_data_cmd_o[280]));
 BUF_X4 _48129_ (.A(_20607_),
    .Z(_20662_));
 OAI21_X1 _48130_ (.A(_20662_),
    .B1(_20652_),
    .B2(\icache.lce.lce_cmd_inst.data_r [275]),
    .ZN(_20663_));
 AOI21_X4 _48131_ (.A(_20663_),
    .B1(_19232_),
    .B2(_20657_),
    .ZN(lce_data_cmd_o[281]));
 OAI21_X2 _48132_ (.A(_20662_),
    .B1(_20652_),
    .B2(\icache.lce.lce_cmd_inst.data_r [276]),
    .ZN(_20664_));
 AOI21_X4 _48133_ (.A(_20664_),
    .B1(_19241_),
    .B2(_20657_),
    .ZN(lce_data_cmd_o[282]));
 BUF_X4 _48134_ (.A(_20611_),
    .Z(_20665_));
 OAI21_X2 _48135_ (.A(_20662_),
    .B1(_20665_),
    .B2(\icache.lce.lce_cmd_inst.data_r [277]),
    .ZN(_20666_));
 AOI21_X4 _48136_ (.A(_20666_),
    .B1(_19251_),
    .B2(_20657_),
    .ZN(lce_data_cmd_o[283]));
 OAI21_X2 _48137_ (.A(_20662_),
    .B1(_20665_),
    .B2(\icache.lce.lce_cmd_inst.data_r [278]),
    .ZN(_20667_));
 AOI21_X4 _48138_ (.A(_20667_),
    .B1(_19259_),
    .B2(_20657_),
    .ZN(lce_data_cmd_o[284]));
 OAI21_X2 _48139_ (.A(_20662_),
    .B1(_20665_),
    .B2(\icache.lce.lce_cmd_inst.data_r [279]),
    .ZN(_20668_));
 AOI21_X4 _48140_ (.A(_20668_),
    .B1(_19267_),
    .B2(_20657_),
    .ZN(lce_data_cmd_o[285]));
 OAI21_X2 _48141_ (.A(_20662_),
    .B1(_20665_),
    .B2(\icache.lce.lce_cmd_inst.data_r [280]),
    .ZN(_20669_));
 BUF_X8 _48142_ (.A(_20630_),
    .Z(_20670_));
 AOI21_X4 _48143_ (.A(_20669_),
    .B1(_19275_),
    .B2(_20670_),
    .ZN(lce_data_cmd_o[286]));
 OAI21_X2 _48144_ (.A(_20662_),
    .B1(_20665_),
    .B2(\icache.lce.lce_cmd_inst.data_r [281]),
    .ZN(_20671_));
 AOI21_X4 _48145_ (.A(_20671_),
    .B1(_19283_),
    .B2(_20670_),
    .ZN(lce_data_cmd_o[287]));
 OAI21_X2 _48146_ (.A(_20662_),
    .B1(_20665_),
    .B2(\icache.lce.lce_cmd_inst.data_r [282]),
    .ZN(_20672_));
 AOI21_X4 _48147_ (.A(_20672_),
    .B1(_19292_),
    .B2(_20670_),
    .ZN(lce_data_cmd_o[288]));
 OAI21_X2 _48148_ (.A(_20662_),
    .B1(_20665_),
    .B2(\icache.lce.lce_cmd_inst.data_r [283]),
    .ZN(_20673_));
 AOI21_X4 _48149_ (.A(_20673_),
    .B1(_19300_),
    .B2(_20670_),
    .ZN(lce_data_cmd_o[289]));
 OAI21_X2 _48150_ (.A(_20662_),
    .B1(_20665_),
    .B2(\icache.lce.lce_cmd_inst.data_r [284]),
    .ZN(_20674_));
 AOI21_X4 _48151_ (.A(_20674_),
    .B1(_19310_),
    .B2(_20670_),
    .ZN(lce_data_cmd_o[290]));
 BUF_X8 _48152_ (.A(_20607_),
    .Z(_20675_));
 OAI21_X2 _48153_ (.A(_20675_),
    .B1(_20665_),
    .B2(\icache.lce.lce_cmd_inst.data_r [285]),
    .ZN(_20676_));
 AOI21_X4 _48154_ (.A(_20676_),
    .B1(_19319_),
    .B2(_20670_),
    .ZN(lce_data_cmd_o[291]));
 OAI21_X2 _48155_ (.A(_20675_),
    .B1(_20665_),
    .B2(\icache.lce.lce_cmd_inst.data_r [286]),
    .ZN(_20677_));
 AOI21_X4 _48156_ (.A(_20677_),
    .B1(_19328_),
    .B2(_20670_),
    .ZN(lce_data_cmd_o[292]));
 BUF_X16 _48157_ (.A(_20611_),
    .Z(_20678_));
 OAI21_X2 _48158_ (.A(_20675_),
    .B1(_20678_),
    .B2(\icache.lce.lce_cmd_inst.data_r [287]),
    .ZN(_20679_));
 AOI21_X4 _48159_ (.A(_20679_),
    .B1(_19338_),
    .B2(_20670_),
    .ZN(lce_data_cmd_o[293]));
 OAI21_X1 _48160_ (.A(_20675_),
    .B1(_20678_),
    .B2(\icache.lce.lce_cmd_inst.data_r [288]),
    .ZN(_20680_));
 AOI21_X4 _48161_ (.A(_20680_),
    .B1(_19346_),
    .B2(_20670_),
    .ZN(lce_data_cmd_o[294]));
 OAI21_X1 _48162_ (.A(_20675_),
    .B1(_20678_),
    .B2(\icache.lce.lce_cmd_inst.data_r [289]),
    .ZN(_20681_));
 AOI21_X4 _48163_ (.A(_20681_),
    .B1(_19355_),
    .B2(_20670_),
    .ZN(lce_data_cmd_o[295]));
 OAI21_X2 _48164_ (.A(_20675_),
    .B1(_20678_),
    .B2(\icache.lce.lce_cmd_inst.data_r [290]),
    .ZN(_20682_));
 BUF_X16 _48165_ (.A(_20630_),
    .Z(_20683_));
 AOI21_X4 _48166_ (.A(_20682_),
    .B1(_19364_),
    .B2(_20683_),
    .ZN(lce_data_cmd_o[296]));
 OAI21_X2 _48167_ (.A(_20675_),
    .B1(_20678_),
    .B2(\icache.lce.lce_cmd_inst.data_r [291]),
    .ZN(_20684_));
 AOI21_X4 _48168_ (.A(_20684_),
    .B1(_19374_),
    .B2(_20683_),
    .ZN(lce_data_cmd_o[297]));
 OAI21_X2 _48169_ (.A(_20675_),
    .B1(_20678_),
    .B2(\icache.lce.lce_cmd_inst.data_r [292]),
    .ZN(_20685_));
 AOI21_X4 _48170_ (.A(_20685_),
    .B1(_18862_),
    .B2(_20683_),
    .ZN(lce_data_cmd_o[298]));
 OAI21_X2 _48171_ (.A(_20675_),
    .B1(_20678_),
    .B2(\icache.lce.lce_cmd_inst.data_r [293]),
    .ZN(_20686_));
 AOI21_X4 _48172_ (.A(_20686_),
    .B1(_18871_),
    .B2(_20683_),
    .ZN(lce_data_cmd_o[299]));
 OAI21_X1 _48173_ (.A(_20675_),
    .B1(_20678_),
    .B2(\icache.lce.lce_cmd_inst.data_r [294]),
    .ZN(_20687_));
 AOI21_X4 _48174_ (.A(_20687_),
    .B1(_18880_),
    .B2(_20683_),
    .ZN(lce_data_cmd_o[300]));
 BUF_X8 _48175_ (.A(_20607_),
    .Z(_20688_));
 OAI21_X2 _48176_ (.A(_20688_),
    .B1(_20678_),
    .B2(\icache.lce.lce_cmd_inst.data_r [295]),
    .ZN(_20689_));
 AOI21_X4 _48177_ (.A(_20689_),
    .B1(_18697_),
    .B2(_20683_),
    .ZN(lce_data_cmd_o[301]));
 OAI21_X2 _48178_ (.A(_20688_),
    .B1(_20678_),
    .B2(\icache.lce.lce_cmd_inst.data_r [296]),
    .ZN(_20690_));
 AOI21_X4 _48179_ (.A(_20690_),
    .B1(_18705_),
    .B2(_20683_),
    .ZN(lce_data_cmd_o[302]));
 BUF_X4 _48180_ (.A(_20611_),
    .Z(_20691_));
 OAI21_X2 _48181_ (.A(_20688_),
    .B1(_20691_),
    .B2(\icache.lce.lce_cmd_inst.data_r [297]),
    .ZN(_20692_));
 AOI21_X4 _48182_ (.A(_20692_),
    .B1(_18715_),
    .B2(_20683_),
    .ZN(lce_data_cmd_o[303]));
 OAI21_X2 _48183_ (.A(_20688_),
    .B1(_20691_),
    .B2(\icache.lce.lce_cmd_inst.data_r [298]),
    .ZN(_20693_));
 AOI21_X4 _48184_ (.A(_20693_),
    .B1(_18723_),
    .B2(_20683_),
    .ZN(lce_data_cmd_o[304]));
 OAI21_X2 _48185_ (.A(_20688_),
    .B1(_20691_),
    .B2(\icache.lce.lce_cmd_inst.data_r [299]),
    .ZN(_20694_));
 AOI21_X4 _48186_ (.A(_20694_),
    .B1(_18731_),
    .B2(_20683_),
    .ZN(lce_data_cmd_o[305]));
 OAI21_X2 _48187_ (.A(_20688_),
    .B1(_20691_),
    .B2(\icache.lce.lce_cmd_inst.data_r [300]),
    .ZN(_20695_));
 BUF_X8 _48188_ (.A(_20630_),
    .Z(_20696_));
 AOI21_X4 _48189_ (.A(_20695_),
    .B1(_18740_),
    .B2(_20696_),
    .ZN(lce_data_cmd_o[306]));
 OAI21_X2 _48190_ (.A(_20688_),
    .B1(_20691_),
    .B2(\icache.lce.lce_cmd_inst.data_r [301]),
    .ZN(_20697_));
 AOI21_X4 _48191_ (.A(_20697_),
    .B1(_18750_),
    .B2(_20696_),
    .ZN(lce_data_cmd_o[307]));
 OAI21_X2 _48192_ (.A(_20688_),
    .B1(_20691_),
    .B2(\icache.lce.lce_cmd_inst.data_r [302]),
    .ZN(_20698_));
 AOI21_X4 _48193_ (.A(_20698_),
    .B1(_18758_),
    .B2(_20696_),
    .ZN(lce_data_cmd_o[308]));
 OAI21_X2 _48194_ (.A(_20688_),
    .B1(_20691_),
    .B2(\icache.lce.lce_cmd_inst.data_r [303]),
    .ZN(_20699_));
 AOI21_X4 _48195_ (.A(_20699_),
    .B1(_18767_),
    .B2(_20696_),
    .ZN(lce_data_cmd_o[309]));
 OAI21_X2 _48196_ (.A(_20688_),
    .B1(_20691_),
    .B2(\icache.lce.lce_cmd_inst.data_r [304]),
    .ZN(_20700_));
 AOI21_X4 _48197_ (.A(_20700_),
    .B1(_18777_),
    .B2(_20696_),
    .ZN(lce_data_cmd_o[310]));
 BUF_X8 _48198_ (.A(_20607_),
    .Z(_20701_));
 OAI21_X2 _48199_ (.A(_20701_),
    .B1(_20691_),
    .B2(\icache.lce.lce_cmd_inst.data_r [305]),
    .ZN(_20702_));
 AOI21_X4 _48200_ (.A(_20702_),
    .B1(_18785_),
    .B2(_20696_),
    .ZN(lce_data_cmd_o[311]));
 OAI21_X2 _48201_ (.A(_20701_),
    .B1(_20691_),
    .B2(\icache.lce.lce_cmd_inst.data_r [306]),
    .ZN(_20703_));
 AOI21_X4 _48202_ (.A(_20703_),
    .B1(_18793_),
    .B2(_20696_),
    .ZN(lce_data_cmd_o[312]));
 BUF_X16 _48203_ (.A(_20611_),
    .Z(_20704_));
 OAI21_X2 _48204_ (.A(_20701_),
    .B1(_20704_),
    .B2(\icache.lce.lce_cmd_inst.data_r [307]),
    .ZN(_20705_));
 AOI21_X4 _48205_ (.A(_20705_),
    .B1(_18802_),
    .B2(_20696_),
    .ZN(lce_data_cmd_o[313]));
 OAI21_X2 _48206_ (.A(_20701_),
    .B1(_20704_),
    .B2(\icache.lce.lce_cmd_inst.data_r [308]),
    .ZN(_20706_));
 AOI21_X4 _48207_ (.A(_20706_),
    .B1(_18812_),
    .B2(_20696_),
    .ZN(lce_data_cmd_o[314]));
 OAI21_X2 _48208_ (.A(_20701_),
    .B1(_20704_),
    .B2(\icache.lce.lce_cmd_inst.data_r [309]),
    .ZN(_20707_));
 AOI21_X4 _48209_ (.A(_20707_),
    .B1(_18821_),
    .B2(_20696_),
    .ZN(lce_data_cmd_o[315]));
 OAI21_X2 _48210_ (.A(_20701_),
    .B1(_20704_),
    .B2(\icache.lce.lce_cmd_inst.data_r [310]),
    .ZN(_20708_));
 BUF_X32 _48211_ (.A(_20630_),
    .Z(_20709_));
 AOI21_X4 _48212_ (.A(_20708_),
    .B1(_18829_),
    .B2(_20709_),
    .ZN(lce_data_cmd_o[316]));
 OAI21_X2 _48213_ (.A(_20701_),
    .B1(_20704_),
    .B2(\icache.lce.lce_cmd_inst.data_r [311]),
    .ZN(_20710_));
 AOI21_X4 _48214_ (.A(_20710_),
    .B1(_18837_),
    .B2(_20709_),
    .ZN(lce_data_cmd_o[317]));
 OAI21_X1 _48215_ (.A(_20701_),
    .B1(_20704_),
    .B2(\icache.lce.lce_cmd_inst.data_r [312]),
    .ZN(_20711_));
 AOI21_X4 _48216_ (.A(_20711_),
    .B1(_18845_),
    .B2(_20709_),
    .ZN(lce_data_cmd_o[318]));
 OAI21_X2 _48217_ (.A(_20701_),
    .B1(_20704_),
    .B2(\icache.lce.lce_cmd_inst.data_r [313]),
    .ZN(_20712_));
 AOI21_X4 _48218_ (.A(_20712_),
    .B1(_18853_),
    .B2(_20709_),
    .ZN(lce_data_cmd_o[319]));
 OAI21_X2 _48219_ (.A(_20701_),
    .B1(_20704_),
    .B2(\icache.lce.lce_cmd_inst.data_r [314]),
    .ZN(_20713_));
 AOI21_X4 _48220_ (.A(_20713_),
    .B1(_17955_),
    .B2(_20709_),
    .ZN(lce_data_cmd_o[320]));
 BUF_X8 _48221_ (.A(_20607_),
    .Z(_20714_));
 OAI21_X2 _48222_ (.A(_20714_),
    .B1(_20704_),
    .B2(\icache.lce.lce_cmd_inst.data_r [315]),
    .ZN(_20715_));
 AOI21_X4 _48223_ (.A(_20715_),
    .B1(_17966_),
    .B2(_20709_),
    .ZN(lce_data_cmd_o[321]));
 OAI21_X2 _48224_ (.A(_20714_),
    .B1(_20704_),
    .B2(\icache.lce.lce_cmd_inst.data_r [316]),
    .ZN(_20716_));
 AOI21_X4 _48225_ (.A(_20716_),
    .B1(_17975_),
    .B2(_20709_),
    .ZN(lce_data_cmd_o[322]));
 BUF_X4 _48226_ (.A(_20611_),
    .Z(_20717_));
 OAI21_X2 _48227_ (.A(_20714_),
    .B1(_20717_),
    .B2(\icache.lce.lce_cmd_inst.data_r [317]),
    .ZN(_20718_));
 AOI21_X4 _48228_ (.A(_20718_),
    .B1(_17985_),
    .B2(_20709_),
    .ZN(lce_data_cmd_o[323]));
 OAI21_X1 _48229_ (.A(_20714_),
    .B1(_20717_),
    .B2(\icache.lce.lce_cmd_inst.data_r [318]),
    .ZN(_20719_));
 AOI21_X4 _48230_ (.A(_20719_),
    .B1(_17995_),
    .B2(_20709_),
    .ZN(lce_data_cmd_o[324]));
 OAI21_X2 _48231_ (.A(_20714_),
    .B1(_20717_),
    .B2(\icache.lce.lce_cmd_inst.data_r [319]),
    .ZN(_20720_));
 AOI21_X4 _48232_ (.A(_20720_),
    .B1(_18003_),
    .B2(_20709_),
    .ZN(lce_data_cmd_o[325]));
 OAI21_X2 _48233_ (.A(_20714_),
    .B1(_20717_),
    .B2(\icache.lce.lce_cmd_inst.data_r [320]),
    .ZN(_20721_));
 BUF_X8 _48234_ (.A(_20630_),
    .Z(_20722_));
 AOI21_X4 _48235_ (.A(_20721_),
    .B1(_18013_),
    .B2(_20722_),
    .ZN(lce_data_cmd_o[326]));
 OAI21_X2 _48236_ (.A(_20714_),
    .B1(_20717_),
    .B2(\icache.lce.lce_cmd_inst.data_r [321]),
    .ZN(_20723_));
 AOI21_X4 _48237_ (.A(_20723_),
    .B1(_18023_),
    .B2(_20722_),
    .ZN(lce_data_cmd_o[327]));
 OAI21_X2 _48238_ (.A(_20714_),
    .B1(_20717_),
    .B2(\icache.lce.lce_cmd_inst.data_r [322]),
    .ZN(_20724_));
 AOI21_X4 _48239_ (.A(_20724_),
    .B1(_18032_),
    .B2(_20722_),
    .ZN(lce_data_cmd_o[328]));
 OAI21_X2 _48240_ (.A(_20714_),
    .B1(_20717_),
    .B2(\icache.lce.lce_cmd_inst.data_r [323]),
    .ZN(_20725_));
 AOI21_X4 _48241_ (.A(_20725_),
    .B1(_18041_),
    .B2(_20722_),
    .ZN(lce_data_cmd_o[329]));
 OAI21_X2 _48242_ (.A(_20714_),
    .B1(_20717_),
    .B2(\icache.lce.lce_cmd_inst.data_r [324]),
    .ZN(_20726_));
 AOI21_X4 _48243_ (.A(_20726_),
    .B1(_18049_),
    .B2(_20722_),
    .ZN(lce_data_cmd_o[330]));
 BUF_X8 _48244_ (.A(_20607_),
    .Z(_20727_));
 OAI21_X1 _48245_ (.A(_20727_),
    .B1(_20717_),
    .B2(\icache.lce.lce_cmd_inst.data_r [325]),
    .ZN(_20728_));
 AOI21_X4 _48246_ (.A(_20728_),
    .B1(_18057_),
    .B2(_20722_),
    .ZN(lce_data_cmd_o[331]));
 OAI21_X2 _48247_ (.A(_20727_),
    .B1(_20717_),
    .B2(\icache.lce.lce_cmd_inst.data_r [326]),
    .ZN(_20729_));
 AOI21_X4 _48248_ (.A(_20729_),
    .B1(_18065_),
    .B2(_20722_),
    .ZN(lce_data_cmd_o[332]));
 BUF_X8 _48249_ (.A(_20611_),
    .Z(_20730_));
 OAI21_X2 _48250_ (.A(_20727_),
    .B1(_20730_),
    .B2(\icache.lce.lce_cmd_inst.data_r [327]),
    .ZN(_20731_));
 AOI21_X4 _48251_ (.A(_20731_),
    .B1(_18073_),
    .B2(_20722_),
    .ZN(lce_data_cmd_o[333]));
 OAI21_X2 _48252_ (.A(_20727_),
    .B1(_20730_),
    .B2(\icache.lce.lce_cmd_inst.data_r [328]),
    .ZN(_20732_));
 AOI21_X4 _48253_ (.A(_20732_),
    .B1(_18081_),
    .B2(_20722_),
    .ZN(lce_data_cmd_o[334]));
 OAI21_X2 _48254_ (.A(_20727_),
    .B1(_20730_),
    .B2(\icache.lce.lce_cmd_inst.data_r [329]),
    .ZN(_20733_));
 AOI21_X4 _48255_ (.A(_20733_),
    .B1(_18090_),
    .B2(_20722_),
    .ZN(lce_data_cmd_o[335]));
 OAI21_X2 _48256_ (.A(_20727_),
    .B1(_20730_),
    .B2(\icache.lce.lce_cmd_inst.data_r [330]),
    .ZN(_20734_));
 BUF_X16 _48257_ (.A(_20630_),
    .Z(_20735_));
 AOI21_X4 _48258_ (.A(_20734_),
    .B1(_18100_),
    .B2(_20735_),
    .ZN(lce_data_cmd_o[336]));
 OAI21_X2 _48259_ (.A(_20727_),
    .B1(_20730_),
    .B2(\icache.lce.lce_cmd_inst.data_r [331]),
    .ZN(_20736_));
 AOI21_X4 _48260_ (.A(_20736_),
    .B1(_18109_),
    .B2(_20735_),
    .ZN(lce_data_cmd_o[337]));
 OAI21_X2 _48261_ (.A(_20727_),
    .B1(_20730_),
    .B2(\icache.lce.lce_cmd_inst.data_r [332]),
    .ZN(_20737_));
 AOI21_X4 _48262_ (.A(_20737_),
    .B1(_18119_),
    .B2(_20735_),
    .ZN(lce_data_cmd_o[338]));
 OAI21_X2 _48263_ (.A(_20727_),
    .B1(_20730_),
    .B2(\icache.lce.lce_cmd_inst.data_r [333]),
    .ZN(_20738_));
 AOI21_X4 _48264_ (.A(_20738_),
    .B1(_18128_),
    .B2(_20735_),
    .ZN(lce_data_cmd_o[339]));
 OAI21_X2 _48265_ (.A(_20727_),
    .B1(_20730_),
    .B2(\icache.lce.lce_cmd_inst.data_r [334]),
    .ZN(_20739_));
 AOI21_X4 _48266_ (.A(_20739_),
    .B1(_18137_),
    .B2(_20735_),
    .ZN(lce_data_cmd_o[340]));
 BUF_X32 _48267_ (.A(_07607_),
    .Z(_20740_));
 BUF_X8 _48268_ (.A(_20740_),
    .Z(_20741_));
 OAI21_X2 _48269_ (.A(_20741_),
    .B1(_20730_),
    .B2(\icache.lce.lce_cmd_inst.data_r [335]),
    .ZN(_20742_));
 AOI21_X4 _48270_ (.A(_20742_),
    .B1(_18145_),
    .B2(_20735_),
    .ZN(lce_data_cmd_o[341]));
 OAI21_X2 _48271_ (.A(_20741_),
    .B1(_20730_),
    .B2(\icache.lce.lce_cmd_inst.data_r [336]),
    .ZN(_20743_));
 AOI21_X4 _48272_ (.A(_20743_),
    .B1(_18153_),
    .B2(_20735_),
    .ZN(lce_data_cmd_o[342]));
 BUF_X32 _48273_ (.A(_15295_),
    .Z(_20744_));
 BUF_X8 _48274_ (.A(_20744_),
    .Z(_20745_));
 OAI21_X2 _48275_ (.A(_20741_),
    .B1(_20745_),
    .B2(\icache.lce.lce_cmd_inst.data_r [337]),
    .ZN(_20746_));
 AOI21_X4 _48276_ (.A(_20746_),
    .B1(_18161_),
    .B2(_20735_),
    .ZN(lce_data_cmd_o[343]));
 OAI21_X2 _48277_ (.A(_20741_),
    .B1(_20745_),
    .B2(\icache.lce.lce_cmd_inst.data_r [338]),
    .ZN(_20747_));
 AOI21_X4 _48278_ (.A(_20747_),
    .B1(_18170_),
    .B2(_20735_),
    .ZN(lce_data_cmd_o[344]));
 OAI21_X2 _48279_ (.A(_20741_),
    .B1(_20745_),
    .B2(\icache.lce.lce_cmd_inst.data_r [339]),
    .ZN(_20748_));
 AOI21_X4 _48280_ (.A(_20748_),
    .B1(_18178_),
    .B2(_20735_),
    .ZN(lce_data_cmd_o[345]));
 OAI21_X2 _48281_ (.A(_20741_),
    .B1(_20745_),
    .B2(\icache.lce.lce_cmd_inst.data_r [340]),
    .ZN(_20749_));
 BUF_X16 _48282_ (.A(_20630_),
    .Z(_20750_));
 AOI21_X4 _48283_ (.A(_20749_),
    .B1(_18188_),
    .B2(_20750_),
    .ZN(lce_data_cmd_o[346]));
 OAI21_X2 _48284_ (.A(_20741_),
    .B1(_20745_),
    .B2(\icache.lce.lce_cmd_inst.data_r [341]),
    .ZN(_20751_));
 AOI21_X4 _48285_ (.A(_20751_),
    .B1(_18197_),
    .B2(_20750_),
    .ZN(lce_data_cmd_o[347]));
 OAI21_X2 _48286_ (.A(_20741_),
    .B1(_20745_),
    .B2(\icache.lce.lce_cmd_inst.data_r [342]),
    .ZN(_20752_));
 AOI21_X4 _48287_ (.A(_20752_),
    .B1(_18205_),
    .B2(_20750_),
    .ZN(lce_data_cmd_o[348]));
 OAI21_X2 _48288_ (.A(_20741_),
    .B1(_20745_),
    .B2(\icache.lce.lce_cmd_inst.data_r [343]),
    .ZN(_20753_));
 AOI21_X4 _48289_ (.A(_20753_),
    .B1(_18216_),
    .B2(_20750_),
    .ZN(lce_data_cmd_o[349]));
 OAI21_X2 _48290_ (.A(_20741_),
    .B1(_20745_),
    .B2(\icache.lce.lce_cmd_inst.data_r [344]),
    .ZN(_20754_));
 AOI21_X4 _48291_ (.A(_20754_),
    .B1(_18224_),
    .B2(_20750_),
    .ZN(lce_data_cmd_o[350]));
 BUF_X8 _48292_ (.A(_20740_),
    .Z(_20755_));
 OAI21_X2 _48293_ (.A(_20755_),
    .B1(_20745_),
    .B2(\icache.lce.lce_cmd_inst.data_r [345]),
    .ZN(_20756_));
 AOI21_X4 _48294_ (.A(_20756_),
    .B1(_18233_),
    .B2(_20750_),
    .ZN(lce_data_cmd_o[351]));
 OAI21_X2 _48295_ (.A(_20755_),
    .B1(_20745_),
    .B2(\icache.lce.lce_cmd_inst.data_r [346]),
    .ZN(_20757_));
 AOI21_X4 _48296_ (.A(_20757_),
    .B1(_18243_),
    .B2(_20750_),
    .ZN(lce_data_cmd_o[352]));
 BUF_X8 _48297_ (.A(_20744_),
    .Z(_20758_));
 OAI21_X2 _48298_ (.A(_20755_),
    .B1(_20758_),
    .B2(\icache.lce.lce_cmd_inst.data_r [347]),
    .ZN(_20759_));
 AOI21_X4 _48299_ (.A(_20759_),
    .B1(_18251_),
    .B2(_20750_),
    .ZN(lce_data_cmd_o[353]));
 OAI21_X2 _48300_ (.A(_20755_),
    .B1(_20758_),
    .B2(\icache.lce.lce_cmd_inst.data_r [348]),
    .ZN(_20760_));
 AOI21_X4 _48301_ (.A(_20760_),
    .B1(_18259_),
    .B2(_20750_),
    .ZN(lce_data_cmd_o[354]));
 OAI21_X2 _48302_ (.A(_20755_),
    .B1(_20758_),
    .B2(\icache.lce.lce_cmd_inst.data_r [349]),
    .ZN(_20761_));
 AOI21_X4 _48303_ (.A(_20761_),
    .B1(_18267_),
    .B2(_20750_),
    .ZN(lce_data_cmd_o[355]));
 OAI21_X2 _48304_ (.A(_20755_),
    .B1(_20758_),
    .B2(\icache.lce.lce_cmd_inst.data_r [350]),
    .ZN(_20762_));
 BUF_X32 _48305_ (.A(_15295_),
    .Z(_20763_));
 BUF_X16 _48306_ (.A(_20763_),
    .Z(_20764_));
 AOI21_X4 _48307_ (.A(_20762_),
    .B1(_18277_),
    .B2(_20764_),
    .ZN(lce_data_cmd_o[356]));
 OAI21_X1 _48308_ (.A(_20755_),
    .B1(_20758_),
    .B2(\icache.lce.lce_cmd_inst.data_r [351]),
    .ZN(_20765_));
 AOI21_X4 _48309_ (.A(_20765_),
    .B1(_18285_),
    .B2(_20764_),
    .ZN(lce_data_cmd_o[357]));
 OAI21_X2 _48310_ (.A(_20755_),
    .B1(_20758_),
    .B2(\icache.lce.lce_cmd_inst.data_r [352]),
    .ZN(_20766_));
 AOI21_X4 _48311_ (.A(_20766_),
    .B1(_18293_),
    .B2(_20764_),
    .ZN(lce_data_cmd_o[358]));
 OAI21_X2 _48312_ (.A(_20755_),
    .B1(_20758_),
    .B2(\icache.lce.lce_cmd_inst.data_r [353]),
    .ZN(_20767_));
 AOI21_X4 _48313_ (.A(_20767_),
    .B1(_18304_),
    .B2(_20764_),
    .ZN(lce_data_cmd_o[359]));
 OAI21_X2 _48314_ (.A(_20755_),
    .B1(_20758_),
    .B2(\icache.lce.lce_cmd_inst.data_r [354]),
    .ZN(_20768_));
 AOI21_X4 _48315_ (.A(_20768_),
    .B1(_18314_),
    .B2(_20764_),
    .ZN(lce_data_cmd_o[360]));
 BUF_X16 _48316_ (.A(_20740_),
    .Z(_20769_));
 OAI21_X2 _48317_ (.A(_20769_),
    .B1(_20758_),
    .B2(\icache.lce.lce_cmd_inst.data_r [355]),
    .ZN(_20770_));
 AOI21_X4 _48318_ (.A(_20770_),
    .B1(_18322_),
    .B2(_20764_),
    .ZN(lce_data_cmd_o[361]));
 OAI21_X2 _48319_ (.A(_20769_),
    .B1(_20758_),
    .B2(\icache.lce.lce_cmd_inst.data_r [356]),
    .ZN(_20771_));
 AOI21_X4 _48320_ (.A(_20771_),
    .B1(_18332_),
    .B2(_20764_),
    .ZN(lce_data_cmd_o[362]));
 BUF_X8 _48321_ (.A(_20744_),
    .Z(_20772_));
 OAI21_X2 _48322_ (.A(_20769_),
    .B1(_20772_),
    .B2(\icache.lce.lce_cmd_inst.data_r [357]),
    .ZN(_20773_));
 AOI21_X4 _48323_ (.A(_20773_),
    .B1(_18341_),
    .B2(_20764_),
    .ZN(lce_data_cmd_o[363]));
 OAI21_X2 _48324_ (.A(_20769_),
    .B1(_20772_),
    .B2(\icache.lce.lce_cmd_inst.data_r [358]),
    .ZN(_20774_));
 AOI21_X4 _48325_ (.A(_20774_),
    .B1(_18349_),
    .B2(_20764_),
    .ZN(lce_data_cmd_o[364]));
 OAI21_X2 _48326_ (.A(_20769_),
    .B1(_20772_),
    .B2(\icache.lce.lce_cmd_inst.data_r [359]),
    .ZN(_20775_));
 AOI21_X4 _48327_ (.A(_20775_),
    .B1(_18359_),
    .B2(_20764_),
    .ZN(lce_data_cmd_o[365]));
 OAI21_X1 _48328_ (.A(_20769_),
    .B1(_20772_),
    .B2(\icache.lce.lce_cmd_inst.data_r [360]),
    .ZN(_20776_));
 BUF_X8 _48329_ (.A(_20763_),
    .Z(_20777_));
 AOI21_X4 _48330_ (.A(_20776_),
    .B1(_18370_),
    .B2(_20777_),
    .ZN(lce_data_cmd_o[366]));
 OAI21_X2 _48331_ (.A(_20769_),
    .B1(_20772_),
    .B2(\icache.lce.lce_cmd_inst.data_r [361]),
    .ZN(_20778_));
 AOI21_X4 _48332_ (.A(_20778_),
    .B1(_18380_),
    .B2(_20777_),
    .ZN(lce_data_cmd_o[367]));
 OAI21_X2 _48333_ (.A(_20769_),
    .B1(_20772_),
    .B2(\icache.lce.lce_cmd_inst.data_r [362]),
    .ZN(_20779_));
 AOI21_X4 _48334_ (.A(_20779_),
    .B1(_18389_),
    .B2(_20777_),
    .ZN(lce_data_cmd_o[368]));
 OAI21_X2 _48335_ (.A(_20769_),
    .B1(_20772_),
    .B2(\icache.lce.lce_cmd_inst.data_r [363]),
    .ZN(_20780_));
 AOI21_X4 _48336_ (.A(_20780_),
    .B1(_18398_),
    .B2(_20777_),
    .ZN(lce_data_cmd_o[369]));
 OAI21_X2 _48337_ (.A(_20769_),
    .B1(_20772_),
    .B2(\icache.lce.lce_cmd_inst.data_r [364]),
    .ZN(_20781_));
 AOI21_X4 _48338_ (.A(_20781_),
    .B1(_18406_),
    .B2(_20777_),
    .ZN(lce_data_cmd_o[370]));
 BUF_X8 _48339_ (.A(_20740_),
    .Z(_20782_));
 OAI21_X2 _48340_ (.A(_20782_),
    .B1(_20772_),
    .B2(\icache.lce.lce_cmd_inst.data_r [365]),
    .ZN(_20783_));
 AOI21_X4 _48341_ (.A(_20783_),
    .B1(_18414_),
    .B2(_20777_),
    .ZN(lce_data_cmd_o[371]));
 OAI21_X2 _48342_ (.A(_20782_),
    .B1(_20772_),
    .B2(\icache.lce.lce_cmd_inst.data_r [366]),
    .ZN(_20784_));
 AOI21_X4 _48343_ (.A(_20784_),
    .B1(_18423_),
    .B2(_20777_),
    .ZN(lce_data_cmd_o[372]));
 BUF_X8 _48344_ (.A(_20744_),
    .Z(_20785_));
 OAI21_X2 _48345_ (.A(_20782_),
    .B1(_20785_),
    .B2(\icache.lce.lce_cmd_inst.data_r [367]),
    .ZN(_20786_));
 AOI21_X4 _48346_ (.A(_20786_),
    .B1(_18433_),
    .B2(_20777_),
    .ZN(lce_data_cmd_o[373]));
 OAI21_X2 _48347_ (.A(_20782_),
    .B1(_20785_),
    .B2(\icache.lce.lce_cmd_inst.data_r [368]),
    .ZN(_20787_));
 AOI21_X4 _48348_ (.A(_20787_),
    .B1(_18442_),
    .B2(_20777_),
    .ZN(lce_data_cmd_o[374]));
 OAI21_X2 _48349_ (.A(_20782_),
    .B1(_20785_),
    .B2(\icache.lce.lce_cmd_inst.data_r [369]),
    .ZN(_20788_));
 AOI21_X4 _48350_ (.A(_20788_),
    .B1(_18450_),
    .B2(_20777_),
    .ZN(lce_data_cmd_o[375]));
 OAI21_X2 _48351_ (.A(_20782_),
    .B1(_20785_),
    .B2(\icache.lce.lce_cmd_inst.data_r [370]),
    .ZN(_20789_));
 BUF_X8 _48352_ (.A(_20763_),
    .Z(_20790_));
 AOI21_X4 _48353_ (.A(_20789_),
    .B1(_18462_),
    .B2(_20790_),
    .ZN(lce_data_cmd_o[376]));
 OAI21_X2 _48354_ (.A(_20782_),
    .B1(_20785_),
    .B2(\icache.lce.lce_cmd_inst.data_r [371]),
    .ZN(_20791_));
 AOI21_X4 _48355_ (.A(_20791_),
    .B1(_18472_),
    .B2(_20790_),
    .ZN(lce_data_cmd_o[377]));
 OAI21_X2 _48356_ (.A(_20782_),
    .B1(_20785_),
    .B2(\icache.lce.lce_cmd_inst.data_r [372]),
    .ZN(_20792_));
 AOI21_X4 _48357_ (.A(_20792_),
    .B1(_18482_),
    .B2(_20790_),
    .ZN(lce_data_cmd_o[378]));
 OAI21_X2 _48358_ (.A(_20782_),
    .B1(_20785_),
    .B2(\icache.lce.lce_cmd_inst.data_r [373]),
    .ZN(_20793_));
 AOI21_X4 _48359_ (.A(_20793_),
    .B1(_18491_),
    .B2(_20790_),
    .ZN(lce_data_cmd_o[379]));
 OAI21_X2 _48360_ (.A(_20782_),
    .B1(_20785_),
    .B2(\icache.lce.lce_cmd_inst.data_r [374]),
    .ZN(_20794_));
 AOI21_X4 _48361_ (.A(_20794_),
    .B1(_18499_),
    .B2(_20790_),
    .ZN(lce_data_cmd_o[380]));
 BUF_X8 _48362_ (.A(_20740_),
    .Z(_20795_));
 OAI21_X2 _48363_ (.A(_20795_),
    .B1(_20785_),
    .B2(\icache.lce.lce_cmd_inst.data_r [375]),
    .ZN(_20796_));
 AOI21_X4 _48364_ (.A(_20796_),
    .B1(_18508_),
    .B2(_20790_),
    .ZN(lce_data_cmd_o[381]));
 OAI21_X2 _48365_ (.A(_20795_),
    .B1(_20785_),
    .B2(\icache.lce.lce_cmd_inst.data_r [376]),
    .ZN(_20797_));
 AOI21_X4 _48366_ (.A(_20797_),
    .B1(_18518_),
    .B2(_20790_),
    .ZN(lce_data_cmd_o[382]));
 BUF_X8 _48367_ (.A(_20744_),
    .Z(_20798_));
 OAI21_X2 _48368_ (.A(_20795_),
    .B1(_20798_),
    .B2(\icache.lce.lce_cmd_inst.data_r [377]),
    .ZN(_20799_));
 AOI21_X4 _48369_ (.A(_20799_),
    .B1(_18526_),
    .B2(_20790_),
    .ZN(lce_data_cmd_o[383]));
 OAI21_X2 _48370_ (.A(_20795_),
    .B1(_20798_),
    .B2(\icache.lce.lce_cmd_inst.data_r [378]),
    .ZN(_20800_));
 AOI21_X4 _48371_ (.A(_20800_),
    .B1(_18535_),
    .B2(_20790_),
    .ZN(lce_data_cmd_o[384]));
 OAI21_X2 _48372_ (.A(_20795_),
    .B1(_20798_),
    .B2(\icache.lce.lce_cmd_inst.data_r [379]),
    .ZN(_20801_));
 AOI21_X4 _48373_ (.A(_20801_),
    .B1(_18543_),
    .B2(_20790_),
    .ZN(lce_data_cmd_o[385]));
 OAI21_X2 _48374_ (.A(_20795_),
    .B1(_20798_),
    .B2(\icache.lce.lce_cmd_inst.data_r [380]),
    .ZN(_20802_));
 BUF_X8 _48375_ (.A(_20763_),
    .Z(_20803_));
 AOI21_X4 _48376_ (.A(_20802_),
    .B1(_18553_),
    .B2(_20803_),
    .ZN(lce_data_cmd_o[386]));
 OAI21_X1 _48377_ (.A(_20795_),
    .B1(_20798_),
    .B2(\icache.lce.lce_cmd_inst.data_r [381]),
    .ZN(_20804_));
 AOI21_X4 _48378_ (.A(_20804_),
    .B1(_18561_),
    .B2(_20803_),
    .ZN(lce_data_cmd_o[387]));
 OAI21_X1 _48379_ (.A(_20795_),
    .B1(_20798_),
    .B2(\icache.lce.lce_cmd_inst.data_r [382]),
    .ZN(_20805_));
 AOI21_X4 _48380_ (.A(_20805_),
    .B1(_18571_),
    .B2(_20803_),
    .ZN(lce_data_cmd_o[388]));
 OAI21_X2 _48381_ (.A(_20795_),
    .B1(_20798_),
    .B2(\icache.lce.lce_cmd_inst.data_r [383]),
    .ZN(_20806_));
 AOI21_X4 _48382_ (.A(_20806_),
    .B1(_18580_),
    .B2(_20803_),
    .ZN(lce_data_cmd_o[389]));
 OAI21_X1 _48383_ (.A(_20795_),
    .B1(_20798_),
    .B2(\icache.lce.lce_cmd_inst.data_r [384]),
    .ZN(_20807_));
 AOI21_X4 _48384_ (.A(_20807_),
    .B1(_18589_),
    .B2(_20803_),
    .ZN(lce_data_cmd_o[390]));
 BUF_X16 _48385_ (.A(_20740_),
    .Z(_20808_));
 OAI21_X2 _48386_ (.A(_20808_),
    .B1(_20798_),
    .B2(\icache.lce.lce_cmd_inst.data_r [385]),
    .ZN(_20809_));
 AOI21_X4 _48387_ (.A(_20809_),
    .B1(_18607_),
    .B2(_20803_),
    .ZN(lce_data_cmd_o[391]));
 OAI21_X2 _48388_ (.A(_20808_),
    .B1(_20798_),
    .B2(\icache.lce.lce_cmd_inst.data_r [386]),
    .ZN(_20810_));
 AOI21_X4 _48389_ (.A(_20810_),
    .B1(_18623_),
    .B2(_20803_),
    .ZN(lce_data_cmd_o[392]));
 BUF_X16 _48390_ (.A(_20744_),
    .Z(_20811_));
 OAI21_X2 _48391_ (.A(_20808_),
    .B1(_20811_),
    .B2(\icache.lce.lce_cmd_inst.data_r [387]),
    .ZN(_20812_));
 AOI21_X4 _48392_ (.A(_20812_),
    .B1(_18638_),
    .B2(_20803_),
    .ZN(lce_data_cmd_o[393]));
 OAI21_X2 _48393_ (.A(_20808_),
    .B1(_20811_),
    .B2(\icache.lce.lce_cmd_inst.data_r [388]),
    .ZN(_20813_));
 AOI21_X4 _48394_ (.A(_20813_),
    .B1(_18653_),
    .B2(_20803_),
    .ZN(lce_data_cmd_o[394]));
 OAI21_X1 _48395_ (.A(_20808_),
    .B1(_20811_),
    .B2(\icache.lce.lce_cmd_inst.data_r [389]),
    .ZN(_20814_));
 AOI21_X4 _48396_ (.A(_20814_),
    .B1(_18671_),
    .B2(_20803_),
    .ZN(lce_data_cmd_o[395]));
 OAI21_X2 _48397_ (.A(_20808_),
    .B1(_20811_),
    .B2(\icache.lce.lce_cmd_inst.data_r [390]),
    .ZN(_20815_));
 BUF_X8 _48398_ (.A(_20763_),
    .Z(_20816_));
 AOI21_X4 _48399_ (.A(_20815_),
    .B1(_18689_),
    .B2(_20816_),
    .ZN(lce_data_cmd_o[396]));
 OAI21_X2 _48400_ (.A(_20808_),
    .B1(_20811_),
    .B2(\icache.lce.lce_cmd_inst.data_r [391]),
    .ZN(_20817_));
 AOI21_X4 _48401_ (.A(_20817_),
    .B1(_17913_),
    .B2(_20816_),
    .ZN(lce_data_cmd_o[397]));
 OAI21_X2 _48402_ (.A(_20808_),
    .B1(_20811_),
    .B2(\icache.lce.lce_cmd_inst.data_r [392]),
    .ZN(_20818_));
 AOI21_X4 _48403_ (.A(_20818_),
    .B1(_17930_),
    .B2(_20816_),
    .ZN(lce_data_cmd_o[398]));
 OAI21_X2 _48404_ (.A(_20808_),
    .B1(_20811_),
    .B2(\icache.lce.lce_cmd_inst.data_r [393]),
    .ZN(_20819_));
 AOI21_X4 _48405_ (.A(_20819_),
    .B1(_17947_),
    .B2(_20816_),
    .ZN(lce_data_cmd_o[399]));
 OAI21_X2 _48406_ (.A(_20808_),
    .B1(_20811_),
    .B2(\icache.lce.lce_cmd_inst.data_r [394]),
    .ZN(_20820_));
 AOI21_X4 _48407_ (.A(_20820_),
    .B1(_17579_),
    .B2(_20816_),
    .ZN(lce_data_cmd_o[400]));
 BUF_X8 _48408_ (.A(_20740_),
    .Z(_20821_));
 OAI21_X2 _48409_ (.A(_20821_),
    .B1(_20811_),
    .B2(\icache.lce.lce_cmd_inst.data_r [395]),
    .ZN(_20822_));
 AOI21_X4 _48410_ (.A(_20822_),
    .B1(_17598_),
    .B2(_20816_),
    .ZN(lce_data_cmd_o[401]));
 OAI21_X2 _48411_ (.A(_20821_),
    .B1(_20811_),
    .B2(\icache.lce.lce_cmd_inst.data_r [396]),
    .ZN(_20823_));
 AOI21_X4 _48412_ (.A(_20823_),
    .B1(_17614_),
    .B2(_20816_),
    .ZN(lce_data_cmd_o[402]));
 BUF_X4 _48413_ (.A(_20744_),
    .Z(_20824_));
 OAI21_X2 _48414_ (.A(_20821_),
    .B1(_20824_),
    .B2(\icache.lce.lce_cmd_inst.data_r [397]),
    .ZN(_20825_));
 AOI21_X4 _48415_ (.A(_20825_),
    .B1(_17636_),
    .B2(_20816_),
    .ZN(lce_data_cmd_o[403]));
 OAI21_X2 _48416_ (.A(_20821_),
    .B1(_20824_),
    .B2(\icache.lce.lce_cmd_inst.data_r [398]),
    .ZN(_20826_));
 AOI21_X4 _48417_ (.A(_20826_),
    .B1(_17652_),
    .B2(_20816_),
    .ZN(lce_data_cmd_o[404]));
 OAI21_X2 _48418_ (.A(_20821_),
    .B1(_20824_),
    .B2(\icache.lce.lce_cmd_inst.data_r [399]),
    .ZN(_20827_));
 AOI21_X4 _48419_ (.A(_20827_),
    .B1(_17668_),
    .B2(_20816_),
    .ZN(lce_data_cmd_o[405]));
 OAI21_X1 _48420_ (.A(_20821_),
    .B1(_20824_),
    .B2(\icache.lce.lce_cmd_inst.data_r [400]),
    .ZN(_20828_));
 BUF_X8 _48421_ (.A(_20763_),
    .Z(_20829_));
 AOI21_X4 _48422_ (.A(_20828_),
    .B1(_17686_),
    .B2(_20829_),
    .ZN(lce_data_cmd_o[406]));
 OAI21_X1 _48423_ (.A(_20821_),
    .B1(_20824_),
    .B2(\icache.lce.lce_cmd_inst.data_r [401]),
    .ZN(_20830_));
 AOI21_X4 _48424_ (.A(_20830_),
    .B1(_17704_),
    .B2(_20829_),
    .ZN(lce_data_cmd_o[407]));
 OAI21_X1 _48425_ (.A(_20821_),
    .B1(_20824_),
    .B2(\icache.lce.lce_cmd_inst.data_r [402]),
    .ZN(_20831_));
 AOI21_X4 _48426_ (.A(_20831_),
    .B1(_17722_),
    .B2(_20829_),
    .ZN(lce_data_cmd_o[408]));
 OAI21_X2 _48427_ (.A(_20821_),
    .B1(_20824_),
    .B2(\icache.lce.lce_cmd_inst.data_r [403]),
    .ZN(_20832_));
 AOI21_X4 _48428_ (.A(_20832_),
    .B1(_17740_),
    .B2(_20829_),
    .ZN(lce_data_cmd_o[409]));
 OAI21_X2 _48429_ (.A(_20821_),
    .B1(_20824_),
    .B2(\icache.lce.lce_cmd_inst.data_r [404]),
    .ZN(_20833_));
 AOI21_X4 _48430_ (.A(_20833_),
    .B1(_17756_),
    .B2(_20829_),
    .ZN(lce_data_cmd_o[410]));
 BUF_X8 _48431_ (.A(_20740_),
    .Z(_20834_));
 OAI21_X2 _48432_ (.A(_20834_),
    .B1(_20824_),
    .B2(\icache.lce.lce_cmd_inst.data_r [405]),
    .ZN(_20835_));
 AOI21_X4 _48433_ (.A(_20835_),
    .B1(_17771_),
    .B2(_20829_),
    .ZN(lce_data_cmd_o[411]));
 OAI21_X2 _48434_ (.A(_20834_),
    .B1(_20824_),
    .B2(\icache.lce.lce_cmd_inst.data_r [406]),
    .ZN(_20836_));
 AOI21_X4 _48435_ (.A(_20836_),
    .B1(_17791_),
    .B2(_20829_),
    .ZN(lce_data_cmd_o[412]));
 BUF_X8 _48436_ (.A(_20744_),
    .Z(_20837_));
 OAI21_X2 _48437_ (.A(_20834_),
    .B1(_20837_),
    .B2(\icache.lce.lce_cmd_inst.data_r [407]),
    .ZN(_20838_));
 AOI21_X4 _48438_ (.A(_20838_),
    .B1(_17808_),
    .B2(_20829_),
    .ZN(lce_data_cmd_o[413]));
 OAI21_X2 _48439_ (.A(_20834_),
    .B1(_20837_),
    .B2(\icache.lce.lce_cmd_inst.data_r [408]),
    .ZN(_20839_));
 AOI21_X4 _48440_ (.A(_20839_),
    .B1(_17825_),
    .B2(_20829_),
    .ZN(lce_data_cmd_o[414]));
 OAI21_X2 _48441_ (.A(_20834_),
    .B1(_20837_),
    .B2(\icache.lce.lce_cmd_inst.data_r [409]),
    .ZN(_20840_));
 AOI21_X4 _48442_ (.A(_20840_),
    .B1(_17843_),
    .B2(_20829_),
    .ZN(lce_data_cmd_o[415]));
 OAI21_X2 _48443_ (.A(_20834_),
    .B1(_20837_),
    .B2(\icache.lce.lce_cmd_inst.data_r [410]),
    .ZN(_20841_));
 BUF_X8 _48444_ (.A(_20763_),
    .Z(_20842_));
 AOI21_X4 _48445_ (.A(_20841_),
    .B1(_17860_),
    .B2(_20842_),
    .ZN(lce_data_cmd_o[416]));
 OAI21_X2 _48446_ (.A(_20834_),
    .B1(_20837_),
    .B2(\icache.lce.lce_cmd_inst.data_r [411]),
    .ZN(_20843_));
 AOI21_X4 _48447_ (.A(_20843_),
    .B1(_17876_),
    .B2(_20842_),
    .ZN(lce_data_cmd_o[417]));
 OAI21_X2 _48448_ (.A(_20834_),
    .B1(_20837_),
    .B2(\icache.lce.lce_cmd_inst.data_r [412]),
    .ZN(_20844_));
 AOI21_X4 _48449_ (.A(_20844_),
    .B1(_17896_),
    .B2(_20842_),
    .ZN(lce_data_cmd_o[418]));
 OAI21_X2 _48450_ (.A(_20834_),
    .B1(_20837_),
    .B2(\icache.lce.lce_cmd_inst.data_r [413]),
    .ZN(_20845_));
 AOI21_X4 _48451_ (.A(_20845_),
    .B1(_15926_),
    .B2(_20842_),
    .ZN(lce_data_cmd_o[419]));
 OAI21_X2 _48452_ (.A(_20834_),
    .B1(_20837_),
    .B2(\icache.lce.lce_cmd_inst.data_r [414]),
    .ZN(_20846_));
 AOI21_X4 _48453_ (.A(_20846_),
    .B1(_15950_),
    .B2(_20842_),
    .ZN(lce_data_cmd_o[420]));
 BUF_X8 _48454_ (.A(_20740_),
    .Z(_20847_));
 OAI21_X2 _48455_ (.A(_20847_),
    .B1(_20837_),
    .B2(\icache.lce.lce_cmd_inst.data_r [415]),
    .ZN(_20848_));
 AOI21_X4 _48456_ (.A(_20848_),
    .B1(_15972_),
    .B2(_20842_),
    .ZN(lce_data_cmd_o[421]));
 OAI21_X2 _48457_ (.A(_20847_),
    .B1(_20837_),
    .B2(\icache.lce.lce_cmd_inst.data_r [416]),
    .ZN(_20849_));
 AOI21_X4 _48458_ (.A(_20849_),
    .B1(_15998_),
    .B2(_20842_),
    .ZN(lce_data_cmd_o[422]));
 BUF_X8 _48459_ (.A(_20744_),
    .Z(_20850_));
 OAI21_X2 _48460_ (.A(_20847_),
    .B1(_20850_),
    .B2(\icache.lce.lce_cmd_inst.data_r [417]),
    .ZN(_20851_));
 AOI21_X4 _48461_ (.A(_20851_),
    .B1(_16028_),
    .B2(_20842_),
    .ZN(lce_data_cmd_o[423]));
 OAI21_X2 _48462_ (.A(_20847_),
    .B1(_20850_),
    .B2(\icache.lce.lce_cmd_inst.data_r [418]),
    .ZN(_20852_));
 AOI21_X4 _48463_ (.A(_20852_),
    .B1(_16047_),
    .B2(_20842_),
    .ZN(lce_data_cmd_o[424]));
 OAI21_X1 _48464_ (.A(_20847_),
    .B1(_20850_),
    .B2(\icache.lce.lce_cmd_inst.data_r [419]),
    .ZN(_20853_));
 AOI21_X4 _48465_ (.A(_20853_),
    .B1(_16071_),
    .B2(_20842_),
    .ZN(lce_data_cmd_o[425]));
 OAI21_X2 _48466_ (.A(_20847_),
    .B1(_20850_),
    .B2(\icache.lce.lce_cmd_inst.data_r [420]),
    .ZN(_20854_));
 BUF_X16 _48467_ (.A(_20763_),
    .Z(_20855_));
 AOI21_X4 _48468_ (.A(_20854_),
    .B1(_16094_),
    .B2(_20855_),
    .ZN(lce_data_cmd_o[426]));
 OAI21_X2 _48469_ (.A(_20847_),
    .B1(_20850_),
    .B2(\icache.lce.lce_cmd_inst.data_r [421]),
    .ZN(_20856_));
 AOI21_X4 _48470_ (.A(_20856_),
    .B1(_16116_),
    .B2(_20855_),
    .ZN(lce_data_cmd_o[427]));
 OAI21_X2 _48471_ (.A(_20847_),
    .B1(_20850_),
    .B2(\icache.lce.lce_cmd_inst.data_r [422]),
    .ZN(_20857_));
 AOI21_X4 _48472_ (.A(_20857_),
    .B1(_16134_),
    .B2(_20855_),
    .ZN(lce_data_cmd_o[428]));
 OAI21_X2 _48473_ (.A(_20847_),
    .B1(_20850_),
    .B2(\icache.lce.lce_cmd_inst.data_r [423]),
    .ZN(_20858_));
 AOI21_X4 _48474_ (.A(_20858_),
    .B1(_16153_),
    .B2(_20855_),
    .ZN(lce_data_cmd_o[429]));
 OAI21_X2 _48475_ (.A(_20847_),
    .B1(_20850_),
    .B2(\icache.lce.lce_cmd_inst.data_r [424]),
    .ZN(_20859_));
 AOI21_X4 _48476_ (.A(_20859_),
    .B1(_16173_),
    .B2(_20855_),
    .ZN(lce_data_cmd_o[430]));
 BUF_X8 _48477_ (.A(_20740_),
    .Z(_20860_));
 OAI21_X1 _48478_ (.A(_20860_),
    .B1(_20850_),
    .B2(\icache.lce.lce_cmd_inst.data_r [425]),
    .ZN(_20861_));
 AOI21_X4 _48479_ (.A(_20861_),
    .B1(_16198_),
    .B2(_20855_),
    .ZN(lce_data_cmd_o[431]));
 OAI21_X2 _48480_ (.A(_20860_),
    .B1(_20850_),
    .B2(\icache.lce.lce_cmd_inst.data_r [426]),
    .ZN(_20862_));
 AOI21_X4 _48481_ (.A(_20862_),
    .B1(_16220_),
    .B2(_20855_),
    .ZN(lce_data_cmd_o[432]));
 BUF_X16 _48482_ (.A(_20744_),
    .Z(_20863_));
 OAI21_X2 _48483_ (.A(_20860_),
    .B1(_20863_),
    .B2(\icache.lce.lce_cmd_inst.data_r [427]),
    .ZN(_20864_));
 AOI21_X4 _48484_ (.A(_20864_),
    .B1(_16249_),
    .B2(_20855_),
    .ZN(lce_data_cmd_o[433]));
 OAI21_X2 _48485_ (.A(_20860_),
    .B1(_20863_),
    .B2(\icache.lce.lce_cmd_inst.data_r [428]),
    .ZN(_20865_));
 AOI21_X4 _48486_ (.A(_20865_),
    .B1(_16278_),
    .B2(_20855_),
    .ZN(lce_data_cmd_o[434]));
 OAI21_X2 _48487_ (.A(_20860_),
    .B1(_20863_),
    .B2(\icache.lce.lce_cmd_inst.data_r [429]),
    .ZN(_20866_));
 AOI21_X4 _48488_ (.A(_20866_),
    .B1(_16296_),
    .B2(_20855_),
    .ZN(lce_data_cmd_o[435]));
 OAI21_X2 _48489_ (.A(_20860_),
    .B1(_20863_),
    .B2(\icache.lce.lce_cmd_inst.data_r [430]),
    .ZN(_20867_));
 BUF_X16 _48490_ (.A(_20763_),
    .Z(_20868_));
 AOI21_X4 _48491_ (.A(_20867_),
    .B1(_16316_),
    .B2(_20868_),
    .ZN(lce_data_cmd_o[436]));
 OAI21_X2 _48492_ (.A(_20860_),
    .B1(_20863_),
    .B2(\icache.lce.lce_cmd_inst.data_r [431]),
    .ZN(_20869_));
 AOI21_X4 _48493_ (.A(_20869_),
    .B1(_16335_),
    .B2(_20868_),
    .ZN(lce_data_cmd_o[437]));
 OAI21_X2 _48494_ (.A(_20860_),
    .B1(_20863_),
    .B2(\icache.lce.lce_cmd_inst.data_r [432]),
    .ZN(_20870_));
 AOI21_X4 _48495_ (.A(_20870_),
    .B1(_16358_),
    .B2(_20868_),
    .ZN(lce_data_cmd_o[438]));
 OAI21_X2 _48496_ (.A(_20860_),
    .B1(_20863_),
    .B2(\icache.lce.lce_cmd_inst.data_r [433]),
    .ZN(_20871_));
 AOI21_X4 _48497_ (.A(_20871_),
    .B1(_16377_),
    .B2(_20868_),
    .ZN(lce_data_cmd_o[439]));
 OAI21_X2 _48498_ (.A(_20860_),
    .B1(_20863_),
    .B2(\icache.lce.lce_cmd_inst.data_r [434]),
    .ZN(_20872_));
 AOI21_X4 _48499_ (.A(_20872_),
    .B1(_16399_),
    .B2(_20868_),
    .ZN(lce_data_cmd_o[440]));
 BUF_X8 _48500_ (.A(_07608_),
    .Z(_20873_));
 OAI21_X2 _48501_ (.A(_20873_),
    .B1(_20863_),
    .B2(\icache.lce.lce_cmd_inst.data_r [435]),
    .ZN(_20874_));
 AOI21_X4 _48502_ (.A(_20874_),
    .B1(_16421_),
    .B2(_20868_),
    .ZN(lce_data_cmd_o[441]));
 OAI21_X2 _48503_ (.A(_20873_),
    .B1(_20863_),
    .B2(\icache.lce.lce_cmd_inst.data_r [436]),
    .ZN(_20875_));
 AOI21_X4 _48504_ (.A(_20875_),
    .B1(_16436_),
    .B2(_20868_),
    .ZN(lce_data_cmd_o[442]));
 BUF_X16 _48505_ (.A(_20363_),
    .Z(_20876_));
 OAI21_X1 _48506_ (.A(_20873_),
    .B1(_20876_),
    .B2(\icache.lce.lce_cmd_inst.data_r [437]),
    .ZN(_20877_));
 AOI21_X4 _48507_ (.A(_20877_),
    .B1(_16454_),
    .B2(_20868_),
    .ZN(lce_data_cmd_o[443]));
 OAI21_X2 _48508_ (.A(_20873_),
    .B1(_20876_),
    .B2(\icache.lce.lce_cmd_inst.data_r [438]),
    .ZN(_20878_));
 AOI21_X4 _48509_ (.A(_20878_),
    .B1(_16473_),
    .B2(_20868_),
    .ZN(lce_data_cmd_o[444]));
 OAI21_X2 _48510_ (.A(_20873_),
    .B1(_20876_),
    .B2(\icache.lce.lce_cmd_inst.data_r [439]),
    .ZN(_20879_));
 AOI21_X4 _48511_ (.A(_20879_),
    .B1(_16489_),
    .B2(_20868_),
    .ZN(lce_data_cmd_o[445]));
 OAI21_X2 _48512_ (.A(_20873_),
    .B1(_20876_),
    .B2(\icache.lce.lce_cmd_inst.data_r [440]),
    .ZN(_20880_));
 BUF_X16 _48513_ (.A(_20763_),
    .Z(_20881_));
 AOI21_X4 _48514_ (.A(_20880_),
    .B1(_16507_),
    .B2(_20881_),
    .ZN(lce_data_cmd_o[446]));
 OAI21_X2 _48515_ (.A(_20873_),
    .B1(_20876_),
    .B2(\icache.lce.lce_cmd_inst.data_r [441]),
    .ZN(_20882_));
 AOI21_X4 _48516_ (.A(_20882_),
    .B1(_16527_),
    .B2(_20881_),
    .ZN(lce_data_cmd_o[447]));
 OAI21_X2 _48517_ (.A(_20873_),
    .B1(_20876_),
    .B2(\icache.lce.lce_cmd_inst.data_r [442]),
    .ZN(_20883_));
 AOI21_X4 _48518_ (.A(_20883_),
    .B1(_16549_),
    .B2(_20881_),
    .ZN(lce_data_cmd_o[448]));
 OAI21_X2 _48519_ (.A(_20873_),
    .B1(_20876_),
    .B2(\icache.lce.lce_cmd_inst.data_r [443]),
    .ZN(_20884_));
 AOI21_X4 _48520_ (.A(_20884_),
    .B1(_16574_),
    .B2(_20881_),
    .ZN(lce_data_cmd_o[449]));
 OAI21_X1 _48521_ (.A(_20873_),
    .B1(_20876_),
    .B2(\icache.lce.lce_cmd_inst.data_r [444]),
    .ZN(_20885_));
 AOI21_X4 _48522_ (.A(_20885_),
    .B1(_16594_),
    .B2(_20881_),
    .ZN(lce_data_cmd_o[450]));
 BUF_X8 _48523_ (.A(_07608_),
    .Z(_20886_));
 OAI21_X2 _48524_ (.A(_20886_),
    .B1(_20876_),
    .B2(\icache.lce.lce_cmd_inst.data_r [445]),
    .ZN(_20887_));
 AOI21_X4 _48525_ (.A(_20887_),
    .B1(_16612_),
    .B2(_20881_),
    .ZN(lce_data_cmd_o[451]));
 OAI21_X2 _48526_ (.A(_20886_),
    .B1(_20876_),
    .B2(\icache.lce.lce_cmd_inst.data_r [446]),
    .ZN(_20888_));
 AOI21_X4 _48527_ (.A(_20888_),
    .B1(_16629_),
    .B2(_20881_),
    .ZN(lce_data_cmd_o[452]));
 BUF_X8 _48528_ (.A(_20363_),
    .Z(_20889_));
 OAI21_X2 _48529_ (.A(_20886_),
    .B1(_20889_),
    .B2(\icache.lce.lce_cmd_inst.data_r [447]),
    .ZN(_20890_));
 AOI21_X4 _48530_ (.A(_20890_),
    .B1(_16649_),
    .B2(_20881_),
    .ZN(lce_data_cmd_o[453]));
 OAI21_X4 _48531_ (.A(_20886_),
    .B1(_20889_),
    .B2(\icache.lce.lce_cmd_inst.data_r [448]),
    .ZN(_20891_));
 AOI21_X4 _48532_ (.A(_20891_),
    .B1(_16665_),
    .B2(_20881_),
    .ZN(lce_data_cmd_o[454]));
 OAI21_X2 _48533_ (.A(_20886_),
    .B1(_20889_),
    .B2(\icache.lce.lce_cmd_inst.data_r [449]),
    .ZN(_20892_));
 AOI21_X4 _48534_ (.A(_20892_),
    .B1(_16683_),
    .B2(_20881_),
    .ZN(lce_data_cmd_o[455]));
 OAI21_X2 _48535_ (.A(_20886_),
    .B1(_20889_),
    .B2(\icache.lce.lce_cmd_inst.data_r [450]),
    .ZN(_20893_));
 BUF_X16 _48536_ (.A(_15296_),
    .Z(_20894_));
 AOI21_X4 _48537_ (.A(_20893_),
    .B1(_16702_),
    .B2(_20894_),
    .ZN(lce_data_cmd_o[456]));
 OAI21_X2 _48538_ (.A(_20886_),
    .B1(_20889_),
    .B2(\icache.lce.lce_cmd_inst.data_r [451]),
    .ZN(_20895_));
 AOI21_X4 _48539_ (.A(_20895_),
    .B1(_16723_),
    .B2(_20894_),
    .ZN(lce_data_cmd_o[457]));
 OAI21_X1 _48540_ (.A(_20886_),
    .B1(_20889_),
    .B2(\icache.lce.lce_cmd_inst.data_r [452]),
    .ZN(_20896_));
 AOI21_X4 _48541_ (.A(_20896_),
    .B1(_16746_),
    .B2(_20894_),
    .ZN(lce_data_cmd_o[458]));
 OAI21_X2 _48542_ (.A(_20886_),
    .B1(_20889_),
    .B2(\icache.lce.lce_cmd_inst.data_r [453]),
    .ZN(_20897_));
 AOI21_X4 _48543_ (.A(_20897_),
    .B1(_16766_),
    .B2(_20894_),
    .ZN(lce_data_cmd_o[459]));
 OAI21_X2 _48544_ (.A(_20886_),
    .B1(_20889_),
    .B2(\icache.lce.lce_cmd_inst.data_r [454]),
    .ZN(_20898_));
 AOI21_X4 _48545_ (.A(_20898_),
    .B1(_16784_),
    .B2(_20894_),
    .ZN(lce_data_cmd_o[460]));
 BUF_X4 _48546_ (.A(_07608_),
    .Z(_20899_));
 OAI21_X1 _48547_ (.A(_20899_),
    .B1(_20889_),
    .B2(\icache.lce.lce_cmd_inst.data_r [455]),
    .ZN(_20900_));
 AOI21_X4 _48548_ (.A(_20900_),
    .B1(_16809_),
    .B2(_20894_),
    .ZN(lce_data_cmd_o[461]));
 OAI21_X2 _48549_ (.A(_20899_),
    .B1(_20889_),
    .B2(\icache.lce.lce_cmd_inst.data_r [456]),
    .ZN(_20901_));
 AOI21_X4 _48550_ (.A(_20901_),
    .B1(_16829_),
    .B2(_20894_),
    .ZN(lce_data_cmd_o[462]));
 BUF_X8 _48551_ (.A(_20363_),
    .Z(_20902_));
 OAI21_X2 _48552_ (.A(_20899_),
    .B1(_20902_),
    .B2(\icache.lce.lce_cmd_inst.data_r [457]),
    .ZN(_20903_));
 AOI21_X4 _48553_ (.A(_20903_),
    .B1(_16851_),
    .B2(_20894_),
    .ZN(lce_data_cmd_o[463]));
 OAI21_X2 _48554_ (.A(_20899_),
    .B1(_20902_),
    .B2(\icache.lce.lce_cmd_inst.data_r [458]),
    .ZN(_20904_));
 AOI21_X4 _48555_ (.A(_20904_),
    .B1(_16876_),
    .B2(_20894_),
    .ZN(lce_data_cmd_o[464]));
 OAI21_X2 _48556_ (.A(_20899_),
    .B1(_20902_),
    .B2(\icache.lce.lce_cmd_inst.data_r [459]),
    .ZN(_20905_));
 AOI21_X4 _48557_ (.A(_20905_),
    .B1(_16895_),
    .B2(_20894_),
    .ZN(lce_data_cmd_o[465]));
 OAI21_X2 _48558_ (.A(_20899_),
    .B1(_20902_),
    .B2(\icache.lce.lce_cmd_inst.data_r [460]),
    .ZN(_20906_));
 BUF_X16 _48559_ (.A(_15296_),
    .Z(_20907_));
 AOI21_X4 _48560_ (.A(_20906_),
    .B1(_16913_),
    .B2(_20907_),
    .ZN(lce_data_cmd_o[466]));
 OAI21_X2 _48561_ (.A(_20899_),
    .B1(_20902_),
    .B2(\icache.lce.lce_cmd_inst.data_r [461]),
    .ZN(_20908_));
 AOI21_X4 _48562_ (.A(_20908_),
    .B1(_16934_),
    .B2(_20907_),
    .ZN(lce_data_cmd_o[467]));
 OAI21_X2 _48563_ (.A(_20899_),
    .B1(_20902_),
    .B2(\icache.lce.lce_cmd_inst.data_r [462]),
    .ZN(_20909_));
 AOI21_X4 _48564_ (.A(_20909_),
    .B1(_16954_),
    .B2(_20907_),
    .ZN(lce_data_cmd_o[468]));
 OAI21_X1 _48565_ (.A(_20899_),
    .B1(_20902_),
    .B2(\icache.lce.lce_cmd_inst.data_r [463]),
    .ZN(_20910_));
 AOI21_X4 _48566_ (.A(_20910_),
    .B1(_16976_),
    .B2(_20907_),
    .ZN(lce_data_cmd_o[469]));
 OAI21_X2 _48567_ (.A(_20899_),
    .B1(_20902_),
    .B2(\icache.lce.lce_cmd_inst.data_r [464]),
    .ZN(_20911_));
 AOI21_X4 _48568_ (.A(_20911_),
    .B1(_16996_),
    .B2(_20907_),
    .ZN(lce_data_cmd_o[470]));
 BUF_X8 _48569_ (.A(_07608_),
    .Z(_20912_));
 OAI21_X2 _48570_ (.A(_20912_),
    .B1(_20902_),
    .B2(\icache.lce.lce_cmd_inst.data_r [465]),
    .ZN(_20913_));
 AOI21_X4 _48571_ (.A(_20913_),
    .B1(_17022_),
    .B2(_20907_),
    .ZN(lce_data_cmd_o[471]));
 OAI21_X2 _48572_ (.A(_20912_),
    .B1(_20902_),
    .B2(\icache.lce.lce_cmd_inst.data_r [466]),
    .ZN(_20914_));
 AOI21_X4 _48573_ (.A(_20914_),
    .B1(_17043_),
    .B2(_20907_),
    .ZN(lce_data_cmd_o[472]));
 BUF_X8 _48574_ (.A(_20363_),
    .Z(_20915_));
 OAI21_X2 _48575_ (.A(_20912_),
    .B1(_20915_),
    .B2(\icache.lce.lce_cmd_inst.data_r [467]),
    .ZN(_20916_));
 AOI21_X4 _48576_ (.A(_20916_),
    .B1(_17064_),
    .B2(_20907_),
    .ZN(lce_data_cmd_o[473]));
 OAI21_X2 _48577_ (.A(_20912_),
    .B1(_20915_),
    .B2(\icache.lce.lce_cmd_inst.data_r [468]),
    .ZN(_20917_));
 AOI21_X4 _48578_ (.A(_20917_),
    .B1(_17086_),
    .B2(_20907_),
    .ZN(lce_data_cmd_o[474]));
 OAI21_X2 _48579_ (.A(_20912_),
    .B1(_20915_),
    .B2(\icache.lce.lce_cmd_inst.data_r [469]),
    .ZN(_20918_));
 AOI21_X4 _48580_ (.A(_20918_),
    .B1(_17107_),
    .B2(_20907_),
    .ZN(lce_data_cmd_o[475]));
 OAI21_X2 _48581_ (.A(_20912_),
    .B1(_20915_),
    .B2(\icache.lce.lce_cmd_inst.data_r [470]),
    .ZN(_20919_));
 BUF_X16 _48582_ (.A(_15296_),
    .Z(_20920_));
 AOI21_X4 _48583_ (.A(_20919_),
    .B1(_17125_),
    .B2(_20920_),
    .ZN(lce_data_cmd_o[476]));
 OAI21_X2 _48584_ (.A(_20912_),
    .B1(_20915_),
    .B2(\icache.lce.lce_cmd_inst.data_r [471]),
    .ZN(_20921_));
 AOI21_X4 _48585_ (.A(_20921_),
    .B1(_17148_),
    .B2(_20920_),
    .ZN(lce_data_cmd_o[477]));
 OAI21_X2 _48586_ (.A(_20912_),
    .B1(_20915_),
    .B2(\icache.lce.lce_cmd_inst.data_r [472]),
    .ZN(_20922_));
 AOI21_X4 _48587_ (.A(_20922_),
    .B1(_17171_),
    .B2(_20920_),
    .ZN(lce_data_cmd_o[478]));
 OAI21_X2 _48588_ (.A(_20912_),
    .B1(_20915_),
    .B2(\icache.lce.lce_cmd_inst.data_r [473]),
    .ZN(_20923_));
 AOI21_X4 _48589_ (.A(_20923_),
    .B1(_17195_),
    .B2(_20920_),
    .ZN(lce_data_cmd_o[479]));
 OAI21_X2 _48590_ (.A(_20912_),
    .B1(_20915_),
    .B2(\icache.lce.lce_cmd_inst.data_r [474]),
    .ZN(_20924_));
 AOI21_X4 _48591_ (.A(_20924_),
    .B1(_17216_),
    .B2(_20920_),
    .ZN(lce_data_cmd_o[480]));
 BUF_X8 _48592_ (.A(_07608_),
    .Z(_20925_));
 OAI21_X2 _48593_ (.A(_20925_),
    .B1(_20915_),
    .B2(\icache.lce.lce_cmd_inst.data_r [475]),
    .ZN(_20926_));
 AOI21_X4 _48594_ (.A(_20926_),
    .B1(_17239_),
    .B2(_20920_),
    .ZN(lce_data_cmd_o[481]));
 OAI21_X2 _48595_ (.A(_20925_),
    .B1(_20915_),
    .B2(\icache.lce.lce_cmd_inst.data_r [476]),
    .ZN(_20927_));
 AOI21_X4 _48596_ (.A(_20927_),
    .B1(_17259_),
    .B2(_20920_),
    .ZN(lce_data_cmd_o[482]));
 BUF_X8 _48597_ (.A(_20363_),
    .Z(_20928_));
 OAI21_X2 _48598_ (.A(_20925_),
    .B1(_20928_),
    .B2(\icache.lce.lce_cmd_inst.data_r [477]),
    .ZN(_20929_));
 AOI21_X4 _48599_ (.A(_20929_),
    .B1(_17280_),
    .B2(_20920_),
    .ZN(lce_data_cmd_o[483]));
 OAI21_X2 _48600_ (.A(_20925_),
    .B1(_20928_),
    .B2(\icache.lce.lce_cmd_inst.data_r [478]),
    .ZN(_20930_));
 AOI21_X4 _48601_ (.A(_20930_),
    .B1(_17298_),
    .B2(_20920_),
    .ZN(lce_data_cmd_o[484]));
 OAI21_X2 _48602_ (.A(_20925_),
    .B1(_20928_),
    .B2(\icache.lce.lce_cmd_inst.data_r [479]),
    .ZN(_20931_));
 AOI21_X4 _48603_ (.A(_20931_),
    .B1(_17317_),
    .B2(_20920_),
    .ZN(lce_data_cmd_o[485]));
 OAI21_X2 _48604_ (.A(_20925_),
    .B1(_20928_),
    .B2(\icache.lce.lce_cmd_inst.data_r [480]),
    .ZN(_20932_));
 BUF_X16 _48605_ (.A(_15296_),
    .Z(_20933_));
 AOI21_X4 _48606_ (.A(_20932_),
    .B1(_17336_),
    .B2(_20933_),
    .ZN(lce_data_cmd_o[486]));
 OAI21_X2 _48607_ (.A(_20925_),
    .B1(_20928_),
    .B2(\icache.lce.lce_cmd_inst.data_r [481]),
    .ZN(_20934_));
 AOI21_X4 _48608_ (.A(_20934_),
    .B1(_17353_),
    .B2(_20933_),
    .ZN(lce_data_cmd_o[487]));
 OAI21_X1 _48609_ (.A(_20925_),
    .B1(_20928_),
    .B2(\icache.lce.lce_cmd_inst.data_r [482]),
    .ZN(_20935_));
 AOI21_X4 _48610_ (.A(_20935_),
    .B1(_17368_),
    .B2(_20933_),
    .ZN(lce_data_cmd_o[488]));
 OAI21_X2 _48611_ (.A(_20925_),
    .B1(_20928_),
    .B2(\icache.lce.lce_cmd_inst.data_r [483]),
    .ZN(_20936_));
 AOI21_X4 _48612_ (.A(_20936_),
    .B1(_17388_),
    .B2(_20933_),
    .ZN(lce_data_cmd_o[489]));
 OAI21_X2 _48613_ (.A(_20925_),
    .B1(_20928_),
    .B2(\icache.lce.lce_cmd_inst.data_r [484]),
    .ZN(_20937_));
 AOI21_X4 _48614_ (.A(_20937_),
    .B1(_17403_),
    .B2(_20933_),
    .ZN(lce_data_cmd_o[490]));
 BUF_X8 _48615_ (.A(_07608_),
    .Z(_20938_));
 OAI21_X2 _48616_ (.A(_20938_),
    .B1(_20928_),
    .B2(\icache.lce.lce_cmd_inst.data_r [485]),
    .ZN(_20939_));
 AOI21_X4 _48617_ (.A(_20939_),
    .B1(_17423_),
    .B2(_20933_),
    .ZN(lce_data_cmd_o[491]));
 OAI21_X2 _48618_ (.A(_20938_),
    .B1(_20928_),
    .B2(\icache.lce.lce_cmd_inst.data_r [486]),
    .ZN(_20940_));
 AOI21_X4 _48619_ (.A(_20940_),
    .B1(_17441_),
    .B2(_20933_),
    .ZN(lce_data_cmd_o[492]));
 BUF_X8 _48620_ (.A(_20363_),
    .Z(_20941_));
 OAI21_X2 _48621_ (.A(_20938_),
    .B1(_20941_),
    .B2(\icache.lce.lce_cmd_inst.data_r [487]),
    .ZN(_20942_));
 AOI21_X4 _48622_ (.A(_20942_),
    .B1(_17457_),
    .B2(_20933_),
    .ZN(lce_data_cmd_o[493]));
 OAI21_X2 _48623_ (.A(_20938_),
    .B1(_20941_),
    .B2(\icache.lce.lce_cmd_inst.data_r [488]),
    .ZN(_20943_));
 AOI21_X4 _48624_ (.A(_20943_),
    .B1(_17473_),
    .B2(_20933_),
    .ZN(lce_data_cmd_o[494]));
 OAI21_X2 _48625_ (.A(_20938_),
    .B1(_20941_),
    .B2(\icache.lce.lce_cmd_inst.data_r [489]),
    .ZN(_20944_));
 AOI21_X4 _48626_ (.A(_20944_),
    .B1(_17488_),
    .B2(_20933_),
    .ZN(lce_data_cmd_o[495]));
 OAI21_X2 _48627_ (.A(_20938_),
    .B1(_20941_),
    .B2(\icache.lce.lce_cmd_inst.data_r [490]),
    .ZN(_20945_));
 BUF_X16 _48628_ (.A(_15296_),
    .Z(_20946_));
 AOI21_X4 _48629_ (.A(_20945_),
    .B1(_17525_),
    .B2(_20946_),
    .ZN(lce_data_cmd_o[496]));
 OAI21_X2 _48630_ (.A(_20938_),
    .B1(_20941_),
    .B2(\icache.lce.lce_cmd_inst.data_r [491]),
    .ZN(_20947_));
 AOI21_X4 _48631_ (.A(_20947_),
    .B1(_17545_),
    .B2(_20946_),
    .ZN(lce_data_cmd_o[497]));
 OAI21_X2 _48632_ (.A(_20938_),
    .B1(_20941_),
    .B2(\icache.lce.lce_cmd_inst.data_r [492]),
    .ZN(_20948_));
 AOI21_X4 _48633_ (.A(_20948_),
    .B1(_17562_),
    .B2(_20946_),
    .ZN(lce_data_cmd_o[498]));
 OAI21_X2 _48634_ (.A(_20938_),
    .B1(_20941_),
    .B2(\icache.lce.lce_cmd_inst.data_r [493]),
    .ZN(_20949_));
 AOI21_X4 _48635_ (.A(_20949_),
    .B1(_15530_),
    .B2(_20946_),
    .ZN(lce_data_cmd_o[499]));
 OAI21_X2 _48636_ (.A(_20938_),
    .B1(_20941_),
    .B2(\icache.lce.lce_cmd_inst.data_r [494]),
    .ZN(_20950_));
 AOI21_X4 _48637_ (.A(_20950_),
    .B1(_15560_),
    .B2(_20946_),
    .ZN(lce_data_cmd_o[500]));
 BUF_X8 _48638_ (.A(_07608_),
    .Z(_20951_));
 OAI21_X2 _48639_ (.A(_20951_),
    .B1(_20941_),
    .B2(\icache.lce.lce_cmd_inst.data_r [495]),
    .ZN(_20952_));
 AOI21_X4 _48640_ (.A(_20952_),
    .B1(_15600_),
    .B2(_20946_),
    .ZN(lce_data_cmd_o[501]));
 OAI21_X2 _48641_ (.A(_20951_),
    .B1(_20941_),
    .B2(\icache.lce.lce_cmd_inst.data_r [496]),
    .ZN(_20953_));
 AOI21_X4 _48642_ (.A(_20953_),
    .B1(_15634_),
    .B2(_20946_),
    .ZN(lce_data_cmd_o[502]));
 BUF_X16 _48643_ (.A(_20363_),
    .Z(_20954_));
 OAI21_X2 _48644_ (.A(_20951_),
    .B1(_20954_),
    .B2(\icache.lce.lce_cmd_inst.data_r [497]),
    .ZN(_20955_));
 AOI21_X4 _48645_ (.A(_20955_),
    .B1(_15658_),
    .B2(_20946_),
    .ZN(lce_data_cmd_o[503]));
 OAI21_X2 _48646_ (.A(_20951_),
    .B1(_20954_),
    .B2(\icache.lce.lce_cmd_inst.data_r [498]),
    .ZN(_20956_));
 AOI21_X4 _48647_ (.A(_20956_),
    .B1(_15683_),
    .B2(_20946_),
    .ZN(lce_data_cmd_o[504]));
 OAI21_X1 _48648_ (.A(_20951_),
    .B1(_20954_),
    .B2(\icache.lce.lce_cmd_inst.data_r [499]),
    .ZN(_20957_));
 AOI21_X4 _48649_ (.A(_20957_),
    .B1(_15706_),
    .B2(_20946_),
    .ZN(lce_data_cmd_o[505]));
 OAI21_X1 _48650_ (.A(_20951_),
    .B1(_20954_),
    .B2(\icache.lce.lce_cmd_inst.data_r [500]),
    .ZN(_20958_));
 BUF_X32 _48651_ (.A(_15296_),
    .Z(_20959_));
 AOI21_X4 _48652_ (.A(_20958_),
    .B1(_15732_),
    .B2(_20959_),
    .ZN(lce_data_cmd_o[506]));
 OAI21_X2 _48653_ (.A(_20951_),
    .B1(_20954_),
    .B2(\icache.lce.lce_cmd_inst.data_r [501]),
    .ZN(_20960_));
 AOI21_X4 _48654_ (.A(_20960_),
    .B1(_15764_),
    .B2(_20959_),
    .ZN(lce_data_cmd_o[507]));
 OAI21_X2 _48655_ (.A(_20951_),
    .B1(_20954_),
    .B2(\icache.lce.lce_cmd_inst.data_r [502]),
    .ZN(_20961_));
 AOI21_X4 _48656_ (.A(_20961_),
    .B1(_15792_),
    .B2(_20959_),
    .ZN(lce_data_cmd_o[508]));
 OAI21_X2 _48657_ (.A(_20951_),
    .B1(_20954_),
    .B2(\icache.lce.lce_cmd_inst.data_r [503]),
    .ZN(_20962_));
 AOI21_X4 _48658_ (.A(_20962_),
    .B1(_15821_),
    .B2(_20959_),
    .ZN(lce_data_cmd_o[509]));
 OAI21_X2 _48659_ (.A(_20951_),
    .B1(_20954_),
    .B2(\icache.lce.lce_cmd_inst.data_r [504]),
    .ZN(_20963_));
 AOI21_X4 _48660_ (.A(_20963_),
    .B1(_15851_),
    .B2(_20959_),
    .ZN(lce_data_cmd_o[510]));
 OAI21_X2 _48661_ (.A(_20300_),
    .B1(_20954_),
    .B2(\icache.lce.lce_cmd_inst.data_r [505]),
    .ZN(_20964_));
 AOI21_X4 _48662_ (.A(_20964_),
    .B1(_15872_),
    .B2(_20959_),
    .ZN(lce_data_cmd_o[511]));
 OAI21_X1 _48663_ (.A(_20300_),
    .B1(_20954_),
    .B2(\icache.lce.lce_cmd_inst.data_r [506]),
    .ZN(_20965_));
 AOI21_X4 _48664_ (.A(_20965_),
    .B1(_15899_),
    .B2(_20959_),
    .ZN(lce_data_cmd_o[512]));
 OAI21_X2 _48665_ (.A(_20300_),
    .B1(_20294_),
    .B2(\icache.lce.lce_cmd_inst.data_r [507]),
    .ZN(_20966_));
 AOI21_X4 _48666_ (.A(_20966_),
    .B1(_17508_),
    .B2(_20959_),
    .ZN(lce_data_cmd_o[513]));
 OAI21_X1 _48667_ (.A(_20300_),
    .B1(_20294_),
    .B2(\icache.lce.lce_cmd_inst.data_r [508]),
    .ZN(_20967_));
 AOI21_X4 _48668_ (.A(_20967_),
    .B1(_15500_),
    .B2(_20959_),
    .ZN(lce_data_cmd_o[514]));
 OAI21_X2 _48669_ (.A(_20300_),
    .B1(_20294_),
    .B2(\icache.lce.lce_cmd_inst.data_r [509]),
    .ZN(_20968_));
 AOI21_X4 _48670_ (.A(_20968_),
    .B1(_15467_),
    .B2(_20959_),
    .ZN(lce_data_cmd_o[515]));
 OAI21_X2 _48671_ (.A(_20300_),
    .B1(_20294_),
    .B2(\icache.lce.lce_cmd_inst.data_r [510]),
    .ZN(_20969_));
 AOI21_X4 _48672_ (.A(_20969_),
    .B1(_15428_),
    .B2(_15297_),
    .ZN(lce_data_cmd_o[516]));
 OAI21_X2 _48673_ (.A(_20300_),
    .B1(_20294_),
    .B2(\icache.lce.lce_cmd_inst.data_r [511]),
    .ZN(_20970_));
 AOI21_X4 _48674_ (.A(_20970_),
    .B1(_15385_),
    .B2(_15297_),
    .ZN(lce_data_cmd_o[517]));
 BUF_X8 _48675_ (.A(_07977_),
    .Z(_20971_));
 AND4_X4 _48676_ (.A1(_00001_),
    .A2(_08421_),
    .A3(_20971_),
    .A4(_07972_),
    .ZN(lce_data_resp_v_o));
 AND2_X4 _48677_ (.A1(_08421_),
    .A2(_07977_),
    .ZN(_20972_));
 INV_X4 _48678_ (.A(_20972_),
    .ZN(_20973_));
 BUF_X16 _48679_ (.A(_20973_),
    .Z(_20974_));
 BUF_X16 _48680_ (.A(_07892_),
    .Z(_20975_));
 NOR3_X4 _48681_ (.A1(_20974_),
    .A2(_20975_),
    .A3(_10654_),
    .ZN(lce_data_resp_o[0]));
 NOR3_X4 _48682_ (.A1(_20974_),
    .A2(_20975_),
    .A3(_10661_),
    .ZN(lce_data_resp_o[1]));
 NOR3_X4 _48683_ (.A1(_20974_),
    .A2(_20975_),
    .A3(_10665_),
    .ZN(lce_data_resp_o[2]));
 NOR3_X4 _48684_ (.A1(_20974_),
    .A2(_20975_),
    .A3(_10669_),
    .ZN(lce_data_resp_o[3]));
 BUF_X8 _48685_ (.A(_20972_),
    .Z(_20976_));
 AND4_X4 _48686_ (.A1(_07939_),
    .A2(_20976_),
    .A3(_10672_),
    .A4(_10673_),
    .ZN(lce_data_resp_o[4]));
 AND4_X4 _48687_ (.A1(_07939_),
    .A2(_20976_),
    .A3(_10675_),
    .A4(_10676_),
    .ZN(lce_data_resp_o[5]));
 AND4_X4 _48688_ (.A1(_07626_),
    .A2(_08421_),
    .A3(_20971_),
    .A4(_07896_),
    .ZN(lce_data_resp_o[6]));
 AND4_X4 _48689_ (.A1(_20971_),
    .A2(_08421_),
    .A3(_07632_),
    .A4(_07896_),
    .ZN(lce_data_resp_o[7]));
 AND4_X4 _48690_ (.A1(_20971_),
    .A2(_08421_),
    .A3(_07637_),
    .A4(_07896_),
    .ZN(lce_data_resp_o[8]));
 AND4_X4 _48691_ (.A1(_20971_),
    .A2(_08421_),
    .A3(_07642_),
    .A4(_07896_),
    .ZN(lce_data_resp_o[9]));
 AND4_X4 _48692_ (.A1(_20971_),
    .A2(_08421_),
    .A3(_07647_),
    .A4(_07896_),
    .ZN(lce_data_resp_o[10]));
 AND4_X4 _48693_ (.A1(_20971_),
    .A2(_08421_),
    .A3(_07652_),
    .A4(_07896_),
    .ZN(lce_data_resp_o[11]));
 BUF_X16 _48694_ (.A(_07892_),
    .Z(_20977_));
 NOR3_X4 _48695_ (.A1(_20974_),
    .A2(_07888_),
    .A3(_20977_),
    .ZN(lce_data_resp_o[12]));
 AND4_X4 _48696_ (.A1(_07939_),
    .A2(_20976_),
    .A3(_07901_),
    .A4(_07902_),
    .ZN(lce_data_resp_o[13]));
 NOR3_X4 _48697_ (.A1(_20974_),
    .A2(_20975_),
    .A3(_07905_),
    .ZN(lce_data_resp_o[14]));
 AND4_X4 _48698_ (.A1(_07939_),
    .A2(_20976_),
    .A3(_07907_),
    .A4(_07908_),
    .ZN(lce_data_resp_o[15]));
 AND4_X4 _48699_ (.A1(_07939_),
    .A2(_20976_),
    .A3(_07909_),
    .A4(_07910_),
    .ZN(lce_data_resp_o[16]));
 AND4_X4 _48700_ (.A1(_07939_),
    .A2(_20976_),
    .A3(_07911_),
    .A4(_07912_),
    .ZN(lce_data_resp_o[17]));
 NOR3_X4 _48701_ (.A1(_20974_),
    .A2(_20975_),
    .A3(_07916_),
    .ZN(lce_data_resp_o[18]));
 NOR3_X4 _48702_ (.A1(_20974_),
    .A2(_20975_),
    .A3(_07919_),
    .ZN(lce_data_resp_o[19]));
 AND4_X4 _48703_ (.A1(_07939_),
    .A2(_20976_),
    .A3(_07920_),
    .A4(_07921_),
    .ZN(lce_data_resp_o[20]));
 AND4_X4 _48704_ (.A1(_07972_),
    .A2(_20976_),
    .A3(_07922_),
    .A4(_07923_),
    .ZN(lce_data_resp_o[21]));
 NOR3_X4 _48705_ (.A1(_20974_),
    .A2(_20975_),
    .A3(_07926_),
    .ZN(lce_data_resp_o[22]));
 AND4_X4 _48706_ (.A1(_07972_),
    .A2(_20976_),
    .A3(_07927_),
    .A4(_07928_),
    .ZN(lce_data_resp_o[23]));
 AND4_X4 _48707_ (.A1(_07972_),
    .A2(_20972_),
    .A3(_07929_),
    .A4(_07930_),
    .ZN(lce_data_resp_o[24]));
 NOR3_X4 _48708_ (.A1(_20974_),
    .A2(_20975_),
    .A3(_07933_),
    .ZN(lce_data_resp_o[25]));
 BUF_X16 _48709_ (.A(_20973_),
    .Z(_20978_));
 NOR3_X4 _48710_ (.A1(_20978_),
    .A2(_20975_),
    .A3(_07936_),
    .ZN(lce_data_resp_o[26]));
 AND4_X4 _48711_ (.A1(_07972_),
    .A2(_20972_),
    .A3(_07937_),
    .A4(_07938_),
    .ZN(lce_data_resp_o[27]));
 AND4_X4 _48712_ (.A1(_07972_),
    .A2(_20972_),
    .A3(_07940_),
    .A4(_07941_),
    .ZN(lce_data_resp_o[28]));
 NOR3_X4 _48713_ (.A1(_20978_),
    .A2(_20977_),
    .A3(_07944_),
    .ZN(lce_data_resp_o[29]));
 AND4_X4 _48714_ (.A1(_07972_),
    .A2(_20972_),
    .A3(_07945_),
    .A4(_07946_),
    .ZN(lce_data_resp_o[30]));
 NOR3_X4 _48715_ (.A1(_20978_),
    .A2(_20977_),
    .A3(_07949_),
    .ZN(lce_data_resp_o[31]));
 NOR3_X4 _48716_ (.A1(_20978_),
    .A2(_20977_),
    .A3(_07952_),
    .ZN(lce_data_resp_o[32]));
 NOR3_X4 _48717_ (.A1(_20978_),
    .A2(_20977_),
    .A3(_07955_),
    .ZN(lce_data_resp_o[33]));
 NOR3_X4 _48718_ (.A1(_20978_),
    .A2(_20977_),
    .A3(_07958_),
    .ZN(lce_data_resp_o[34]));
 NOR3_X4 _48719_ (.A1(_20978_),
    .A2(_20977_),
    .A3(_07961_),
    .ZN(lce_data_resp_o[35]));
 AND4_X4 _48720_ (.A1(_07972_),
    .A2(_20972_),
    .A3(_07962_),
    .A4(_07963_),
    .ZN(lce_data_resp_o[36]));
 NOR3_X4 _48721_ (.A1(_20978_),
    .A2(_20977_),
    .A3(_07966_),
    .ZN(lce_data_resp_o[37]));
 NOR3_X4 _48722_ (.A1(_20978_),
    .A2(_20977_),
    .A3(_07969_),
    .ZN(lce_data_resp_o[38]));
 AND2_X4 _48723_ (.A1(_20976_),
    .A2(_07897_),
    .ZN(lce_data_resp_o[39]));
 NOR3_X4 _48724_ (.A1(_20978_),
    .A2(_20977_),
    .A3(_10720_),
    .ZN(lce_data_resp_o[41]));
 NAND2_X4 _48725_ (.A1(net235),
    .A2(_07898_),
    .ZN(_20979_));
 NOR2_X1 _48726_ (.A1(_20979_),
    .A2(_10678_),
    .ZN(_20980_));
 OAI21_X1 _48727_ (.A(_00601_),
    .B1(_20979_),
    .B2(_20971_),
    .ZN(_20981_));
 NOR2_X1 _48728_ (.A1(_15278_),
    .A2(_15281_),
    .ZN(_20982_));
 INV_X1 _48729_ (.A(_20982_),
    .ZN(_20983_));
 NAND2_X1 _48730_ (.A1(_15271_),
    .A2(_15272_),
    .ZN(_20984_));
 NOR3_X2 _48731_ (.A1(_20983_),
    .A2(_15270_),
    .A3(_20984_),
    .ZN(_20985_));
 INV_X1 _48732_ (.A(_00602_),
    .ZN(_20986_));
 OAI21_X1 _48733_ (.A(_20981_),
    .B1(_20985_),
    .B2(_20986_),
    .ZN(_20987_));
 NOR2_X1 _48734_ (.A1(_15278_),
    .A2(_15275_),
    .ZN(_20988_));
 INV_X1 _48735_ (.A(_20988_),
    .ZN(_20989_));
 AOI21_X1 _48736_ (.A(_20980_),
    .B1(_20987_),
    .B2(_20989_),
    .ZN(_20990_));
 AND2_X1 _48737_ (.A1(_08021_),
    .A2(\icache.lce.lce_req_inst.state_r [0]),
    .ZN(_20991_));
 INV_X1 _48738_ (.A(_20991_),
    .ZN(_20992_));
 OAI22_X2 _48739_ (.A1(_20990_),
    .A2(_20992_),
    .B1(lce_resp_ready_i),
    .B2(_10716_),
    .ZN(_20993_));
 AND2_X4 _48740_ (.A1(_08021_),
    .A2(_00002_),
    .ZN(lce_req_o[2]));
 INV_X2 _48741_ (.A(lce_req_o[2]),
    .ZN(_20994_));
 NAND2_X1 _48742_ (.A1(_20993_),
    .A2(_20994_),
    .ZN(_20995_));
 INV_X1 _48743_ (.A(_08016_),
    .ZN(_20996_));
 NOR3_X2 _48744_ (.A1(_07879_),
    .A2(\icache.N8 ),
    .A3(_20996_),
    .ZN(_20997_));
 AOI221_X4 _48745_ (.A(_20997_),
    .B1(\icache.lce.lce_req_inst.state_r [0]),
    .B2(_08014_),
    .C1(lce_req_ready_i),
    .C2(lce_req_o[2]),
    .ZN(_20998_));
 AOI21_X1 _48746_ (.A(_08651_),
    .B1(_20995_),
    .B2(_20998_),
    .ZN(_06589_));
 AND3_X1 _48747_ (.A1(_08013_),
    .A2(_00604_),
    .A3(_08016_),
    .ZN(_20999_));
 NOR2_X1 _48748_ (.A1(_20983_),
    .A2(_20984_),
    .ZN(_21000_));
 INV_X1 _48749_ (.A(_21000_),
    .ZN(_21001_));
 AND3_X1 _48750_ (.A1(_21001_),
    .A2(_00602_),
    .A3(_00603_),
    .ZN(_21002_));
 INV_X1 _48751_ (.A(_20981_),
    .ZN(_21003_));
 OAI21_X1 _48752_ (.A(_20989_),
    .B1(_10678_),
    .B2(_20979_),
    .ZN(_21004_));
 NOR3_X1 _48753_ (.A1(_21002_),
    .A2(_21003_),
    .A3(_21004_),
    .ZN(_21005_));
 OR3_X1 _48754_ (.A1(_21005_),
    .A2(_20992_),
    .A3(_20980_),
    .ZN(_21006_));
 AOI21_X1 _48755_ (.A(lce_resp_ready_i),
    .B1(_10648_),
    .B2(_10649_),
    .ZN(_21007_));
 OAI211_X2 _48756_ (.A(_21006_),
    .B(_20994_),
    .C1(_20991_),
    .C2(_21007_),
    .ZN(_21008_));
 INV_X1 _48757_ (.A(_08017_),
    .ZN(_21009_));
 AOI211_X1 _48758_ (.A(_11219_),
    .B(_20999_),
    .C1(_21008_),
    .C2(_21009_),
    .ZN(_06590_));
 AND3_X1 _48759_ (.A1(_08013_),
    .A2(_00605_),
    .A3(_08016_),
    .ZN(_21010_));
 OR4_X1 _48760_ (.A1(\icache.lce.lce_req_inst.state_r [2]),
    .A2(\icache.lce.lce_req_inst.state_r [1]),
    .A3(_00002_),
    .A4(lce_req_ready_i),
    .ZN(_21011_));
 NOR2_X1 _48761_ (.A1(_21002_),
    .A2(_21003_),
    .ZN(_21012_));
 NOR3_X1 _48762_ (.A1(_21012_),
    .A2(_20992_),
    .A3(_21004_),
    .ZN(_21013_));
 AOI21_X1 _48763_ (.A(_08019_),
    .B1(_00002_),
    .B2(_08021_),
    .ZN(_21014_));
 INV_X1 _48764_ (.A(_21014_),
    .ZN(_21015_));
 OAI21_X1 _48765_ (.A(_21011_),
    .B1(_21013_),
    .B2(_21015_),
    .ZN(_21016_));
 MUX2_X1 _48766_ (.A(_08012_),
    .B(_21016_),
    .S(_20996_),
    .Z(_21017_));
 AOI211_X1 _48767_ (.A(_11219_),
    .B(_21010_),
    .C1(_21017_),
    .C2(_21009_),
    .ZN(_06591_));
 NOR2_X1 _48768_ (.A1(_08017_),
    .A2(_21015_),
    .ZN(_21018_));
 AND2_X1 _48769_ (.A1(\icache.lce.lce_req_inst.state_r [2]),
    .A2(\icache.lce.lce_req_inst.state_r [1]),
    .ZN(_21019_));
 INV_X1 _48770_ (.A(_21019_),
    .ZN(_21020_));
 NAND3_X1 _48771_ (.A1(_10648_),
    .A2(_21020_),
    .A3(_10649_),
    .ZN(_21021_));
 INV_X1 _48772_ (.A(_21021_),
    .ZN(_21022_));
 AND2_X1 _48773_ (.A1(_21018_),
    .A2(_21022_),
    .ZN(_21023_));
 AND2_X1 _48774_ (.A1(_21023_),
    .A2(_20992_),
    .ZN(_21024_));
 AND2_X4 _48775_ (.A1(_21024_),
    .A2(_08519_),
    .ZN(_21025_));
 BUF_X8 _48776_ (.A(_21025_),
    .Z(_21026_));
 BUF_X8 _48777_ (.A(_21026_),
    .Z(_21027_));
 MUX2_X1 _48778_ (.A(\icache.lce.lce_data_cmd.miss_addr_i [0]),
    .B(\icache.addr_tv_r [0]),
    .S(_21027_),
    .Z(_06549_));
 MUX2_X1 _48779_ (.A(\icache.lce.lce_data_cmd.miss_addr_i [1]),
    .B(\icache.addr_tv_r [1]),
    .S(_21027_),
    .Z(_06560_));
 MUX2_X1 _48780_ (.A(\icache.lce.lce_data_cmd.miss_addr_i [2]),
    .B(_09308_),
    .S(_21027_),
    .Z(_06571_));
 MUX2_X1 _48781_ (.A(lce_req_o[10]),
    .B(\icache.addr_tv_r [3]),
    .S(_21027_),
    .Z(_06581_));
 MUX2_X1 _48782_ (.A(lce_req_o[11]),
    .B(\icache.addr_tv_r [4]),
    .S(_21027_),
    .Z(_06582_));
 MUX2_X1 _48783_ (.A(lce_req_o[12]),
    .B(\icache.addr_tv_r [5]),
    .S(_21027_),
    .Z(_06583_));
 MUX2_X1 _48784_ (.A(lce_req_o[13]),
    .B(\icache.addr_tv_r [6]),
    .S(_21027_),
    .Z(_06584_));
 MUX2_X1 _48785_ (.A(lce_req_o[14]),
    .B(\icache.addr_tv_r [7]),
    .S(_21027_),
    .Z(_06585_));
 MUX2_X1 _48786_ (.A(lce_req_o[15]),
    .B(\icache.addr_tv_r [8]),
    .S(_21027_),
    .Z(_06586_));
 MUX2_X1 _48787_ (.A(lce_req_o[16]),
    .B(\icache.addr_tv_r [9]),
    .S(_21027_),
    .Z(_06587_));
 BUF_X8 _48788_ (.A(_21025_),
    .Z(_21028_));
 MUX2_X1 _48789_ (.A(lce_req_o[17]),
    .B(\icache.addr_tv_r [10]),
    .S(_21028_),
    .Z(_06550_));
 MUX2_X1 _48790_ (.A(lce_req_o[18]),
    .B(\icache.addr_tv_r [11]),
    .S(_21028_),
    .Z(_06551_));
 MUX2_X1 _48791_ (.A(lce_req_o[19]),
    .B(_07193_),
    .S(_21028_),
    .Z(_06552_));
 MUX2_X1 _48792_ (.A(lce_req_o[20]),
    .B(net1380),
    .S(_21028_),
    .Z(_06553_));
 MUX2_X1 _48793_ (.A(lce_req_o[21]),
    .B(_07370_),
    .S(_21028_),
    .Z(_06554_));
 MUX2_X1 _48794_ (.A(lce_req_o[22]),
    .B(_07186_),
    .S(_21028_),
    .Z(_06555_));
 MUX2_X1 _48795_ (.A(lce_req_o[23]),
    .B(_07123_),
    .S(_21028_),
    .Z(_06556_));
 MUX2_X1 _48796_ (.A(lce_req_o[24]),
    .B(net1369),
    .S(_21028_),
    .Z(_06557_));
 MUX2_X1 _48797_ (.A(lce_req_o[25]),
    .B(_07113_),
    .S(_21028_),
    .Z(_06558_));
 MUX2_X1 _48798_ (.A(lce_req_o[26]),
    .B(net1362),
    .S(_21028_),
    .Z(_06559_));
 BUF_X8 _48799_ (.A(_21025_),
    .Z(_21029_));
 MUX2_X1 _48800_ (.A(lce_req_o[27]),
    .B(_07128_),
    .S(_21029_),
    .Z(_06561_));
 MUX2_X1 _48801_ (.A(lce_req_o[28]),
    .B(net1356),
    .S(_21029_),
    .Z(_06562_));
 MUX2_X1 _48802_ (.A(lce_req_o[29]),
    .B(_07118_),
    .S(_21029_),
    .Z(_06563_));
 MUX2_X1 _48803_ (.A(lce_req_o[30]),
    .B(net1353),
    .S(_21029_),
    .Z(_06564_));
 MUX2_X1 _48804_ (.A(lce_req_o[31]),
    .B(_07105_),
    .S(_21029_),
    .Z(_06565_));
 MUX2_X1 _48805_ (.A(lce_req_o[32]),
    .B(_07135_),
    .S(_21029_),
    .Z(_06566_));
 MUX2_X1 _48806_ (.A(lce_req_o[33]),
    .B(_07107_),
    .S(_21029_),
    .Z(_06567_));
 MUX2_X1 _48807_ (.A(lce_req_o[34]),
    .B(_07190_),
    .S(_21029_),
    .Z(_06568_));
 MUX2_X1 _48808_ (.A(lce_req_o[35]),
    .B(net1346),
    .S(_21029_),
    .Z(_06569_));
 MUX2_X1 _48809_ (.A(lce_req_o[36]),
    .B(_07248_),
    .S(_21029_),
    .Z(_06570_));
 MUX2_X1 _48810_ (.A(lce_req_o[37]),
    .B(_07130_),
    .S(_21026_),
    .Z(_06572_));
 MUX2_X1 _48811_ (.A(lce_req_o[38]),
    .B(net1336),
    .S(_21026_),
    .Z(_06573_));
 MUX2_X1 _48812_ (.A(lce_req_o[39]),
    .B(_07133_),
    .S(_21026_),
    .Z(_06574_));
 MUX2_X1 _48813_ (.A(lce_req_o[40]),
    .B(net1333),
    .S(_21026_),
    .Z(_06575_));
 MUX2_X1 _48814_ (.A(lce_req_o[41]),
    .B(_07156_),
    .S(_21026_),
    .Z(_06576_));
 MUX2_X1 _48815_ (.A(lce_req_o[42]),
    .B(net1326),
    .S(_21026_),
    .Z(_06577_));
 MUX2_X1 _48816_ (.A(lce_req_o[43]),
    .B(_07092_),
    .S(_21026_),
    .Z(_06578_));
 MUX2_X1 _48817_ (.A(lce_req_o[44]),
    .B(net1321),
    .S(_21026_),
    .Z(_06579_));
 MUX2_X1 _48818_ (.A(lce_req_o[45]),
    .B(_07160_),
    .S(_21026_),
    .Z(_06580_));
 OR2_X1 _48819_ (.A1(_21024_),
    .A2(_08650_),
    .ZN(_21030_));
 NOR3_X1 _48820_ (.A1(_20985_),
    .A2(_20986_),
    .A3(_20992_),
    .ZN(_21031_));
 INV_X1 _48821_ (.A(_21023_),
    .ZN(_21032_));
 AOI211_X1 _48822_ (.A(_21030_),
    .B(_21031_),
    .C1(_00602_),
    .C2(_21032_),
    .ZN(_06592_));
 NAND3_X1 _48823_ (.A1(_21000_),
    .A2(_15270_),
    .A3(_21023_),
    .ZN(_21033_));
 AOI21_X1 _48824_ (.A(_21030_),
    .B1(_21033_),
    .B2(_00603_),
    .ZN(_06548_));
 OR3_X1 _48825_ (.A1(_20979_),
    .A2(_20971_),
    .A3(_21032_),
    .ZN(_21034_));
 AOI21_X1 _48826_ (.A(_21030_),
    .B1(_21034_),
    .B2(_00601_),
    .ZN(_06588_));
 NOR2_X2 _48827_ (.A1(_07255_),
    .A2(_07333_),
    .ZN(_21035_));
 NOR2_X1 _48828_ (.A1(_07350_),
    .A2(_07425_),
    .ZN(_21036_));
 AND2_X4 _48829_ (.A1(_21035_),
    .A2(_21036_),
    .ZN(_21037_));
 NOR2_X4 _48830_ (.A1(_07198_),
    .A2(_07094_),
    .ZN(_21038_));
 AND2_X4 _48831_ (.A1(_21037_),
    .A2(_21038_),
    .ZN(_21039_));
 INV_X1 _48832_ (.A(\icache.lru_encoder.lru_i [1]),
    .ZN(_21040_));
 INV_X1 _48833_ (.A(\icache.lru_encode [2]),
    .ZN(_21041_));
 NAND3_X1 _48834_ (.A1(_21040_),
    .A2(_21041_),
    .A3(\icache.lru_encoder.lru_i [3]),
    .ZN(_21042_));
 NOR2_X1 _48835_ (.A1(_21041_),
    .A2(\icache.lru_encoder.lru_i [2]),
    .ZN(_21043_));
 NAND2_X1 _48836_ (.A1(_21043_),
    .A2(\icache.lru_encoder.lru_i [5]),
    .ZN(_21044_));
 NOR2_X4 _48837_ (.A1(_07501_),
    .A2(_07562_),
    .ZN(_21045_));
 NAND4_X2 _48838_ (.A1(_21039_),
    .A2(_21042_),
    .A3(_21044_),
    .A4(_21045_),
    .ZN(_21046_));
 AND3_X1 _48839_ (.A1(\icache.lru_encode [2]),
    .A2(\icache.lru_encoder.lru_i [2]),
    .A3(\icache.lru_encoder.lru_i [6]),
    .ZN(_21047_));
 AND3_X1 _48840_ (.A1(_21041_),
    .A2(\icache.lru_encoder.lru_i [1]),
    .A3(\icache.lru_encoder.lru_i [4]),
    .ZN(_21048_));
 NOR3_X4 _48841_ (.A1(_21046_),
    .A2(_21047_),
    .A3(_21048_),
    .ZN(_21049_));
 OAI21_X1 _48842_ (.A(_20994_),
    .B1(_21021_),
    .B2(_20991_),
    .ZN(_21050_));
 OAI21_X1 _48843_ (.A(_08014_),
    .B1(_08015_),
    .B2(_08018_),
    .ZN(_21051_));
 AND2_X4 _48844_ (.A1(_21050_),
    .A2(_21051_),
    .ZN(_21052_));
 OAI211_X4 _48845_ (.A(_07351_),
    .B(_07095_),
    .C1(_07502_),
    .C2(_07198_),
    .ZN(_21053_));
 AOI21_X1 _48846_ (.A(_07425_),
    .B1(_21037_),
    .B2(_21053_),
    .ZN(_21054_));
 NOR2_X1 _48847_ (.A1(_21054_),
    .A2(_07333_),
    .ZN(_21055_));
 NOR4_X4 _48848_ (.A1(_21049_),
    .A2(_21052_),
    .A3(_07255_),
    .A4(_21055_),
    .ZN(lce_req_o[4]));
 OAI211_X2 _48849_ (.A(_21039_),
    .B(_21045_),
    .C1(_21040_),
    .C2(\icache.lru_encode [2]),
    .ZN(_21056_));
 AOI21_X4 _48850_ (.A(_21056_),
    .B1(\icache.lru_encode [2]),
    .B2(\icache.lru_encoder.lru_i [2]),
    .ZN(_21057_));
 INV_X1 _48851_ (.A(_21039_),
    .ZN(_21058_));
 OAI21_X4 _48852_ (.A(_21035_),
    .B1(_07350_),
    .B2(_07425_),
    .ZN(_21059_));
 AOI211_X2 _48853_ (.A(_21052_),
    .B(_21057_),
    .C1(_21058_),
    .C2(_21059_),
    .ZN(lce_req_o[5]));
 NAND3_X1 _48854_ (.A1(_21039_),
    .A2(_21041_),
    .A3(_21045_),
    .ZN(_21060_));
 NAND2_X2 _48855_ (.A1(_21060_),
    .A2(_21037_),
    .ZN(_21061_));
 NOR2_X4 _48856_ (.A1(_21052_),
    .A2(_21061_),
    .ZN(lce_req_o[6]));
 AOI21_X1 _48857_ (.A(_00606_),
    .B1(_00002_),
    .B2(_00604_),
    .ZN(_21062_));
 MUX2_X2 _48858_ (.A(_21062_),
    .B(\icache.lce.lce_data_cmd.miss_addr_i [0]),
    .S(_08016_),
    .Z(lce_req_o[7]));
 AOI21_X1 _48859_ (.A(_00607_),
    .B1(_00002_),
    .B2(_00604_),
    .ZN(_21063_));
 MUX2_X2 _48860_ (.A(_21063_),
    .B(\icache.lce.lce_data_cmd.miss_addr_i [1]),
    .S(_08016_),
    .Z(lce_req_o[8]));
 AOI21_X1 _48861_ (.A(_00608_),
    .B1(_00002_),
    .B2(_00604_),
    .ZN(_21064_));
 MUX2_X2 _48862_ (.A(_21064_),
    .B(\icache.lce.lce_data_cmd.miss_addr_i [2]),
    .S(_08016_),
    .Z(lce_req_o[9]));
 NAND2_X1 _48863_ (.A1(_08014_),
    .A2(\icache.lce.lce_req_inst.state_r [0]),
    .ZN(_21065_));
 NAND2_X4 _48864_ (.A1(_20994_),
    .A2(_21065_),
    .ZN(lce_req_v_o));
 AOI21_X2 _48865_ (.A(_08031_),
    .B1(_10320_),
    .B2(_10372_),
    .ZN(_21066_));
 AND4_X1 _48866_ (.A1(_00004_),
    .A2(_08029_),
    .A3(_10518_),
    .A4(_10520_),
    .ZN(_21067_));
 NOR2_X2 _48867_ (.A1(_21066_),
    .A2(_21067_),
    .ZN(_21068_));
 OAI21_X2 _48868_ (.A(_08032_),
    .B1(_10501_),
    .B2(_10502_),
    .ZN(_21069_));
 NAND3_X2 _48869_ (.A1(_08029_),
    .A2(_00004_),
    .A3(_10558_),
    .ZN(_21070_));
 AND3_X2 _48870_ (.A1(_21068_),
    .A2(_21069_),
    .A3(_21070_),
    .ZN(_21071_));
 AND3_X1 _48871_ (.A1(_10159_),
    .A2(_08032_),
    .A3(_10265_),
    .ZN(_21072_));
 AND2_X4 _48872_ (.A1(_08031_),
    .A2(_10480_),
    .ZN(_21073_));
 NOR2_X2 _48873_ (.A1(_21072_),
    .A2(_21073_),
    .ZN(_21074_));
 BUF_X4 _48874_ (.A(_21074_),
    .Z(_21075_));
 AND2_X2 _48875_ (.A1(_21071_),
    .A2(_21075_),
    .ZN(_21076_));
 NAND2_X4 _48876_ (.A1(_21076_),
    .A2(_08031_),
    .ZN(_21077_));
 BUF_X8 _48877_ (.A(_21077_),
    .Z(_21078_));
 MUX2_X1 _48878_ (.A(fe_cmd_i[1]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [132]),
    .S(_21078_),
    .Z(_06624_));
 MUX2_X1 _48879_ (.A(fe_cmd_i[7]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [138]),
    .S(_21078_),
    .Z(_06625_));
 MUX2_X1 _48880_ (.A(fe_cmd_i[8]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [139]),
    .S(_21078_),
    .Z(_06626_));
 MUX2_X1 _48881_ (.A(fe_cmd_i[9]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [140]),
    .S(_21078_),
    .Z(_06628_));
 MUX2_X1 _48882_ (.A(fe_cmd_i[10]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [141]),
    .S(_21078_),
    .Z(_06629_));
 MUX2_X1 _48883_ (.A(fe_cmd_i[11]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [142]),
    .S(_21078_),
    .Z(_06630_));
 MUX2_X1 _48884_ (.A(fe_cmd_i[12]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [143]),
    .S(_21078_),
    .Z(_06631_));
 MUX2_X1 _48885_ (.A(fe_cmd_i[13]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [144]),
    .S(_21078_),
    .Z(_06632_));
 MUX2_X1 _48886_ (.A(fe_cmd_i[14]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [145]),
    .S(_21078_),
    .Z(_06633_));
 MUX2_X1 _48887_ (.A(fe_cmd_i[15]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [146]),
    .S(_21078_),
    .Z(_06634_));
 BUF_X8 _48888_ (.A(_21077_),
    .Z(_21079_));
 MUX2_X1 _48889_ (.A(fe_cmd_i[16]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [147]),
    .S(_21079_),
    .Z(_06635_));
 MUX2_X1 _48890_ (.A(fe_cmd_i[17]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [148]),
    .S(_21079_),
    .Z(_06636_));
 MUX2_X1 _48891_ (.A(fe_cmd_i[18]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [149]),
    .S(_21079_),
    .Z(_06637_));
 MUX2_X1 _48892_ (.A(fe_cmd_i[19]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [150]),
    .S(_21079_),
    .Z(_06639_));
 MUX2_X1 _48893_ (.A(fe_cmd_i[20]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [151]),
    .S(_21079_),
    .Z(_06640_));
 MUX2_X1 _48894_ (.A(fe_cmd_i[21]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [152]),
    .S(_21079_),
    .Z(_06641_));
 MUX2_X1 _48895_ (.A(fe_cmd_i[22]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [153]),
    .S(_21079_),
    .Z(_06642_));
 MUX2_X1 _48896_ (.A(fe_cmd_i[23]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [154]),
    .S(_21079_),
    .Z(_06643_));
 MUX2_X1 _48897_ (.A(fe_cmd_i[24]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [155]),
    .S(_21079_),
    .Z(_06644_));
 MUX2_X1 _48898_ (.A(fe_cmd_i[25]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [156]),
    .S(_21079_),
    .Z(_06645_));
 MUX2_X1 _48899_ (.A(fe_cmd_i[26]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [157]),
    .S(_21077_),
    .Z(_06646_));
 MUX2_X1 _48900_ (.A(fe_cmd_i[27]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [158]),
    .S(_21077_),
    .Z(_06647_));
 MUX2_X1 _48901_ (.A(fe_cmd_i[28]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [159]),
    .S(_21077_),
    .Z(_06648_));
 MUX2_X1 _48902_ (.A(fe_cmd_i[29]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [160]),
    .S(_21077_),
    .Z(_06650_));
 MUX2_X1 _48903_ (.A(fe_cmd_i[30]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [161]),
    .S(_21077_),
    .Z(_06651_));
 MUX2_X1 _48904_ (.A(fe_cmd_i[31]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [162]),
    .S(_21077_),
    .Z(_06652_));
 MUX2_X1 _48905_ (.A(fe_cmd_i[32]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [163]),
    .S(_21077_),
    .Z(_06653_));
 MUX2_X1 _48906_ (.A(_10741_),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [164]),
    .S(_21077_),
    .Z(_06654_));
 AOI21_X4 _48907_ (.A(_21068_),
    .B1(_21069_),
    .B2(_21070_),
    .ZN(_21080_));
 AND2_X4 _48908_ (.A1(_21080_),
    .A2(_21075_),
    .ZN(_21081_));
 NAND2_X4 _48909_ (.A1(_21081_),
    .A2(_08031_),
    .ZN(_21082_));
 BUF_X8 _48910_ (.A(_21082_),
    .Z(_21083_));
 MUX2_X1 _48911_ (.A(fe_cmd_i[1]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [231]),
    .S(_21083_),
    .Z(_06718_));
 MUX2_X1 _48912_ (.A(fe_cmd_i[7]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [237]),
    .S(_21083_),
    .Z(_06719_));
 MUX2_X1 _48913_ (.A(fe_cmd_i[8]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [238]),
    .S(_21083_),
    .Z(_06720_));
 MUX2_X1 _48914_ (.A(fe_cmd_i[9]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [239]),
    .S(_21083_),
    .Z(_06721_));
 MUX2_X1 _48915_ (.A(fe_cmd_i[10]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [240]),
    .S(_21083_),
    .Z(_06723_));
 MUX2_X1 _48916_ (.A(fe_cmd_i[11]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [241]),
    .S(_21083_),
    .Z(_06724_));
 MUX2_X1 _48917_ (.A(fe_cmd_i[12]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [242]),
    .S(_21083_),
    .Z(_06725_));
 MUX2_X1 _48918_ (.A(fe_cmd_i[13]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [243]),
    .S(_21083_),
    .Z(_06726_));
 MUX2_X1 _48919_ (.A(fe_cmd_i[14]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [244]),
    .S(_21083_),
    .Z(_06727_));
 MUX2_X1 _48920_ (.A(fe_cmd_i[15]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [245]),
    .S(_21083_),
    .Z(_06728_));
 BUF_X8 _48921_ (.A(_21082_),
    .Z(_21084_));
 MUX2_X1 _48922_ (.A(fe_cmd_i[16]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [246]),
    .S(_21084_),
    .Z(_06729_));
 MUX2_X1 _48923_ (.A(fe_cmd_i[17]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [247]),
    .S(_21084_),
    .Z(_06730_));
 MUX2_X1 _48924_ (.A(fe_cmd_i[18]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [248]),
    .S(_21084_),
    .Z(_06731_));
 MUX2_X1 _48925_ (.A(fe_cmd_i[19]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [249]),
    .S(_21084_),
    .Z(_06732_));
 MUX2_X1 _48926_ (.A(fe_cmd_i[20]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [250]),
    .S(_21084_),
    .Z(_06734_));
 MUX2_X1 _48927_ (.A(fe_cmd_i[21]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [251]),
    .S(_21084_),
    .Z(_06735_));
 MUX2_X1 _48928_ (.A(fe_cmd_i[22]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [252]),
    .S(_21084_),
    .Z(_06736_));
 MUX2_X1 _48929_ (.A(fe_cmd_i[23]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [253]),
    .S(_21084_),
    .Z(_06737_));
 MUX2_X1 _48930_ (.A(fe_cmd_i[24]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [254]),
    .S(_21084_),
    .Z(_06738_));
 MUX2_X1 _48931_ (.A(fe_cmd_i[25]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [255]),
    .S(_21084_),
    .Z(_06739_));
 MUX2_X1 _48932_ (.A(fe_cmd_i[26]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [256]),
    .S(_21082_),
    .Z(_06740_));
 MUX2_X1 _48933_ (.A(fe_cmd_i[27]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [257]),
    .S(_21082_),
    .Z(_06741_));
 MUX2_X1 _48934_ (.A(fe_cmd_i[28]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [258]),
    .S(_21082_),
    .Z(_06742_));
 MUX2_X1 _48935_ (.A(fe_cmd_i[29]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [259]),
    .S(_21082_),
    .Z(_06743_));
 MUX2_X1 _48936_ (.A(fe_cmd_i[30]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [260]),
    .S(_21082_),
    .Z(_06745_));
 MUX2_X1 _48937_ (.A(fe_cmd_i[31]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [261]),
    .S(_21082_),
    .Z(_06746_));
 MUX2_X1 _48938_ (.A(fe_cmd_i[32]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [262]),
    .S(_21082_),
    .Z(_06747_));
 MUX2_X1 _48939_ (.A(_10741_),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [263]),
    .S(_21082_),
    .Z(_06748_));
 AND2_X1 _48940_ (.A1(_21069_),
    .A2(_21070_),
    .ZN(_21085_));
 INV_X1 _48941_ (.A(_21068_),
    .ZN(_21086_));
 NOR2_X2 _48942_ (.A1(_21085_),
    .A2(_21086_),
    .ZN(_21087_));
 AND2_X2 _48943_ (.A1(_21087_),
    .A2(_21074_),
    .ZN(_21088_));
 NAND2_X4 _48944_ (.A1(_21088_),
    .A2(_08031_),
    .ZN(_21089_));
 BUF_X8 _48945_ (.A(_21089_),
    .Z(_21090_));
 MUX2_X1 _48946_ (.A(fe_cmd_i[1]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [198]),
    .S(_21090_),
    .Z(_06686_));
 MUX2_X1 _48947_ (.A(fe_cmd_i[7]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [204]),
    .S(_21090_),
    .Z(_06688_));
 MUX2_X1 _48948_ (.A(fe_cmd_i[8]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [205]),
    .S(_21090_),
    .Z(_06689_));
 MUX2_X1 _48949_ (.A(fe_cmd_i[9]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [206]),
    .S(_21090_),
    .Z(_06690_));
 MUX2_X1 _48950_ (.A(fe_cmd_i[10]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [207]),
    .S(_21090_),
    .Z(_06691_));
 MUX2_X1 _48951_ (.A(fe_cmd_i[11]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [208]),
    .S(_21090_),
    .Z(_06692_));
 MUX2_X1 _48952_ (.A(fe_cmd_i[12]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [209]),
    .S(_21090_),
    .Z(_06693_));
 MUX2_X1 _48953_ (.A(fe_cmd_i[13]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [210]),
    .S(_21090_),
    .Z(_06695_));
 MUX2_X1 _48954_ (.A(fe_cmd_i[14]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [211]),
    .S(_21090_),
    .Z(_06696_));
 MUX2_X1 _48955_ (.A(fe_cmd_i[15]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [212]),
    .S(_21090_),
    .Z(_06697_));
 BUF_X4 _48956_ (.A(_21089_),
    .Z(_21091_));
 MUX2_X1 _48957_ (.A(fe_cmd_i[16]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [213]),
    .S(_21091_),
    .Z(_06698_));
 MUX2_X1 _48958_ (.A(fe_cmd_i[17]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [214]),
    .S(_21091_),
    .Z(_06699_));
 MUX2_X1 _48959_ (.A(fe_cmd_i[18]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [215]),
    .S(_21091_),
    .Z(_06700_));
 MUX2_X1 _48960_ (.A(fe_cmd_i[19]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [216]),
    .S(_21091_),
    .Z(_06701_));
 MUX2_X1 _48961_ (.A(fe_cmd_i[20]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [217]),
    .S(_21091_),
    .Z(_06702_));
 MUX2_X1 _48962_ (.A(fe_cmd_i[21]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [218]),
    .S(_21091_),
    .Z(_06703_));
 MUX2_X1 _48963_ (.A(fe_cmd_i[22]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [219]),
    .S(_21091_),
    .Z(_06704_));
 MUX2_X1 _48964_ (.A(fe_cmd_i[23]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [220]),
    .S(_21091_),
    .Z(_06706_));
 MUX2_X1 _48965_ (.A(fe_cmd_i[24]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [221]),
    .S(_21091_),
    .Z(_06707_));
 MUX2_X1 _48966_ (.A(fe_cmd_i[25]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [222]),
    .S(_21091_),
    .Z(_06708_));
 MUX2_X1 _48967_ (.A(fe_cmd_i[26]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [223]),
    .S(_21089_),
    .Z(_06709_));
 MUX2_X1 _48968_ (.A(fe_cmd_i[27]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [224]),
    .S(_21089_),
    .Z(_06710_));
 MUX2_X1 _48969_ (.A(fe_cmd_i[28]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [225]),
    .S(_21089_),
    .Z(_06711_));
 MUX2_X1 _48970_ (.A(fe_cmd_i[29]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [226]),
    .S(_21089_),
    .Z(_06712_));
 MUX2_X1 _48971_ (.A(fe_cmd_i[30]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [227]),
    .S(_21089_),
    .Z(_06713_));
 MUX2_X1 _48972_ (.A(fe_cmd_i[31]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [228]),
    .S(_21089_),
    .Z(_06714_));
 MUX2_X1 _48973_ (.A(fe_cmd_i[32]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [229]),
    .S(_21089_),
    .Z(_06715_));
 MUX2_X1 _48974_ (.A(_10741_),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [230]),
    .S(_21089_),
    .Z(_06717_));
 AND2_X1 _48975_ (.A1(_21085_),
    .A2(_21086_),
    .ZN(_21092_));
 AND2_X1 _48976_ (.A1(_21092_),
    .A2(_21074_),
    .ZN(_21093_));
 BUF_X8 _48977_ (.A(_21093_),
    .Z(_21094_));
 NAND2_X4 _48978_ (.A1(_21094_),
    .A2(_08031_),
    .ZN(_21095_));
 BUF_X8 _48979_ (.A(_21095_),
    .Z(_21096_));
 MUX2_X1 _48980_ (.A(fe_cmd_i[1]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [165]),
    .S(_21096_),
    .Z(_06655_));
 MUX2_X1 _48981_ (.A(fe_cmd_i[7]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [171]),
    .S(_21096_),
    .Z(_06657_));
 MUX2_X1 _48982_ (.A(fe_cmd_i[8]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [172]),
    .S(_21096_),
    .Z(_06658_));
 MUX2_X1 _48983_ (.A(fe_cmd_i[9]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [173]),
    .S(_21096_),
    .Z(_06659_));
 MUX2_X1 _48984_ (.A(fe_cmd_i[10]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [174]),
    .S(_21096_),
    .Z(_06660_));
 MUX2_X1 _48985_ (.A(fe_cmd_i[11]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [175]),
    .S(_21096_),
    .Z(_06661_));
 MUX2_X1 _48986_ (.A(fe_cmd_i[12]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [176]),
    .S(_21096_),
    .Z(_06662_));
 MUX2_X1 _48987_ (.A(fe_cmd_i[13]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [177]),
    .S(_21096_),
    .Z(_06663_));
 MUX2_X1 _48988_ (.A(fe_cmd_i[14]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [178]),
    .S(_21096_),
    .Z(_06664_));
 MUX2_X1 _48989_ (.A(fe_cmd_i[15]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [179]),
    .S(_21096_),
    .Z(_06665_));
 BUF_X8 _48990_ (.A(_21095_),
    .Z(_21097_));
 MUX2_X1 _48991_ (.A(fe_cmd_i[16]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [180]),
    .S(_21097_),
    .Z(_06667_));
 MUX2_X1 _48992_ (.A(fe_cmd_i[17]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [181]),
    .S(_21097_),
    .Z(_06668_));
 MUX2_X1 _48993_ (.A(fe_cmd_i[18]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [182]),
    .S(_21097_),
    .Z(_06669_));
 MUX2_X1 _48994_ (.A(fe_cmd_i[19]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [183]),
    .S(_21097_),
    .Z(_06670_));
 MUX2_X1 _48995_ (.A(fe_cmd_i[20]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [184]),
    .S(_21097_),
    .Z(_06671_));
 MUX2_X1 _48996_ (.A(fe_cmd_i[21]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [185]),
    .S(_21097_),
    .Z(_06672_));
 MUX2_X1 _48997_ (.A(fe_cmd_i[22]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [186]),
    .S(_21097_),
    .Z(_06673_));
 MUX2_X1 _48998_ (.A(fe_cmd_i[23]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [187]),
    .S(_21097_),
    .Z(_06674_));
 MUX2_X1 _48999_ (.A(fe_cmd_i[24]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [188]),
    .S(_21097_),
    .Z(_06675_));
 MUX2_X1 _49000_ (.A(fe_cmd_i[25]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [189]),
    .S(_21097_),
    .Z(_06676_));
 MUX2_X1 _49001_ (.A(fe_cmd_i[26]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [190]),
    .S(_21095_),
    .Z(_06678_));
 MUX2_X1 _49002_ (.A(fe_cmd_i[27]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [191]),
    .S(_21095_),
    .Z(_06679_));
 MUX2_X1 _49003_ (.A(fe_cmd_i[28]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [192]),
    .S(_21095_),
    .Z(_06680_));
 MUX2_X1 _49004_ (.A(fe_cmd_i[29]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [193]),
    .S(_21095_),
    .Z(_06681_));
 MUX2_X1 _49005_ (.A(fe_cmd_i[30]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [194]),
    .S(_21095_),
    .Z(_06682_));
 MUX2_X1 _49006_ (.A(fe_cmd_i[31]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [195]),
    .S(_21095_),
    .Z(_06683_));
 MUX2_X1 _49007_ (.A(fe_cmd_i[32]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [196]),
    .S(_21095_),
    .Z(_06684_));
 MUX2_X1 _49008_ (.A(_10741_),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [197]),
    .S(_21095_),
    .Z(_06685_));
 AND2_X1 _49009_ (.A1(_21080_),
    .A2(_21073_),
    .ZN(_21098_));
 BUF_X8 _49010_ (.A(_21098_),
    .Z(_21099_));
 BUF_X8 _49011_ (.A(_21099_),
    .Z(_21100_));
 MUX2_X1 _49012_ (.A(\itlb.entry_ram.z_s1r1w_mem.synth.mem [99]),
    .B(fe_cmd_i[1]),
    .S(_21100_),
    .Z(_06815_));
 MUX2_X1 _49013_ (.A(\itlb.entry_ram.z_s1r1w_mem.synth.mem [105]),
    .B(fe_cmd_i[7]),
    .S(_21100_),
    .Z(_06594_));
 MUX2_X1 _49014_ (.A(\itlb.entry_ram.z_s1r1w_mem.synth.mem [106]),
    .B(fe_cmd_i[8]),
    .S(_21100_),
    .Z(_06595_));
 MUX2_X1 _49015_ (.A(\itlb.entry_ram.z_s1r1w_mem.synth.mem [107]),
    .B(fe_cmd_i[9]),
    .S(_21100_),
    .Z(_06596_));
 MUX2_X1 _49016_ (.A(\itlb.entry_ram.z_s1r1w_mem.synth.mem [108]),
    .B(fe_cmd_i[10]),
    .S(_21100_),
    .Z(_06597_));
 MUX2_X1 _49017_ (.A(\itlb.entry_ram.z_s1r1w_mem.synth.mem [109]),
    .B(fe_cmd_i[11]),
    .S(_21100_),
    .Z(_06598_));
 MUX2_X1 _49018_ (.A(\itlb.entry_ram.z_s1r1w_mem.synth.mem [110]),
    .B(fe_cmd_i[12]),
    .S(_21100_),
    .Z(_06600_));
 MUX2_X1 _49019_ (.A(\itlb.entry_ram.z_s1r1w_mem.synth.mem [111]),
    .B(fe_cmd_i[13]),
    .S(_21100_),
    .Z(_06601_));
 MUX2_X1 _49020_ (.A(\itlb.entry_ram.z_s1r1w_mem.synth.mem [112]),
    .B(fe_cmd_i[14]),
    .S(_21100_),
    .Z(_06602_));
 MUX2_X1 _49021_ (.A(\itlb.entry_ram.z_s1r1w_mem.synth.mem [113]),
    .B(fe_cmd_i[15]),
    .S(_21100_),
    .Z(_06603_));
 BUF_X4 _49022_ (.A(_21099_),
    .Z(_21101_));
 MUX2_X1 _49023_ (.A(\itlb.entry_ram.z_s1r1w_mem.synth.mem [114]),
    .B(fe_cmd_i[16]),
    .S(_21101_),
    .Z(_06604_));
 MUX2_X1 _49024_ (.A(\itlb.entry_ram.z_s1r1w_mem.synth.mem [115]),
    .B(fe_cmd_i[17]),
    .S(_21101_),
    .Z(_06605_));
 MUX2_X1 _49025_ (.A(\itlb.entry_ram.z_s1r1w_mem.synth.mem [116]),
    .B(fe_cmd_i[18]),
    .S(_21101_),
    .Z(_06606_));
 MUX2_X1 _49026_ (.A(\itlb.entry_ram.z_s1r1w_mem.synth.mem [117]),
    .B(fe_cmd_i[19]),
    .S(_21101_),
    .Z(_06607_));
 MUX2_X1 _49027_ (.A(\itlb.entry_ram.z_s1r1w_mem.synth.mem [118]),
    .B(fe_cmd_i[20]),
    .S(_21101_),
    .Z(_06608_));
 MUX2_X1 _49028_ (.A(\itlb.entry_ram.z_s1r1w_mem.synth.mem [119]),
    .B(fe_cmd_i[21]),
    .S(_21101_),
    .Z(_06609_));
 MUX2_X1 _49029_ (.A(\itlb.entry_ram.z_s1r1w_mem.synth.mem [120]),
    .B(fe_cmd_i[22]),
    .S(_21101_),
    .Z(_06611_));
 MUX2_X1 _49030_ (.A(\itlb.entry_ram.z_s1r1w_mem.synth.mem [121]),
    .B(fe_cmd_i[23]),
    .S(_21101_),
    .Z(_06612_));
 MUX2_X1 _49031_ (.A(\itlb.entry_ram.z_s1r1w_mem.synth.mem [122]),
    .B(fe_cmd_i[24]),
    .S(_21101_),
    .Z(_06613_));
 MUX2_X1 _49032_ (.A(\itlb.entry_ram.z_s1r1w_mem.synth.mem [123]),
    .B(fe_cmd_i[25]),
    .S(_21101_),
    .Z(_06614_));
 MUX2_X1 _49033_ (.A(\itlb.entry_ram.z_s1r1w_mem.synth.mem [124]),
    .B(fe_cmd_i[26]),
    .S(_21099_),
    .Z(_06615_));
 MUX2_X1 _49034_ (.A(\itlb.entry_ram.z_s1r1w_mem.synth.mem [125]),
    .B(fe_cmd_i[27]),
    .S(_21099_),
    .Z(_06616_));
 MUX2_X1 _49035_ (.A(\itlb.entry_ram.z_s1r1w_mem.synth.mem [126]),
    .B(fe_cmd_i[28]),
    .S(_21099_),
    .Z(_06617_));
 MUX2_X1 _49036_ (.A(\itlb.entry_ram.z_s1r1w_mem.synth.mem [127]),
    .B(fe_cmd_i[29]),
    .S(_21099_),
    .Z(_06618_));
 MUX2_X1 _49037_ (.A(\itlb.entry_ram.z_s1r1w_mem.synth.mem [128]),
    .B(fe_cmd_i[30]),
    .S(_21099_),
    .Z(_06619_));
 MUX2_X1 _49038_ (.A(\itlb.entry_ram.z_s1r1w_mem.synth.mem [129]),
    .B(fe_cmd_i[31]),
    .S(_21099_),
    .Z(_06620_));
 MUX2_X1 _49039_ (.A(\itlb.entry_ram.z_s1r1w_mem.synth.mem [130]),
    .B(fe_cmd_i[32]),
    .S(_21099_),
    .Z(_06622_));
 MUX2_X1 _49040_ (.A(\itlb.entry_ram.z_s1r1w_mem.synth.mem [131]),
    .B(_10741_),
    .S(_21099_),
    .Z(_06623_));
 NAND2_X4 _49041_ (.A1(_21087_),
    .A2(_21073_),
    .ZN(_21102_));
 BUF_X8 _49042_ (.A(_21102_),
    .Z(_21103_));
 MUX2_X1 _49043_ (.A(fe_cmd_i[1]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [66]),
    .S(_21103_),
    .Z(_06784_));
 MUX2_X1 _49044_ (.A(fe_cmd_i[7]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [72]),
    .S(_21103_),
    .Z(_06786_));
 MUX2_X1 _49045_ (.A(fe_cmd_i[8]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [73]),
    .S(_21103_),
    .Z(_06787_));
 MUX2_X1 _49046_ (.A(fe_cmd_i[9]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [74]),
    .S(_21103_),
    .Z(_06788_));
 MUX2_X1 _49047_ (.A(fe_cmd_i[10]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [75]),
    .S(_21103_),
    .Z(_06789_));
 MUX2_X1 _49048_ (.A(fe_cmd_i[11]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [76]),
    .S(_21103_),
    .Z(_06790_));
 MUX2_X1 _49049_ (.A(fe_cmd_i[12]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [77]),
    .S(_21103_),
    .Z(_06791_));
 MUX2_X1 _49050_ (.A(fe_cmd_i[13]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [78]),
    .S(_21103_),
    .Z(_06792_));
 MUX2_X1 _49051_ (.A(fe_cmd_i[14]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [79]),
    .S(_21103_),
    .Z(_06793_));
 MUX2_X1 _49052_ (.A(fe_cmd_i[15]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [80]),
    .S(_21103_),
    .Z(_06795_));
 BUF_X4 _49053_ (.A(_21102_),
    .Z(_21104_));
 MUX2_X1 _49054_ (.A(fe_cmd_i[16]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [81]),
    .S(_21104_),
    .Z(_06796_));
 MUX2_X1 _49055_ (.A(fe_cmd_i[17]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [82]),
    .S(_21104_),
    .Z(_06797_));
 MUX2_X1 _49056_ (.A(fe_cmd_i[18]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [83]),
    .S(_21104_),
    .Z(_06798_));
 MUX2_X1 _49057_ (.A(fe_cmd_i[19]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [84]),
    .S(_21104_),
    .Z(_06799_));
 MUX2_X1 _49058_ (.A(fe_cmd_i[20]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [85]),
    .S(_21104_),
    .Z(_06800_));
 MUX2_X1 _49059_ (.A(fe_cmd_i[21]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [86]),
    .S(_21104_),
    .Z(_06801_));
 MUX2_X1 _49060_ (.A(fe_cmd_i[22]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [87]),
    .S(_21104_),
    .Z(_06802_));
 MUX2_X1 _49061_ (.A(fe_cmd_i[23]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [88]),
    .S(_21104_),
    .Z(_06803_));
 MUX2_X1 _49062_ (.A(fe_cmd_i[24]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [89]),
    .S(_21104_),
    .Z(_06804_));
 MUX2_X1 _49063_ (.A(fe_cmd_i[25]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [90]),
    .S(_21104_),
    .Z(_06806_));
 MUX2_X1 _49064_ (.A(fe_cmd_i[26]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [91]),
    .S(_21102_),
    .Z(_06807_));
 MUX2_X1 _49065_ (.A(fe_cmd_i[27]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [92]),
    .S(_21102_),
    .Z(_06808_));
 MUX2_X1 _49066_ (.A(fe_cmd_i[28]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [93]),
    .S(_21102_),
    .Z(_06809_));
 MUX2_X1 _49067_ (.A(fe_cmd_i[29]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [94]),
    .S(_21102_),
    .Z(_06810_));
 MUX2_X1 _49068_ (.A(fe_cmd_i[30]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [95]),
    .S(_21102_),
    .Z(_06811_));
 MUX2_X1 _49069_ (.A(fe_cmd_i[31]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [96]),
    .S(_21102_),
    .Z(_06812_));
 MUX2_X1 _49070_ (.A(fe_cmd_i[32]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [97]),
    .S(_21102_),
    .Z(_06813_));
 MUX2_X1 _49071_ (.A(_10741_),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [98]),
    .S(_21102_),
    .Z(_06814_));
 NAND2_X4 _49072_ (.A1(_21071_),
    .A2(_21073_),
    .ZN(_21105_));
 BUF_X4 _49073_ (.A(_21105_),
    .Z(_21106_));
 MUX2_X1 _49074_ (.A(fe_cmd_i[1]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [0]),
    .S(_21106_),
    .Z(_06593_));
 MUX2_X1 _49075_ (.A(fe_cmd_i[7]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [6]),
    .S(_21106_),
    .Z(_06785_));
 MUX2_X1 _49076_ (.A(fe_cmd_i[8]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [7]),
    .S(_21106_),
    .Z(_06794_));
 MUX2_X1 _49077_ (.A(fe_cmd_i[9]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [8]),
    .S(_21106_),
    .Z(_06805_));
 MUX2_X1 _49078_ (.A(fe_cmd_i[10]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [9]),
    .S(_21106_),
    .Z(_06816_));
 MUX2_X1 _49079_ (.A(fe_cmd_i[11]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [10]),
    .S(_21106_),
    .Z(_06599_));
 MUX2_X1 _49080_ (.A(fe_cmd_i[12]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [11]),
    .S(_21106_),
    .Z(_06610_));
 MUX2_X1 _49081_ (.A(fe_cmd_i[13]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [12]),
    .S(_21106_),
    .Z(_06621_));
 MUX2_X1 _49082_ (.A(fe_cmd_i[14]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [13]),
    .S(_21106_),
    .Z(_06627_));
 MUX2_X1 _49083_ (.A(fe_cmd_i[15]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [14]),
    .S(_21106_),
    .Z(_06638_));
 BUF_X4 _49084_ (.A(_21105_),
    .Z(_21107_));
 MUX2_X1 _49085_ (.A(fe_cmd_i[16]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [15]),
    .S(_21107_),
    .Z(_06649_));
 MUX2_X1 _49086_ (.A(fe_cmd_i[17]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [16]),
    .S(_21107_),
    .Z(_06656_));
 MUX2_X1 _49087_ (.A(fe_cmd_i[18]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [17]),
    .S(_21107_),
    .Z(_06666_));
 MUX2_X1 _49088_ (.A(fe_cmd_i[19]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [18]),
    .S(_21107_),
    .Z(_06677_));
 MUX2_X1 _49089_ (.A(fe_cmd_i[20]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [19]),
    .S(_21107_),
    .Z(_06687_));
 MUX2_X1 _49090_ (.A(fe_cmd_i[21]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [20]),
    .S(_21107_),
    .Z(_06694_));
 MUX2_X1 _49091_ (.A(fe_cmd_i[22]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [21]),
    .S(_21107_),
    .Z(_06705_));
 MUX2_X1 _49092_ (.A(fe_cmd_i[23]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [22]),
    .S(_21107_),
    .Z(_06716_));
 MUX2_X1 _49093_ (.A(fe_cmd_i[24]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [23]),
    .S(_21107_),
    .Z(_06722_));
 MUX2_X1 _49094_ (.A(fe_cmd_i[25]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [24]),
    .S(_21107_),
    .Z(_06733_));
 MUX2_X1 _49095_ (.A(fe_cmd_i[26]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [25]),
    .S(_21105_),
    .Z(_06744_));
 MUX2_X1 _49096_ (.A(fe_cmd_i[27]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [26]),
    .S(_21105_),
    .Z(_06749_));
 MUX2_X1 _49097_ (.A(fe_cmd_i[28]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [27]),
    .S(_21105_),
    .Z(_06750_));
 MUX2_X1 _49098_ (.A(fe_cmd_i[29]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [28]),
    .S(_21105_),
    .Z(_06751_));
 MUX2_X1 _49099_ (.A(fe_cmd_i[30]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [29]),
    .S(_21105_),
    .Z(_06752_));
 MUX2_X1 _49100_ (.A(fe_cmd_i[31]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [30]),
    .S(_21105_),
    .Z(_06753_));
 MUX2_X1 _49101_ (.A(fe_cmd_i[32]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [31]),
    .S(_21105_),
    .Z(_06754_));
 MUX2_X1 _49102_ (.A(_10741_),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [32]),
    .S(_21105_),
    .Z(_06755_));
 NAND2_X4 _49103_ (.A1(_21092_),
    .A2(_21073_),
    .ZN(_21108_));
 BUF_X8 _49104_ (.A(_21108_),
    .Z(_21109_));
 MUX2_X1 _49105_ (.A(fe_cmd_i[1]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [33]),
    .S(_21109_),
    .Z(_06756_));
 MUX2_X1 _49106_ (.A(fe_cmd_i[7]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [39]),
    .S(_21109_),
    .Z(_06757_));
 MUX2_X1 _49107_ (.A(fe_cmd_i[8]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [40]),
    .S(_21109_),
    .Z(_06758_));
 MUX2_X1 _49108_ (.A(fe_cmd_i[9]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [41]),
    .S(_21109_),
    .Z(_06759_));
 MUX2_X1 _49109_ (.A(fe_cmd_i[10]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [42]),
    .S(_21109_),
    .Z(_06760_));
 MUX2_X1 _49110_ (.A(fe_cmd_i[11]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [43]),
    .S(_21109_),
    .Z(_06761_));
 MUX2_X1 _49111_ (.A(fe_cmd_i[12]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [44]),
    .S(_21109_),
    .Z(_06762_));
 MUX2_X1 _49112_ (.A(fe_cmd_i[13]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [45]),
    .S(_21109_),
    .Z(_06763_));
 MUX2_X1 _49113_ (.A(fe_cmd_i[14]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [46]),
    .S(_21109_),
    .Z(_06764_));
 MUX2_X1 _49114_ (.A(fe_cmd_i[15]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [47]),
    .S(_21109_),
    .Z(_06765_));
 BUF_X4 _49115_ (.A(_21108_),
    .Z(_21110_));
 MUX2_X1 _49116_ (.A(fe_cmd_i[16]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [48]),
    .S(_21110_),
    .Z(_06766_));
 MUX2_X1 _49117_ (.A(fe_cmd_i[17]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [49]),
    .S(_21110_),
    .Z(_06767_));
 MUX2_X1 _49118_ (.A(fe_cmd_i[18]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [50]),
    .S(_21110_),
    .Z(_06768_));
 MUX2_X1 _49119_ (.A(fe_cmd_i[19]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [51]),
    .S(_21110_),
    .Z(_06769_));
 MUX2_X1 _49120_ (.A(fe_cmd_i[20]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [52]),
    .S(_21110_),
    .Z(_06770_));
 MUX2_X1 _49121_ (.A(fe_cmd_i[21]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [53]),
    .S(_21110_),
    .Z(_06771_));
 MUX2_X1 _49122_ (.A(fe_cmd_i[22]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [54]),
    .S(_21110_),
    .Z(_06772_));
 MUX2_X1 _49123_ (.A(fe_cmd_i[23]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [55]),
    .S(_21110_),
    .Z(_06773_));
 MUX2_X1 _49124_ (.A(fe_cmd_i[24]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [56]),
    .S(_21110_),
    .Z(_06774_));
 MUX2_X1 _49125_ (.A(fe_cmd_i[25]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [57]),
    .S(_21110_),
    .Z(_06775_));
 MUX2_X1 _49126_ (.A(fe_cmd_i[26]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [58]),
    .S(_21108_),
    .Z(_06776_));
 MUX2_X1 _49127_ (.A(fe_cmd_i[27]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [59]),
    .S(_21108_),
    .Z(_06777_));
 MUX2_X1 _49128_ (.A(fe_cmd_i[28]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [60]),
    .S(_21108_),
    .Z(_06778_));
 MUX2_X1 _49129_ (.A(fe_cmd_i[29]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [61]),
    .S(_21108_),
    .Z(_06779_));
 MUX2_X1 _49130_ (.A(fe_cmd_i[30]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [62]),
    .S(_21108_),
    .Z(_06780_));
 MUX2_X1 _49131_ (.A(fe_cmd_i[31]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [63]),
    .S(_21108_),
    .Z(_06781_));
 MUX2_X1 _49132_ (.A(fe_cmd_i[32]),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [64]),
    .S(_21108_),
    .Z(_06782_));
 MUX2_X1 _49133_ (.A(_10741_),
    .B(\itlb.entry_ram.z_s1r1w_mem.synth.mem [65]),
    .S(_21108_),
    .Z(_06783_));
 INV_X1 _49134_ (.A(_21074_),
    .ZN(_21111_));
 AND2_X1 _49135_ (.A1(_21092_),
    .A2(_21111_),
    .ZN(_21112_));
 BUF_X8 _49136_ (.A(_21112_),
    .Z(_21113_));
 BUF_X8 _49137_ (.A(_21113_),
    .Z(_21114_));
 AND2_X1 _49138_ (.A1(_21080_),
    .A2(_21111_),
    .ZN(_21115_));
 BUF_X8 _49139_ (.A(_21115_),
    .Z(_21116_));
 BUF_X8 _49140_ (.A(_21116_),
    .Z(_21117_));
 AOI22_X1 _49141_ (.A1(_21114_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [33]),
    .B1(\itlb.entry_ram.z_s1r1w_mem.synth.mem [99]),
    .B2(_21117_),
    .ZN(_21118_));
 AND2_X1 _49142_ (.A1(_21087_),
    .A2(_21111_),
    .ZN(_21119_));
 BUF_X8 _49143_ (.A(_21119_),
    .Z(_21120_));
 BUF_X8 _49144_ (.A(_21120_),
    .Z(_21121_));
 AND2_X1 _49145_ (.A1(_21071_),
    .A2(_21111_),
    .ZN(_21122_));
 BUF_X8 _49146_ (.A(_21122_),
    .Z(_21123_));
 BUF_X8 _49147_ (.A(_21123_),
    .Z(_21124_));
 AOI22_X1 _49148_ (.A1(_21121_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [66]),
    .B1(_21124_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [0]),
    .ZN(_21125_));
 AND3_X1 _49149_ (.A1(_21080_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [231]),
    .A3(_21075_),
    .ZN(_21126_));
 BUF_X16 _49150_ (.A(_21088_),
    .Z(_21127_));
 BUF_X8 _49151_ (.A(_21127_),
    .Z(_21128_));
 AOI21_X1 _49152_ (.A(_21126_),
    .B1(_21128_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [198]),
    .ZN(_21129_));
 AND4_X1 _49153_ (.A1(\itlb.entry_ram.z_s1r1w_mem.synth.mem [165]),
    .A2(_21085_),
    .A3(_21086_),
    .A4(_21075_),
    .ZN(_21130_));
 BUF_X8 _49154_ (.A(_21076_),
    .Z(_21131_));
 BUF_X8 _49155_ (.A(_21131_),
    .Z(_21132_));
 AOI21_X1 _49156_ (.A(_21130_),
    .B1(_21132_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [132]),
    .ZN(_21133_));
 NAND4_X1 _49157_ (.A1(_21118_),
    .A2(_21125_),
    .A3(_21129_),
    .A4(_21133_),
    .ZN(\itlb.entry_ram.z_s1r1w_data_lo [0]));
 BUF_X8 _49158_ (.A(_21094_),
    .Z(_21134_));
 BUF_X8 _49159_ (.A(_21081_),
    .Z(_21135_));
 AOI22_X2 _49160_ (.A1(_21134_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [171]),
    .B1(\itlb.entry_ram.z_s1r1w_mem.synth.mem [237]),
    .B2(_21135_),
    .ZN(_21136_));
 AOI22_X2 _49161_ (.A1(_21114_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [39]),
    .B1(\itlb.entry_ram.z_s1r1w_mem.synth.mem [105]),
    .B2(_21117_),
    .ZN(_21137_));
 AOI22_X2 _49162_ (.A1(_21121_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [72]),
    .B1(_21131_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [138]),
    .ZN(_21138_));
 AOI22_X2 _49163_ (.A1(_21127_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [204]),
    .B1(_21124_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [6]),
    .ZN(_21139_));
 NAND4_X2 _49164_ (.A1(_21136_),
    .A2(_21137_),
    .A3(_21138_),
    .A4(_21139_),
    .ZN(\itlb.entry_ram.z_s1r1w_data_lo [6]));
 AOI22_X1 _49165_ (.A1(_21134_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [172]),
    .B1(\itlb.entry_ram.z_s1r1w_mem.synth.mem [238]),
    .B2(_21135_),
    .ZN(_21140_));
 AOI22_X1 _49166_ (.A1(_21114_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [40]),
    .B1(\itlb.entry_ram.z_s1r1w_mem.synth.mem [106]),
    .B2(_21117_),
    .ZN(_21141_));
 AOI22_X1 _49167_ (.A1(_21121_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [73]),
    .B1(_21131_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [139]),
    .ZN(_21142_));
 AOI22_X2 _49168_ (.A1(_21127_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [205]),
    .B1(_21124_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [7]),
    .ZN(_21143_));
 NAND4_X1 _49169_ (.A1(_21140_),
    .A2(_21141_),
    .A3(_21142_),
    .A4(_21143_),
    .ZN(\itlb.entry_ram.z_s1r1w_data_lo [7]));
 AOI22_X1 _49170_ (.A1(_21134_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [173]),
    .B1(_21132_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [140]),
    .ZN(_21144_));
 AOI22_X2 _49171_ (.A1(_21114_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [41]),
    .B1(\itlb.entry_ram.z_s1r1w_mem.synth.mem [107]),
    .B2(_21117_),
    .ZN(_21145_));
 AOI22_X2 _49172_ (.A1(_21128_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [206]),
    .B1(_21135_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [239]),
    .ZN(_21146_));
 BUF_X8 _49173_ (.A(_21120_),
    .Z(_21147_));
 AOI22_X2 _49174_ (.A1(_21147_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [74]),
    .B1(_21124_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [8]),
    .ZN(_21148_));
 NAND4_X2 _49175_ (.A1(_21144_),
    .A2(_21145_),
    .A3(_21146_),
    .A4(_21148_),
    .ZN(\itlb.entry_ram.z_s1r1w_data_lo [8]));
 AOI22_X2 _49176_ (.A1(_21114_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [42]),
    .B1(\itlb.entry_ram.z_s1r1w_mem.synth.mem [108]),
    .B2(_21117_),
    .ZN(_21149_));
 AOI22_X1 _49177_ (.A1(_21128_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [207]),
    .B1(_21135_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [240]),
    .ZN(_21150_));
 AOI22_X2 _49178_ (.A1(_21121_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [75]),
    .B1(_21124_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [9]),
    .ZN(_21151_));
 AND4_X1 _49179_ (.A1(\itlb.entry_ram.z_s1r1w_mem.synth.mem [174]),
    .A2(_21085_),
    .A3(_21086_),
    .A4(_21075_),
    .ZN(_21152_));
 AOI21_X1 _49180_ (.A(_21152_),
    .B1(_21132_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [141]),
    .ZN(_21153_));
 NAND4_X1 _49181_ (.A1(_21149_),
    .A2(_21150_),
    .A3(_21151_),
    .A4(_21153_),
    .ZN(\itlb.entry_ram.z_s1r1w_data_lo [9]));
 AOI22_X1 _49182_ (.A1(_21134_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [175]),
    .B1(_21132_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [142]),
    .ZN(_21154_));
 AOI22_X1 _49183_ (.A1(_21114_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [43]),
    .B1(\itlb.entry_ram.z_s1r1w_mem.synth.mem [109]),
    .B2(_21117_),
    .ZN(_21155_));
 AOI22_X2 _49184_ (.A1(_21128_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [208]),
    .B1(_21135_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [241]),
    .ZN(_21156_));
 BUF_X8 _49185_ (.A(_21123_),
    .Z(_21157_));
 AOI22_X2 _49186_ (.A1(_21147_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [76]),
    .B1(_21157_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [10]),
    .ZN(_21158_));
 NAND4_X1 _49187_ (.A1(_21154_),
    .A2(_21155_),
    .A3(_21156_),
    .A4(_21158_),
    .ZN(\itlb.entry_ram.z_s1r1w_data_lo [10]));
 AOI22_X1 _49188_ (.A1(_21134_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [176]),
    .B1(_21132_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [143]),
    .ZN(_21159_));
 AOI22_X1 _49189_ (.A1(_21114_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [44]),
    .B1(\itlb.entry_ram.z_s1r1w_mem.synth.mem [110]),
    .B2(_21117_),
    .ZN(_21160_));
 AOI22_X1 _49190_ (.A1(_21128_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [209]),
    .B1(_21135_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [242]),
    .ZN(_21161_));
 AOI22_X2 _49191_ (.A1(_21147_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [77]),
    .B1(_21157_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [11]),
    .ZN(_21162_));
 NAND4_X1 _49192_ (.A1(_21159_),
    .A2(_21160_),
    .A3(_21161_),
    .A4(_21162_),
    .ZN(\itlb.entry_ram.z_s1r1w_data_lo [11]));
 AOI22_X1 _49193_ (.A1(_21134_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [177]),
    .B1(_21132_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [144]),
    .ZN(_21163_));
 AOI22_X2 _49194_ (.A1(_21114_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [45]),
    .B1(\itlb.entry_ram.z_s1r1w_mem.synth.mem [111]),
    .B2(_21117_),
    .ZN(_21164_));
 BUF_X8 _49195_ (.A(_21127_),
    .Z(_21165_));
 BUF_X8 _49196_ (.A(_21081_),
    .Z(_21166_));
 AOI22_X2 _49197_ (.A1(_21165_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [210]),
    .B1(_21166_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [243]),
    .ZN(_21167_));
 AOI22_X2 _49198_ (.A1(_21147_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [78]),
    .B1(_21157_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [12]),
    .ZN(_21168_));
 NAND4_X2 _49199_ (.A1(_21163_),
    .A2(_21164_),
    .A3(_21167_),
    .A4(_21168_),
    .ZN(\itlb.entry_ram.z_s1r1w_data_lo [12]));
 AOI22_X1 _49200_ (.A1(_21134_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [178]),
    .B1(\itlb.entry_ram.z_s1r1w_mem.synth.mem [244]),
    .B2(_21135_),
    .ZN(_21169_));
 AOI22_X2 _49201_ (.A1(_21114_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [46]),
    .B1(\itlb.entry_ram.z_s1r1w_mem.synth.mem [112]),
    .B2(_21117_),
    .ZN(_21170_));
 AOI22_X1 _49202_ (.A1(_21121_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [79]),
    .B1(_21131_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [145]),
    .ZN(_21171_));
 AOI22_X2 _49203_ (.A1(_21127_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [211]),
    .B1(_21157_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [13]),
    .ZN(_21172_));
 NAND4_X1 _49204_ (.A1(_21169_),
    .A2(_21170_),
    .A3(_21171_),
    .A4(_21172_),
    .ZN(\itlb.entry_ram.z_s1r1w_data_lo [13]));
 AOI22_X1 _49205_ (.A1(_21134_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [179]),
    .B1(_21132_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [146]),
    .ZN(_21173_));
 AOI22_X1 _49206_ (.A1(_21114_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [47]),
    .B1(\itlb.entry_ram.z_s1r1w_mem.synth.mem [113]),
    .B2(_21117_),
    .ZN(_21174_));
 AOI22_X4 _49207_ (.A1(_21165_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [212]),
    .B1(_21166_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [245]),
    .ZN(_21175_));
 AOI22_X1 _49208_ (.A1(_21147_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [80]),
    .B1(_21157_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [14]),
    .ZN(_21176_));
 NAND4_X1 _49209_ (.A1(_21173_),
    .A2(_21174_),
    .A3(_21175_),
    .A4(_21176_),
    .ZN(\itlb.entry_ram.z_s1r1w_data_lo [14]));
 AOI22_X1 _49210_ (.A1(_21134_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [180]),
    .B1(\itlb.entry_ram.z_s1r1w_mem.synth.mem [246]),
    .B2(_21135_),
    .ZN(_21177_));
 BUF_X8 _49211_ (.A(_21113_),
    .Z(_21178_));
 BUF_X8 _49212_ (.A(_21116_),
    .Z(_21179_));
 AOI22_X4 _49213_ (.A1(_21178_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [48]),
    .B1(\itlb.entry_ram.z_s1r1w_mem.synth.mem [114]),
    .B2(_21179_),
    .ZN(_21180_));
 AOI22_X2 _49214_ (.A1(_21121_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [81]),
    .B1(_21131_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [147]),
    .ZN(_21181_));
 AOI22_X1 _49215_ (.A1(_21127_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [213]),
    .B1(_21157_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [15]),
    .ZN(_21182_));
 NAND4_X1 _49216_ (.A1(_21177_),
    .A2(_21180_),
    .A3(_21181_),
    .A4(_21182_),
    .ZN(\itlb.entry_ram.z_s1r1w_data_lo [15]));
 AOI22_X2 _49217_ (.A1(_21134_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [181]),
    .B1(_21132_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [148]),
    .ZN(_21183_));
 AOI22_X4 _49218_ (.A1(_21178_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [49]),
    .B1(\itlb.entry_ram.z_s1r1w_mem.synth.mem [115]),
    .B2(_21179_),
    .ZN(_21184_));
 AOI22_X1 _49219_ (.A1(_21121_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [82]),
    .B1(_21124_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [16]),
    .ZN(_21185_));
 AND3_X1 _49220_ (.A1(_21080_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [247]),
    .A3(_21075_),
    .ZN(_21186_));
 AOI21_X1 _49221_ (.A(_21186_),
    .B1(_21128_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [214]),
    .ZN(_21187_));
 NAND4_X1 _49222_ (.A1(_21183_),
    .A2(_21184_),
    .A3(_21185_),
    .A4(_21187_),
    .ZN(\itlb.entry_ram.z_s1r1w_data_lo [16]));
 BUF_X8 _49223_ (.A(_21094_),
    .Z(_21188_));
 BUF_X8 _49224_ (.A(_21131_),
    .Z(_21189_));
 AOI22_X1 _49225_ (.A1(_21188_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [182]),
    .B1(_21189_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [149]),
    .ZN(_21190_));
 AOI22_X2 _49226_ (.A1(_21178_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [50]),
    .B1(\itlb.entry_ram.z_s1r1w_mem.synth.mem [116]),
    .B2(_21179_),
    .ZN(_21191_));
 AOI22_X1 _49227_ (.A1(_21165_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [215]),
    .B1(_21166_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [248]),
    .ZN(_21192_));
 AOI22_X2 _49228_ (.A1(_21147_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [83]),
    .B1(_21157_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [17]),
    .ZN(_21193_));
 NAND4_X1 _49229_ (.A1(_21190_),
    .A2(_21191_),
    .A3(_21192_),
    .A4(_21193_),
    .ZN(\itlb.entry_ram.z_s1r1w_data_lo [17]));
 AOI22_X2 _49230_ (.A1(_21188_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [183]),
    .B1(_21189_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [150]),
    .ZN(_21194_));
 AOI22_X4 _49231_ (.A1(_21178_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [51]),
    .B1(\itlb.entry_ram.z_s1r1w_mem.synth.mem [117]),
    .B2(_21179_),
    .ZN(_21195_));
 AOI22_X1 _49232_ (.A1(_21165_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [216]),
    .B1(_21166_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [249]),
    .ZN(_21196_));
 AOI22_X1 _49233_ (.A1(_21147_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [84]),
    .B1(_21157_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [18]),
    .ZN(_21197_));
 NAND4_X1 _49234_ (.A1(_21194_),
    .A2(_21195_),
    .A3(_21196_),
    .A4(_21197_),
    .ZN(\itlb.entry_ram.z_s1r1w_data_lo [18]));
 AOI22_X2 _49235_ (.A1(_21188_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [184]),
    .B1(_21189_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [151]),
    .ZN(_21198_));
 AOI22_X4 _49236_ (.A1(_21178_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [52]),
    .B1(\itlb.entry_ram.z_s1r1w_mem.synth.mem [118]),
    .B2(_21179_),
    .ZN(_21199_));
 AOI22_X1 _49237_ (.A1(_21165_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [217]),
    .B1(_21166_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [250]),
    .ZN(_21200_));
 AOI22_X2 _49238_ (.A1(_21120_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [85]),
    .B1(_21157_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [19]),
    .ZN(_21201_));
 NAND4_X2 _49239_ (.A1(_21198_),
    .A2(_21199_),
    .A3(_21200_),
    .A4(_21201_),
    .ZN(\itlb.entry_ram.z_s1r1w_data_lo [19]));
 AOI22_X1 _49240_ (.A1(_21188_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [185]),
    .B1(_21189_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [152]),
    .ZN(_21202_));
 AOI22_X2 _49241_ (.A1(_21178_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [53]),
    .B1(\itlb.entry_ram.z_s1r1w_mem.synth.mem [119]),
    .B2(_21179_),
    .ZN(_21203_));
 AOI22_X1 _49242_ (.A1(_21165_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [218]),
    .B1(_21166_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [251]),
    .ZN(_21204_));
 AOI22_X2 _49243_ (.A1(_21120_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [86]),
    .B1(_21157_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [20]),
    .ZN(_21205_));
 NAND4_X1 _49244_ (.A1(_21202_),
    .A2(_21203_),
    .A3(_21204_),
    .A4(_21205_),
    .ZN(\itlb.entry_ram.z_s1r1w_data_lo [20]));
 AOI22_X1 _49245_ (.A1(_21188_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [186]),
    .B1(_21189_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [153]),
    .ZN(_21206_));
 AOI22_X2 _49246_ (.A1(_21178_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [54]),
    .B1(\itlb.entry_ram.z_s1r1w_mem.synth.mem [120]),
    .B2(_21179_),
    .ZN(_21207_));
 AOI22_X1 _49247_ (.A1(_21165_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [219]),
    .B1(_21166_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [252]),
    .ZN(_21208_));
 AOI22_X2 _49248_ (.A1(_21120_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [87]),
    .B1(_21123_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [21]),
    .ZN(_21209_));
 NAND4_X1 _49249_ (.A1(_21206_),
    .A2(_21207_),
    .A3(_21208_),
    .A4(_21209_),
    .ZN(\itlb.entry_ram.z_s1r1w_data_lo [21]));
 AOI22_X1 _49250_ (.A1(_21188_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [187]),
    .B1(_21189_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [154]),
    .ZN(_21210_));
 AOI22_X2 _49251_ (.A1(_21178_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [55]),
    .B1(\itlb.entry_ram.z_s1r1w_mem.synth.mem [121]),
    .B2(_21179_),
    .ZN(_21211_));
 AOI22_X2 _49252_ (.A1(_21121_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [88]),
    .B1(_21124_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [22]),
    .ZN(_21212_));
 AND3_X1 _49253_ (.A1(_21080_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [253]),
    .A3(_21075_),
    .ZN(_21213_));
 AOI21_X1 _49254_ (.A(_21213_),
    .B1(_21128_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [220]),
    .ZN(_21214_));
 NAND4_X1 _49255_ (.A1(_21210_),
    .A2(_21211_),
    .A3(_21212_),
    .A4(_21214_),
    .ZN(\itlb.entry_ram.z_s1r1w_data_lo [22]));
 AOI22_X2 _49256_ (.A1(_21188_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [188]),
    .B1(\itlb.entry_ram.z_s1r1w_mem.synth.mem [254]),
    .B2(_21135_),
    .ZN(_21215_));
 AOI22_X4 _49257_ (.A1(_21178_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [56]),
    .B1(\itlb.entry_ram.z_s1r1w_mem.synth.mem [122]),
    .B2(_21179_),
    .ZN(_21216_));
 AOI22_X2 _49258_ (.A1(_21121_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [89]),
    .B1(_21131_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [155]),
    .ZN(_21217_));
 AOI22_X2 _49259_ (.A1(_21127_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [221]),
    .B1(_21123_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [23]),
    .ZN(_21218_));
 NAND4_X2 _49260_ (.A1(_21215_),
    .A2(_21216_),
    .A3(_21217_),
    .A4(_21218_),
    .ZN(\itlb.entry_ram.z_s1r1w_data_lo [23]));
 AOI22_X2 _49261_ (.A1(_21188_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [189]),
    .B1(_21189_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [156]),
    .ZN(_21219_));
 AOI22_X4 _49262_ (.A1(_21178_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [57]),
    .B1(\itlb.entry_ram.z_s1r1w_mem.synth.mem [123]),
    .B2(_21179_),
    .ZN(_21220_));
 AOI22_X2 _49263_ (.A1(_21121_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [90]),
    .B1(_21124_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [24]),
    .ZN(_21221_));
 AND3_X1 _49264_ (.A1(_21080_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [255]),
    .A3(_21075_),
    .ZN(_21222_));
 AOI21_X2 _49265_ (.A(_21222_),
    .B1(_21128_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [222]),
    .ZN(_21223_));
 NAND4_X2 _49266_ (.A1(_21219_),
    .A2(_21220_),
    .A3(_21221_),
    .A4(_21223_),
    .ZN(\itlb.entry_ram.z_s1r1w_data_lo [24]));
 AOI22_X1 _49267_ (.A1(_21188_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [190]),
    .B1(_21189_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [157]),
    .ZN(_21224_));
 AOI22_X2 _49268_ (.A1(_21113_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [58]),
    .B1(\itlb.entry_ram.z_s1r1w_mem.synth.mem [124]),
    .B2(_21116_),
    .ZN(_21225_));
 AOI22_X1 _49269_ (.A1(_21147_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [91]),
    .B1(_21124_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [25]),
    .ZN(_21226_));
 AND3_X1 _49270_ (.A1(_21080_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [256]),
    .A3(_21075_),
    .ZN(_21227_));
 AOI21_X1 _49271_ (.A(_21227_),
    .B1(_21128_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [223]),
    .ZN(_21228_));
 NAND4_X1 _49272_ (.A1(_21224_),
    .A2(_21225_),
    .A3(_21226_),
    .A4(_21228_),
    .ZN(\itlb.entry_ram.z_s1r1w_data_lo [25]));
 AOI22_X2 _49273_ (.A1(_21188_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [191]),
    .B1(_21189_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [158]),
    .ZN(_21229_));
 AOI22_X4 _49274_ (.A1(_21113_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [59]),
    .B1(\itlb.entry_ram.z_s1r1w_mem.synth.mem [125]),
    .B2(_21116_),
    .ZN(_21230_));
 AOI22_X2 _49275_ (.A1(_21165_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [224]),
    .B1(_21166_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [257]),
    .ZN(_21231_));
 AOI22_X2 _49276_ (.A1(_21120_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [92]),
    .B1(_21123_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [26]),
    .ZN(_21232_));
 NAND4_X2 _49277_ (.A1(_21229_),
    .A2(_21230_),
    .A3(_21231_),
    .A4(_21232_),
    .ZN(\itlb.entry_ram.z_s1r1w_data_lo [26]));
 AOI22_X2 _49278_ (.A1(_21094_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [192]),
    .B1(_21189_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [159]),
    .ZN(_21233_));
 AOI22_X2 _49279_ (.A1(_21113_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [60]),
    .B1(\itlb.entry_ram.z_s1r1w_mem.synth.mem [126]),
    .B2(_21116_),
    .ZN(_21234_));
 AOI22_X1 _49280_ (.A1(_21165_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [225]),
    .B1(_21166_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [258]),
    .ZN(_21235_));
 AOI22_X1 _49281_ (.A1(_21120_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [93]),
    .B1(_21123_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [27]),
    .ZN(_21236_));
 NAND4_X1 _49282_ (.A1(_21233_),
    .A2(_21234_),
    .A3(_21235_),
    .A4(_21236_),
    .ZN(\itlb.entry_ram.z_s1r1w_data_lo [27]));
 AOI22_X2 _49283_ (.A1(_21094_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [193]),
    .B1(\itlb.entry_ram.z_s1r1w_mem.synth.mem [259]),
    .B2(_21135_),
    .ZN(_21237_));
 AOI22_X2 _49284_ (.A1(_21113_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [61]),
    .B1(\itlb.entry_ram.z_s1r1w_mem.synth.mem [127]),
    .B2(_21116_),
    .ZN(_21238_));
 AOI22_X2 _49285_ (.A1(_21147_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [94]),
    .B1(_21131_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [160]),
    .ZN(_21239_));
 AOI22_X4 _49286_ (.A1(_21127_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [226]),
    .B1(_21123_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [28]),
    .ZN(_21240_));
 NAND4_X4 _49287_ (.A1(_21237_),
    .A2(_21238_),
    .A3(_21239_),
    .A4(_21240_),
    .ZN(\itlb.entry_ram.z_s1r1w_data_lo [28]));
 AOI22_X1 _49288_ (.A1(_21094_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [194]),
    .B1(_21120_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [95]),
    .ZN(_21241_));
 AOI22_X1 _49289_ (.A1(_21113_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [62]),
    .B1(\itlb.entry_ram.z_s1r1w_mem.synth.mem [128]),
    .B2(_21116_),
    .ZN(_21242_));
 AOI22_X1 _49290_ (.A1(\itlb.entry_ram.z_s1r1w_mem.synth.mem [161]),
    .A2(_21132_),
    .B1(_21166_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [260]),
    .ZN(_21243_));
 AOI22_X1 _49291_ (.A1(_21127_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [227]),
    .B1(_21123_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [29]),
    .ZN(_21244_));
 NAND4_X1 _49292_ (.A1(_21241_),
    .A2(_21242_),
    .A3(_21243_),
    .A4(_21244_),
    .ZN(\itlb.entry_ram.z_s1r1w_data_lo [29]));
 AOI22_X2 _49293_ (.A1(_21094_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [195]),
    .B1(_21131_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [162]),
    .ZN(_21245_));
 AOI22_X1 _49294_ (.A1(_21113_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [63]),
    .B1(\itlb.entry_ram.z_s1r1w_mem.synth.mem [129]),
    .B2(_21116_),
    .ZN(_21246_));
 AOI22_X1 _49295_ (.A1(_21165_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [228]),
    .B1(_21081_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [261]),
    .ZN(_21247_));
 AOI22_X2 _49296_ (.A1(_21120_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [96]),
    .B1(_21123_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [30]),
    .ZN(_21248_));
 NAND4_X1 _49297_ (.A1(_21245_),
    .A2(_21246_),
    .A3(_21247_),
    .A4(_21248_),
    .ZN(\itlb.entry_ram.z_s1r1w_data_lo [30]));
 AOI22_X1 _49298_ (.A1(_21094_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [196]),
    .B1(_21120_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [97]),
    .ZN(_21249_));
 AOI22_X4 _49299_ (.A1(_21113_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [64]),
    .B1(\itlb.entry_ram.z_s1r1w_mem.synth.mem [130]),
    .B2(_21116_),
    .ZN(_21250_));
 AOI22_X1 _49300_ (.A1(\itlb.entry_ram.z_s1r1w_mem.synth.mem [163]),
    .A2(_21132_),
    .B1(_21081_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [262]),
    .ZN(_21251_));
 AOI22_X2 _49301_ (.A1(_21127_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [229]),
    .B1(_21123_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [31]),
    .ZN(_21252_));
 NAND4_X1 _49302_ (.A1(_21249_),
    .A2(_21250_),
    .A3(_21251_),
    .A4(_21252_),
    .ZN(\itlb.entry_ram.z_s1r1w_data_lo [31]));
 AOI22_X1 _49303_ (.A1(_21094_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [197]),
    .B1(_21131_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [164]),
    .ZN(_21253_));
 AOI22_X1 _49304_ (.A1(_21113_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [65]),
    .B1(\itlb.entry_ram.z_s1r1w_mem.synth.mem [131]),
    .B2(_21116_),
    .ZN(_21254_));
 AOI22_X1 _49305_ (.A1(_21147_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [98]),
    .B1(_21124_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [32]),
    .ZN(_21255_));
 AND3_X1 _49306_ (.A1(_21080_),
    .A2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [263]),
    .A3(_21075_),
    .ZN(_21256_));
 AOI21_X1 _49307_ (.A(_21256_),
    .B1(_21128_),
    .B2(\itlb.entry_ram.z_s1r1w_mem.synth.mem [230]),
    .ZN(_21257_));
 NAND4_X1 _49308_ (.A1(_21253_),
    .A2(_21254_),
    .A3(_21255_),
    .A4(_21257_),
    .ZN(\itlb.entry_ram.z_s1r1w_data_lo [32]));
 INV_X1 _49309_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.full_r ),
    .ZN(_21258_));
 AND2_X2 _49310_ (.A1(_21258_),
    .A2(lce_cmd_v_i),
    .ZN(_21259_));
 AND2_X1 _49311_ (.A1(_21259_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.w_addr_i ),
    .ZN(_21260_));
 BUF_X4 _49312_ (.A(_21260_),
    .Z(_21261_));
 BUF_X8 _49313_ (.A(_21261_),
    .Z(_21262_));
 OAI21_X1 _49314_ (.A(_10739_),
    .B1(_21259_),
    .B2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.w_addr_i ),
    .ZN(_21263_));
 NOR2_X1 _49315_ (.A1(_21262_),
    .A2(_21263_),
    .ZN(_05407_));
 OR3_X1 _49316_ (.A1(_07604_),
    .A2(_07605_),
    .A3(lce_data_cmd_ready_i),
    .ZN(_21264_));
 INV_X1 _49317_ (.A(\icache.N8 ),
    .ZN(_21265_));
 NAND2_X2 _49318_ (.A1(_21265_),
    .A2(\icache.N10 ),
    .ZN(_21266_));
 AND4_X1 _49319_ (.A1(_00001_),
    .A2(_08480_),
    .A3(_08009_),
    .A4(_21266_),
    .ZN(_21267_));
 NAND3_X1 _49320_ (.A1(_21267_),
    .A2(_07618_),
    .A3(_20971_),
    .ZN(_21268_));
 OAI21_X1 _49321_ (.A(_21268_),
    .B1(_15261_),
    .B2(_15263_),
    .ZN(_21269_));
 OAI21_X1 _49322_ (.A(_21264_),
    .B1(_21269_),
    .B2(_07607_),
    .ZN(_21270_));
 AND2_X1 _49323_ (.A1(_10725_),
    .A2(lce_data_resp_ready_i),
    .ZN(_21271_));
 AND3_X1 _49324_ (.A1(_10732_),
    .A2(_07979_),
    .A3(_10733_),
    .ZN(_21272_));
 NAND2_X1 _49325_ (.A1(_20979_),
    .A2(_20973_),
    .ZN(_21273_));
 OAI221_X2 _49326_ (.A(_07889_),
    .B1(_20973_),
    .B2(_21271_),
    .C1(_21272_),
    .C2(_21273_),
    .ZN(_21274_));
 AND2_X1 _49327_ (.A1(_21270_),
    .A2(_21274_),
    .ZN(_21275_));
 INV_X1 _49328_ (.A(_21275_),
    .ZN(_21276_));
 NAND3_X1 _49329_ (.A1(_21276_),
    .A2(_07884_),
    .A3(_08723_),
    .ZN(_21277_));
 NAND4_X1 _49330_ (.A1(_21270_),
    .A2(_07973_),
    .A3(_21274_),
    .A4(_08662_),
    .ZN(_21278_));
 NAND2_X1 _49331_ (.A1(_21277_),
    .A2(_21278_),
    .ZN(_05406_));
 BUF_X8 _49332_ (.A(_08650_),
    .Z(_21279_));
 NAND3_X1 _49333_ (.A1(_10725_),
    .A2(_21258_),
    .A3(lce_cmd_v_i),
    .ZN(_21280_));
 AOI211_X1 _49334_ (.A(_21279_),
    .B(_21276_),
    .C1(_21258_),
    .C2(_21280_),
    .ZN(\icache.lce.lce_cmd_inst.rv_adapter.N14 ));
 INV_X1 _49335_ (.A(\icache.lce.lce_data_cmd.rv_adapter.full_r ),
    .ZN(_21281_));
 AND2_X2 _49336_ (.A1(_21281_),
    .A2(lce_data_cmd_v_i),
    .ZN(_21282_));
 INV_X1 _49337_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.w_addr_i ),
    .ZN(_21283_));
 OR3_X1 _49338_ (.A1(_21282_),
    .A2(_08650_),
    .A3(_21283_),
    .ZN(_21284_));
 NAND4_X1 _49339_ (.A1(_08723_),
    .A2(_21281_),
    .A3(_21283_),
    .A4(lce_data_cmd_v_i),
    .ZN(_21285_));
 NAND2_X1 _49340_ (.A1(_21284_),
    .A2(_21285_),
    .ZN(_05513_));
 NAND3_X1 _49341_ (.A1(_20982_),
    .A2(_08424_),
    .A3(_08723_),
    .ZN(_21286_));
 OAI211_X2 _49342_ (.A(_11248_),
    .B(_08662_),
    .C1(_15278_),
    .C2(_15281_),
    .ZN(_21287_));
 NAND2_X1 _49343_ (.A1(_21286_),
    .A2(_21287_),
    .ZN(_05512_));
 NAND3_X1 _49344_ (.A1(_08501_),
    .A2(_21281_),
    .A3(lce_data_cmd_v_i),
    .ZN(_21288_));
 AOI221_X4 _49345_ (.A(_08650_),
    .B1(_21281_),
    .B2(_21288_),
    .C1(_15280_),
    .C2(_00075_),
    .ZN(\icache.lce.lce_data_cmd.rv_adapter.N14 ));
 BUF_X8 _49346_ (.A(_10874_),
    .Z(_21289_));
 BUF_X32 _49347_ (.A(_10762_),
    .Z(_21290_));
 AND2_X4 _49348_ (.A1(_21289_),
    .A2(_21290_),
    .ZN(_21291_));
 BUF_X16 _49349_ (.A(_21291_),
    .Z(_21292_));
 BUF_X8 _49350_ (.A(_21292_),
    .Z(_21293_));
 MUX2_X1 _49351_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2744]),
    .B(_08524_),
    .S(_21293_),
    .Z(_02759_));
 MUX2_X1 _49352_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2745]),
    .B(_08529_),
    .S(_21293_),
    .Z(_02760_));
 BUF_X32 _49353_ (.A(fe_cmd_i[36]),
    .Z(_21294_));
 BUF_X8 _49354_ (.A(_21294_),
    .Z(_21295_));
 BUF_X8 _49355_ (.A(_21291_),
    .Z(_21296_));
 MUX2_X1 _49356_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2746]),
    .B(_21295_),
    .S(_21296_),
    .Z(_02761_));
 MUX2_X1 _49357_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2747]),
    .B(_08537_),
    .S(_21296_),
    .Z(_02762_));
 BUF_X32 _49358_ (.A(fe_cmd_i[38]),
    .Z(_21297_));
 BUF_X4 _49359_ (.A(_21297_),
    .Z(_21298_));
 MUX2_X1 _49360_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2748]),
    .B(_21298_),
    .S(_21296_),
    .Z(_02763_));
 BUF_X32 _49361_ (.A(fe_cmd_i[39]),
    .Z(_21299_));
 BUF_X8 _49362_ (.A(_21299_),
    .Z(_21300_));
 MUX2_X1 _49363_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2749]),
    .B(_21300_),
    .S(_21296_),
    .Z(_02764_));
 BUF_X32 _49364_ (.A(fe_cmd_i[40]),
    .Z(_21301_));
 BUF_X8 _49365_ (.A(_21301_),
    .Z(_21302_));
 MUX2_X1 _49366_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2750]),
    .B(_21302_),
    .S(_21296_),
    .Z(_02766_));
 BUF_X32 _49367_ (.A(fe_cmd_i[41]),
    .Z(_21303_));
 BUF_X4 _49368_ (.A(_21303_),
    .Z(_21304_));
 MUX2_X1 _49369_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2751]),
    .B(_21304_),
    .S(_21296_),
    .Z(_02767_));
 BUF_X32 _49370_ (.A(fe_cmd_i[42]),
    .Z(_21305_));
 BUF_X8 _49371_ (.A(_21305_),
    .Z(_21306_));
 MUX2_X1 _49372_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2752]),
    .B(_21306_),
    .S(_21296_),
    .Z(_02768_));
 BUF_X32 _49373_ (.A(fe_cmd_i[43]),
    .Z(_21307_));
 BUF_X8 _49374_ (.A(_21307_),
    .Z(_21308_));
 MUX2_X1 _49375_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2753]),
    .B(_21308_),
    .S(_21296_),
    .Z(_02769_));
 BUF_X32 _49376_ (.A(fe_cmd_i[44]),
    .Z(_21309_));
 BUF_X8 _49377_ (.A(_21309_),
    .Z(_21310_));
 MUX2_X1 _49378_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2754]),
    .B(_21310_),
    .S(_21296_),
    .Z(_02770_));
 BUF_X32 _49379_ (.A(fe_cmd_i[45]),
    .Z(_21311_));
 BUF_X8 _49380_ (.A(_21311_),
    .Z(_21312_));
 MUX2_X1 _49381_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2755]),
    .B(_21312_),
    .S(_21296_),
    .Z(_02771_));
 BUF_X8 _49382_ (.A(_21291_),
    .Z(_21313_));
 MUX2_X1 _49383_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2756]),
    .B(_10515_),
    .S(_21313_),
    .Z(_02772_));
 BUF_X8 _49384_ (.A(_10784_),
    .Z(_21314_));
 BUF_X8 _49385_ (.A(_21314_),
    .Z(_21315_));
 BUF_X8 _49386_ (.A(_10791_),
    .Z(_21316_));
 NAND4_X1 _49387_ (.A1(_10881_),
    .A2(_10569_),
    .A3(_21315_),
    .A4(_21316_),
    .ZN(_21317_));
 INV_X1 _49388_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2757]),
    .ZN(_21318_));
 OAI21_X1 _49389_ (.A(_21317_),
    .B1(_21293_),
    .B2(_21318_),
    .ZN(_02773_));
 MUX2_X1 _49390_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2758]),
    .B(_10529_),
    .S(_21313_),
    .Z(_02774_));
 MUX2_X1 _49391_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2759]),
    .B(_10530_),
    .S(_21313_),
    .Z(_02775_));
 MUX2_X1 _49392_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2760]),
    .B(_10531_),
    .S(_21313_),
    .Z(_02777_));
 MUX2_X1 _49393_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2761]),
    .B(_10532_),
    .S(_21313_),
    .Z(_02778_));
 MUX2_X1 _49394_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2762]),
    .B(_10533_),
    .S(_21313_),
    .Z(_02779_));
 MUX2_X1 _49395_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2763]),
    .B(_10534_),
    .S(_21313_),
    .Z(_02780_));
 MUX2_X1 _49396_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2764]),
    .B(_10535_),
    .S(_21313_),
    .Z(_02781_));
 MUX2_X1 _49397_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2765]),
    .B(_10536_),
    .S(_21313_),
    .Z(_02782_));
 MUX2_X1 _49398_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2766]),
    .B(_10538_),
    .S(_21313_),
    .Z(_02783_));
 BUF_X8 _49399_ (.A(_21291_),
    .Z(_21319_));
 MUX2_X1 _49400_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2767]),
    .B(_10539_),
    .S(_21319_),
    .Z(_02784_));
 MUX2_X1 _49401_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2768]),
    .B(_10540_),
    .S(_21319_),
    .Z(_02785_));
 NAND4_X2 _49402_ (.A1(_10881_),
    .A2(_10582_),
    .A3(_21315_),
    .A4(_21316_),
    .ZN(_21320_));
 INV_X1 _49403_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2769]),
    .ZN(_21321_));
 OAI21_X1 _49404_ (.A(_21320_),
    .B1(_21293_),
    .B2(_21321_),
    .ZN(_02786_));
 MUX2_X1 _49405_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2770]),
    .B(_10542_),
    .S(_21319_),
    .Z(_02788_));
 MUX2_X1 _49406_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2771]),
    .B(_10543_),
    .S(_21319_),
    .Z(_02789_));
 BUF_X8 _49407_ (.A(_10880_),
    .Z(_21322_));
 BUF_X8 _49408_ (.A(_10791_),
    .Z(_21323_));
 NAND4_X1 _49409_ (.A1(_21322_),
    .A2(_10585_),
    .A3(_21315_),
    .A4(_21323_),
    .ZN(_21324_));
 INV_X1 _49410_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2772]),
    .ZN(_21325_));
 OAI21_X1 _49411_ (.A(_21324_),
    .B1(_21293_),
    .B2(_21325_),
    .ZN(_02790_));
 NAND4_X1 _49412_ (.A1(_21322_),
    .A2(_10616_),
    .A3(_21315_),
    .A4(_21323_),
    .ZN(_21326_));
 INV_X1 _49413_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2773]),
    .ZN(_21327_));
 OAI21_X1 _49414_ (.A(_21326_),
    .B1(_21293_),
    .B2(_21327_),
    .ZN(_02791_));
 MUX2_X1 _49415_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2774]),
    .B(_10546_),
    .S(_21319_),
    .Z(_02792_));
 NAND4_X2 _49416_ (.A1(_21322_),
    .A2(_10588_),
    .A3(_21315_),
    .A4(_21323_),
    .ZN(_21328_));
 INV_X2 _49417_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2775]),
    .ZN(_21329_));
 OAI21_X1 _49418_ (.A(_21328_),
    .B1(_21293_),
    .B2(_21329_),
    .ZN(_02793_));
 MUX2_X1 _49419_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2776]),
    .B(_10548_),
    .S(_21319_),
    .Z(_02794_));
 MUX2_X1 _49420_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2777]),
    .B(_10549_),
    .S(_21319_),
    .Z(_02795_));
 MUX2_X1 _49421_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2778]),
    .B(_10550_),
    .S(_21319_),
    .Z(_02796_));
 MUX2_X1 _49422_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2779]),
    .B(_10551_),
    .S(_21319_),
    .Z(_02797_));
 MUX2_X1 _49423_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2780]),
    .B(_10552_),
    .S(_21319_),
    .Z(_02799_));
 BUF_X16 _49424_ (.A(_08632_),
    .Z(_21330_));
 NAND4_X1 _49425_ (.A1(_21322_),
    .A2(_21330_),
    .A3(_21315_),
    .A4(_21323_),
    .ZN(_21331_));
 INV_X1 _49426_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2781]),
    .ZN(_21332_));
 OAI21_X1 _49427_ (.A(_21331_),
    .B1(_21293_),
    .B2(_21332_),
    .ZN(_02800_));
 MUX2_X1 _49428_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2782]),
    .B(_10554_),
    .S(_21292_),
    .Z(_02801_));
 BUF_X4 _49429_ (.A(_08510_),
    .Z(_21333_));
 NAND2_X1 _49430_ (.A1(_21333_),
    .A2(fe_cmd_i[24]),
    .ZN(_21334_));
 BUF_X4 _49431_ (.A(_08326_),
    .Z(_21335_));
 BUF_X4 _49432_ (.A(_08027_),
    .Z(_21336_));
 BUF_X4 _49433_ (.A(fe_cmd_i[73]),
    .Z(_21337_));
 NAND4_X2 _49434_ (.A1(_21335_),
    .A2(_21336_),
    .A3(_21337_),
    .A4(fe_cmd_i[21]),
    .ZN(_21338_));
 NAND2_X4 _49435_ (.A1(_21334_),
    .A2(_21338_),
    .ZN(_21339_));
 BUF_X4 _49436_ (.A(_21339_),
    .Z(_21340_));
 MUX2_X1 _49437_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2783]),
    .B(_21340_),
    .S(_21292_),
    .Z(_02802_));
 NAND2_X1 _49438_ (.A1(_21333_),
    .A2(fe_cmd_i[25]),
    .ZN(_21341_));
 NAND4_X2 _49439_ (.A1(_21335_),
    .A2(_21336_),
    .A3(_21337_),
    .A4(fe_cmd_i[22]),
    .ZN(_21342_));
 NAND2_X4 _49440_ (.A1(_21341_),
    .A2(_21342_),
    .ZN(_21343_));
 BUF_X8 _49441_ (.A(_21343_),
    .Z(_21344_));
 MUX2_X1 _49442_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2784]),
    .B(_21344_),
    .S(_21292_),
    .Z(_02803_));
 NAND2_X1 _49443_ (.A1(_21333_),
    .A2(fe_cmd_i[26]),
    .ZN(_21345_));
 NAND4_X2 _49444_ (.A1(_21335_),
    .A2(_21336_),
    .A3(_21337_),
    .A4(fe_cmd_i[23]),
    .ZN(_21346_));
 NAND2_X4 _49445_ (.A1(_21345_),
    .A2(_21346_),
    .ZN(_21347_));
 BUF_X8 _49446_ (.A(_21347_),
    .Z(_21348_));
 MUX2_X1 _49447_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2785]),
    .B(_21348_),
    .S(_21292_),
    .Z(_02804_));
 NAND2_X1 _49448_ (.A1(_21333_),
    .A2(fe_cmd_i[27]),
    .ZN(_21349_));
 NAND4_X2 _49449_ (.A1(_21335_),
    .A2(_21336_),
    .A3(_21337_),
    .A4(fe_cmd_i[24]),
    .ZN(_21350_));
 NAND2_X4 _49450_ (.A1(_21349_),
    .A2(_21350_),
    .ZN(_21351_));
 BUF_X8 _49451_ (.A(_21351_),
    .Z(_21352_));
 MUX2_X1 _49452_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2786]),
    .B(_21352_),
    .S(_21292_),
    .Z(_02805_));
 NAND2_X1 _49453_ (.A1(_21333_),
    .A2(fe_cmd_i[28]),
    .ZN(_21353_));
 NAND4_X2 _49454_ (.A1(_21335_),
    .A2(_21336_),
    .A3(_21337_),
    .A4(fe_cmd_i[25]),
    .ZN(_21354_));
 NAND2_X4 _49455_ (.A1(_21353_),
    .A2(_21354_),
    .ZN(_21355_));
 BUF_X4 _49456_ (.A(_21355_),
    .Z(_21356_));
 MUX2_X1 _49457_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2787]),
    .B(_21356_),
    .S(_21292_),
    .Z(_02806_));
 NAND2_X1 _49458_ (.A1(_21333_),
    .A2(fe_cmd_i[29]),
    .ZN(_21357_));
 NAND4_X2 _49459_ (.A1(_21335_),
    .A2(_21336_),
    .A3(_21337_),
    .A4(fe_cmd_i[26]),
    .ZN(_21358_));
 NAND2_X4 _49460_ (.A1(_21357_),
    .A2(_21358_),
    .ZN(_21359_));
 BUF_X16 _49461_ (.A(_21359_),
    .Z(_21360_));
 NAND4_X1 _49462_ (.A1(_21322_),
    .A2(_11193_),
    .A3(_10792_),
    .A4(_21360_),
    .ZN(_21361_));
 INV_X1 _49463_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2788]),
    .ZN(_21362_));
 OAI21_X1 _49464_ (.A(_21361_),
    .B1(_21293_),
    .B2(_21362_),
    .ZN(_02807_));
 NAND2_X1 _49465_ (.A1(_21333_),
    .A2(fe_cmd_i[30]),
    .ZN(_21363_));
 NAND4_X2 _49466_ (.A1(_21335_),
    .A2(_21336_),
    .A3(fe_cmd_i[73]),
    .A4(fe_cmd_i[27]),
    .ZN(_21364_));
 NAND2_X4 _49467_ (.A1(_21363_),
    .A2(_21364_),
    .ZN(_21365_));
 BUF_X4 _49468_ (.A(_21365_),
    .Z(_21366_));
 MUX2_X1 _49469_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2789]),
    .B(_21366_),
    .S(_21292_),
    .Z(_02808_));
 NAND2_X1 _49470_ (.A1(_21333_),
    .A2(fe_cmd_i[31]),
    .ZN(_21367_));
 NAND4_X2 _49471_ (.A1(_21335_),
    .A2(_21336_),
    .A3(_21337_),
    .A4(fe_cmd_i[28]),
    .ZN(_21368_));
 NAND2_X4 _49472_ (.A1(_21367_),
    .A2(_21368_),
    .ZN(_21369_));
 BUF_X8 _49473_ (.A(_21369_),
    .Z(_21370_));
 MUX2_X1 _49474_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2790]),
    .B(_21370_),
    .S(_21292_),
    .Z(_02810_));
 NAND2_X1 _49475_ (.A1(_21333_),
    .A2(fe_cmd_i[32]),
    .ZN(_21371_));
 NAND4_X2 _49476_ (.A1(_21335_),
    .A2(_21336_),
    .A3(_21337_),
    .A4(fe_cmd_i[29]),
    .ZN(_21372_));
 NAND2_X4 _49477_ (.A1(_21371_),
    .A2(_21372_),
    .ZN(_21373_));
 BUF_X4 _49478_ (.A(_21373_),
    .Z(_21374_));
 MUX2_X1 _49479_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2791]),
    .B(_21374_),
    .S(_21292_),
    .Z(_02811_));
 NAND2_X1 _49480_ (.A1(_21333_),
    .A2(_10741_),
    .ZN(_21375_));
 NAND4_X2 _49481_ (.A1(_21335_),
    .A2(_21336_),
    .A3(_21337_),
    .A4(fe_cmd_i[30]),
    .ZN(_21376_));
 NAND2_X4 _49482_ (.A1(_21375_),
    .A2(_21376_),
    .ZN(_21377_));
 NAND4_X1 _49483_ (.A1(_21322_),
    .A2(_11193_),
    .A3(_10792_),
    .A4(_21377_),
    .ZN(_21378_));
 INV_X1 _49484_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2792]),
    .ZN(_21379_));
 OAI21_X1 _49485_ (.A(_21378_),
    .B1(_21293_),
    .B2(_21379_),
    .ZN(_02812_));
 AND2_X4 _49486_ (.A1(_10799_),
    .A2(_21290_),
    .ZN(_21380_));
 BUF_X8 _49487_ (.A(_21380_),
    .Z(_21381_));
 BUF_X8 _49488_ (.A(_21381_),
    .Z(_21382_));
 MUX2_X1 _49489_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3087]),
    .B(_08524_),
    .S(_21382_),
    .Z(_03140_));
 MUX2_X1 _49490_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3088]),
    .B(_08529_),
    .S(_21382_),
    .Z(_03141_));
 BUF_X16 _49491_ (.A(_21294_),
    .Z(_21383_));
 NAND4_X1 _49492_ (.A1(_10806_),
    .A2(_21383_),
    .A3(_21315_),
    .A4(_21323_),
    .ZN(_21384_));
 INV_X1 _49493_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3089]),
    .ZN(_21385_));
 OAI21_X1 _49494_ (.A(_21384_),
    .B1(_21382_),
    .B2(_21385_),
    .ZN(_03142_));
 BUF_X8 _49495_ (.A(_21380_),
    .Z(_21386_));
 MUX2_X1 _49496_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3090]),
    .B(_08537_),
    .S(_21386_),
    .Z(_03144_));
 BUF_X16 _49497_ (.A(_21297_),
    .Z(_21387_));
 BUF_X4 _49498_ (.A(_21314_),
    .Z(_21388_));
 NAND4_X1 _49499_ (.A1(_10806_),
    .A2(_21387_),
    .A3(_21388_),
    .A4(_21323_),
    .ZN(_21389_));
 INV_X1 _49500_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3091]),
    .ZN(_21390_));
 OAI21_X1 _49501_ (.A(_21389_),
    .B1(_21382_),
    .B2(_21390_),
    .ZN(_03145_));
 MUX2_X1 _49502_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3092]),
    .B(_21300_),
    .S(_21386_),
    .Z(_03146_));
 MUX2_X1 _49503_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3093]),
    .B(_21302_),
    .S(_21386_),
    .Z(_03147_));
 MUX2_X1 _49504_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3094]),
    .B(_21304_),
    .S(_21386_),
    .Z(_03148_));
 BUF_X8 _49505_ (.A(_10805_),
    .Z(_21391_));
 BUF_X32 _49506_ (.A(_21305_),
    .Z(_21392_));
 NAND4_X1 _49507_ (.A1(_21391_),
    .A2(_21392_),
    .A3(_21388_),
    .A4(_21323_),
    .ZN(_21393_));
 INV_X1 _49508_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3095]),
    .ZN(_21394_));
 OAI21_X1 _49509_ (.A(_21393_),
    .B1(_21382_),
    .B2(_21394_),
    .ZN(_03149_));
 BUF_X16 _49510_ (.A(_21307_),
    .Z(_21395_));
 NAND4_X1 _49511_ (.A1(_21391_),
    .A2(_21395_),
    .A3(_21388_),
    .A4(_21323_),
    .ZN(_21396_));
 INV_X4 _49512_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3096]),
    .ZN(_21397_));
 OAI21_X1 _49513_ (.A(_21396_),
    .B1(_21382_),
    .B2(_21397_),
    .ZN(_03150_));
 MUX2_X1 _49514_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3097]),
    .B(_21310_),
    .S(_21386_),
    .Z(_03151_));
 MUX2_X1 _49515_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3098]),
    .B(_21312_),
    .S(_21386_),
    .Z(_03152_));
 MUX2_X1 _49516_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3099]),
    .B(_10515_),
    .S(_21386_),
    .Z(_03153_));
 MUX2_X1 _49517_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3100]),
    .B(_10528_),
    .S(_21386_),
    .Z(_03156_));
 MUX2_X1 _49518_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3101]),
    .B(_10529_),
    .S(_21386_),
    .Z(_03157_));
 MUX2_X1 _49519_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3102]),
    .B(_10530_),
    .S(_21386_),
    .Z(_03158_));
 BUF_X8 _49520_ (.A(_21380_),
    .Z(_21398_));
 MUX2_X1 _49521_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3103]),
    .B(_10531_),
    .S(_21398_),
    .Z(_03159_));
 MUX2_X1 _49522_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3104]),
    .B(_10532_),
    .S(_21398_),
    .Z(_03160_));
 MUX2_X1 _49523_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3105]),
    .B(_10533_),
    .S(_21398_),
    .Z(_03161_));
 MUX2_X1 _49524_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3106]),
    .B(_10534_),
    .S(_21398_),
    .Z(_03162_));
 MUX2_X1 _49525_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3107]),
    .B(_10535_),
    .S(_21398_),
    .Z(_03163_));
 MUX2_X1 _49526_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3108]),
    .B(_10536_),
    .S(_21398_),
    .Z(_03164_));
 MUX2_X1 _49527_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3109]),
    .B(_10538_),
    .S(_21398_),
    .Z(_03165_));
 NAND4_X1 _49528_ (.A1(_21391_),
    .A2(_10580_),
    .A3(_21388_),
    .A4(_21323_),
    .ZN(_21399_));
 INV_X1 _49529_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3110]),
    .ZN(_21400_));
 OAI21_X1 _49530_ (.A(_21399_),
    .B1(_21382_),
    .B2(_21400_),
    .ZN(_03167_));
 MUX2_X1 _49531_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3111]),
    .B(_10540_),
    .S(_21398_),
    .Z(_03168_));
 NAND4_X1 _49532_ (.A1(_21391_),
    .A2(_10582_),
    .A3(_21388_),
    .A4(_21323_),
    .ZN(_21401_));
 INV_X1 _49533_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3112]),
    .ZN(_21402_));
 OAI21_X1 _49534_ (.A(_21401_),
    .B1(_21382_),
    .B2(_21402_),
    .ZN(_03169_));
 MUX2_X1 _49535_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3113]),
    .B(_10542_),
    .S(_21398_),
    .Z(_03170_));
 MUX2_X1 _49536_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3114]),
    .B(_10543_),
    .S(_21398_),
    .Z(_03171_));
 BUF_X8 _49537_ (.A(_21380_),
    .Z(_21403_));
 MUX2_X1 _49538_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3115]),
    .B(_10544_),
    .S(_21403_),
    .Z(_03172_));
 MUX2_X1 _49539_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3116]),
    .B(_10545_),
    .S(_21403_),
    .Z(_03173_));
 MUX2_X1 _49540_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3117]),
    .B(_10546_),
    .S(_21403_),
    .Z(_03174_));
 MUX2_X1 _49541_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3118]),
    .B(_10547_),
    .S(_21403_),
    .Z(_03175_));
 MUX2_X1 _49542_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3119]),
    .B(_10548_),
    .S(_21403_),
    .Z(_03176_));
 MUX2_X1 _49543_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3120]),
    .B(_10549_),
    .S(_21403_),
    .Z(_03178_));
 BUF_X4 _49544_ (.A(_10791_),
    .Z(_21404_));
 NAND4_X1 _49545_ (.A1(_21391_),
    .A2(_10591_),
    .A3(_21388_),
    .A4(_21404_),
    .ZN(_21405_));
 INV_X1 _49546_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3121]),
    .ZN(_21406_));
 OAI21_X1 _49547_ (.A(_21405_),
    .B1(_21382_),
    .B2(_21406_),
    .ZN(_03179_));
 MUX2_X1 _49548_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3122]),
    .B(_10551_),
    .S(_21403_),
    .Z(_03180_));
 MUX2_X1 _49549_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3123]),
    .B(_10552_),
    .S(_21403_),
    .Z(_03181_));
 MUX2_X1 _49550_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3124]),
    .B(_10553_),
    .S(_21403_),
    .Z(_03182_));
 MUX2_X1 _49551_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3125]),
    .B(_10554_),
    .S(_21403_),
    .Z(_03183_));
 MUX2_X1 _49552_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3126]),
    .B(_21340_),
    .S(_21381_),
    .Z(_03184_));
 MUX2_X1 _49553_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3127]),
    .B(_21344_),
    .S(_21381_),
    .Z(_03185_));
 BUF_X16 _49554_ (.A(_21347_),
    .Z(_21407_));
 NAND4_X1 _49555_ (.A1(_21391_),
    .A2(_11193_),
    .A3(_21316_),
    .A4(_21407_),
    .ZN(_21408_));
 INV_X4 _49556_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3128]),
    .ZN(_21409_));
 OAI21_X1 _49557_ (.A(_21408_),
    .B1(_21382_),
    .B2(_21409_),
    .ZN(_03186_));
 MUX2_X1 _49558_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3129]),
    .B(_21352_),
    .S(_21381_),
    .Z(_03187_));
 MUX2_X1 _49559_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3130]),
    .B(_21356_),
    .S(_21381_),
    .Z(_03189_));
 BUF_X8 _49560_ (.A(_21359_),
    .Z(_21410_));
 MUX2_X1 _49561_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3131]),
    .B(_21410_),
    .S(_21381_),
    .Z(_03190_));
 MUX2_X1 _49562_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3132]),
    .B(_21366_),
    .S(_21381_),
    .Z(_03191_));
 MUX2_X1 _49563_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3133]),
    .B(_21370_),
    .S(_21381_),
    .Z(_03192_));
 MUX2_X1 _49564_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3134]),
    .B(_21374_),
    .S(_21381_),
    .Z(_03193_));
 BUF_X8 _49565_ (.A(_21377_),
    .Z(_21411_));
 MUX2_X1 _49566_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3135]),
    .B(_21411_),
    .S(_21381_),
    .Z(_03194_));
 BUF_X32 _49567_ (.A(_10762_),
    .Z(_21412_));
 AND2_X4 _49568_ (.A1(_10812_),
    .A2(_21412_),
    .ZN(_21413_));
 BUF_X8 _49569_ (.A(_21413_),
    .Z(_21414_));
 BUF_X8 _49570_ (.A(_21414_),
    .Z(_21415_));
 MUX2_X1 _49571_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3038]),
    .B(_08524_),
    .S(_21415_),
    .Z(_03086_));
 MUX2_X1 _49572_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3039]),
    .B(_08529_),
    .S(_21415_),
    .Z(_03087_));
 NAND4_X1 _49573_ (.A1(_10820_),
    .A2(_21383_),
    .A3(_21388_),
    .A4(_21404_),
    .ZN(_21416_));
 INV_X1 _49574_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3040]),
    .ZN(_21417_));
 OAI21_X1 _49575_ (.A(_21416_),
    .B1(_21415_),
    .B2(_21417_),
    .ZN(_03089_));
 MUX2_X1 _49576_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3041]),
    .B(_08537_),
    .S(_21415_),
    .Z(_03090_));
 BUF_X32 _49577_ (.A(_21297_),
    .Z(_21418_));
 NAND4_X1 _49578_ (.A1(_10820_),
    .A2(_21418_),
    .A3(_21388_),
    .A4(_21404_),
    .ZN(_21419_));
 INV_X1 _49579_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3042]),
    .ZN(_21420_));
 OAI21_X1 _49580_ (.A(_21419_),
    .B1(_21415_),
    .B2(_21420_),
    .ZN(_03091_));
 MUX2_X1 _49581_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3043]),
    .B(_21300_),
    .S(_21415_),
    .Z(_03092_));
 MUX2_X1 _49582_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3044]),
    .B(_21302_),
    .S(_21415_),
    .Z(_03093_));
 BUF_X8 _49583_ (.A(_21413_),
    .Z(_21421_));
 MUX2_X1 _49584_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3045]),
    .B(_21304_),
    .S(_21421_),
    .Z(_03094_));
 BUF_X8 _49585_ (.A(_10819_),
    .Z(_21422_));
 NAND4_X1 _49586_ (.A1(_21422_),
    .A2(_21392_),
    .A3(_21388_),
    .A4(_21404_),
    .ZN(_21423_));
 INV_X1 _49587_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3046]),
    .ZN(_21424_));
 OAI21_X1 _49588_ (.A(_21423_),
    .B1(_21415_),
    .B2(_21424_),
    .ZN(_03095_));
 MUX2_X1 _49589_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3047]),
    .B(_21308_),
    .S(_21421_),
    .Z(_03096_));
 MUX2_X1 _49590_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3048]),
    .B(_21310_),
    .S(_21421_),
    .Z(_03097_));
 MUX2_X1 _49591_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3049]),
    .B(_21312_),
    .S(_21421_),
    .Z(_03098_));
 MUX2_X1 _49592_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3050]),
    .B(_10515_),
    .S(_21421_),
    .Z(_03100_));
 MUX2_X1 _49593_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3051]),
    .B(_10528_),
    .S(_21421_),
    .Z(_03101_));
 MUX2_X1 _49594_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3052]),
    .B(_10529_),
    .S(_21421_),
    .Z(_03102_));
 MUX2_X1 _49595_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3053]),
    .B(_10530_),
    .S(_21421_),
    .Z(_03103_));
 MUX2_X1 _49596_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3054]),
    .B(_10531_),
    .S(_21421_),
    .Z(_03104_));
 MUX2_X1 _49597_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3055]),
    .B(_10532_),
    .S(_21421_),
    .Z(_03105_));
 BUF_X8 _49598_ (.A(_21413_),
    .Z(_21425_));
 MUX2_X1 _49599_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3056]),
    .B(_10533_),
    .S(_21425_),
    .Z(_03106_));
 MUX2_X1 _49600_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3057]),
    .B(_10534_),
    .S(_21425_),
    .Z(_03107_));
 MUX2_X1 _49601_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3058]),
    .B(_10535_),
    .S(_21425_),
    .Z(_03108_));
 MUX2_X1 _49602_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3059]),
    .B(_10536_),
    .S(_21425_),
    .Z(_03109_));
 MUX2_X1 _49603_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3060]),
    .B(_10538_),
    .S(_21425_),
    .Z(_03111_));
 MUX2_X1 _49604_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3061]),
    .B(_10539_),
    .S(_21425_),
    .Z(_03112_));
 MUX2_X1 _49605_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3062]),
    .B(_10540_),
    .S(_21425_),
    .Z(_03113_));
 NAND4_X1 _49606_ (.A1(_21422_),
    .A2(_10582_),
    .A3(_21388_),
    .A4(_21404_),
    .ZN(_21426_));
 INV_X1 _49607_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3063]),
    .ZN(_21427_));
 OAI21_X1 _49608_ (.A(_21426_),
    .B1(_21415_),
    .B2(_21427_),
    .ZN(_03114_));
 MUX2_X1 _49609_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3064]),
    .B(_10542_),
    .S(_21425_),
    .Z(_03115_));
 MUX2_X1 _49610_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3065]),
    .B(_10543_),
    .S(_21425_),
    .Z(_03116_));
 MUX2_X1 _49611_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3066]),
    .B(_10544_),
    .S(_21425_),
    .Z(_03117_));
 BUF_X8 _49612_ (.A(_21413_),
    .Z(_21428_));
 MUX2_X1 _49613_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3067]),
    .B(_10545_),
    .S(_21428_),
    .Z(_03118_));
 MUX2_X1 _49614_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3068]),
    .B(_10546_),
    .S(_21428_),
    .Z(_03119_));
 MUX2_X1 _49615_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3069]),
    .B(_10547_),
    .S(_21428_),
    .Z(_03120_));
 MUX2_X1 _49616_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3070]),
    .B(_10548_),
    .S(_21428_),
    .Z(_03122_));
 MUX2_X1 _49617_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3071]),
    .B(_10549_),
    .S(_21428_),
    .Z(_03123_));
 BUF_X8 _49618_ (.A(_21314_),
    .Z(_21429_));
 NAND4_X1 _49619_ (.A1(_21422_),
    .A2(_10591_),
    .A3(_21429_),
    .A4(_21404_),
    .ZN(_21430_));
 INV_X1 _49620_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3072]),
    .ZN(_21431_));
 OAI21_X1 _49621_ (.A(_21430_),
    .B1(_21415_),
    .B2(_21431_),
    .ZN(_03124_));
 MUX2_X1 _49622_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3073]),
    .B(_10551_),
    .S(_21428_),
    .Z(_03125_));
 MUX2_X1 _49623_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3074]),
    .B(_10552_),
    .S(_21428_),
    .Z(_03126_));
 MUX2_X1 _49624_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3075]),
    .B(_10553_),
    .S(_21428_),
    .Z(_03127_));
 MUX2_X1 _49625_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3076]),
    .B(_10554_),
    .S(_21428_),
    .Z(_03128_));
 MUX2_X1 _49626_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3077]),
    .B(_21340_),
    .S(_21428_),
    .Z(_03129_));
 MUX2_X1 _49627_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3078]),
    .B(_21344_),
    .S(_21414_),
    .Z(_03130_));
 MUX2_X1 _49628_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3079]),
    .B(_21348_),
    .S(_21414_),
    .Z(_03131_));
 MUX2_X1 _49629_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3080]),
    .B(_21352_),
    .S(_21414_),
    .Z(_03133_));
 MUX2_X1 _49630_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3081]),
    .B(_21356_),
    .S(_21414_),
    .Z(_03134_));
 MUX2_X1 _49631_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3082]),
    .B(_21410_),
    .S(_21414_),
    .Z(_03135_));
 MUX2_X1 _49632_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3083]),
    .B(_21366_),
    .S(_21414_),
    .Z(_03136_));
 MUX2_X1 _49633_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3084]),
    .B(_21370_),
    .S(_21414_),
    .Z(_03137_));
 MUX2_X1 _49634_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3085]),
    .B(_21374_),
    .S(_21414_),
    .Z(_03138_));
 MUX2_X1 _49635_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3086]),
    .B(_21411_),
    .S(_21414_),
    .Z(_03139_));
 BUF_X32 _49636_ (.A(_10762_),
    .Z(_21432_));
 AND2_X4 _49637_ (.A1(_10826_),
    .A2(_21432_),
    .ZN(_21433_));
 BUF_X8 _49638_ (.A(_21433_),
    .Z(_21434_));
 BUF_X8 _49639_ (.A(_21434_),
    .Z(_21435_));
 MUX2_X1 _49640_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2989]),
    .B(_08524_),
    .S(_21435_),
    .Z(_03030_));
 MUX2_X1 _49641_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2990]),
    .B(_08529_),
    .S(_21435_),
    .Z(_03032_));
 MUX2_X1 _49642_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2991]),
    .B(_21295_),
    .S(_21435_),
    .Z(_03033_));
 MUX2_X1 _49643_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2992]),
    .B(_08537_),
    .S(_21435_),
    .Z(_03034_));
 MUX2_X1 _49644_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2993]),
    .B(_21298_),
    .S(_21435_),
    .Z(_03035_));
 MUX2_X1 _49645_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2994]),
    .B(_21300_),
    .S(_21435_),
    .Z(_03036_));
 MUX2_X1 _49646_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2995]),
    .B(_21302_),
    .S(_21435_),
    .Z(_03037_));
 MUX2_X1 _49647_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2996]),
    .B(_21304_),
    .S(_21435_),
    .Z(_03038_));
 MUX2_X1 _49648_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2997]),
    .B(_21306_),
    .S(_21435_),
    .Z(_03039_));
 BUF_X8 _49649_ (.A(_21433_),
    .Z(_21436_));
 MUX2_X1 _49650_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2998]),
    .B(_21308_),
    .S(_21436_),
    .Z(_03040_));
 MUX2_X1 _49651_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2999]),
    .B(_21310_),
    .S(_21436_),
    .Z(_03041_));
 MUX2_X1 _49652_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3000]),
    .B(_21312_),
    .S(_21436_),
    .Z(_03045_));
 MUX2_X1 _49653_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3001]),
    .B(_10515_),
    .S(_21436_),
    .Z(_03046_));
 MUX2_X1 _49654_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3002]),
    .B(_10528_),
    .S(_21436_),
    .Z(_03047_));
 MUX2_X1 _49655_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3003]),
    .B(_10529_),
    .S(_21436_),
    .Z(_03048_));
 MUX2_X1 _49656_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3004]),
    .B(_10530_),
    .S(_21436_),
    .Z(_03049_));
 MUX2_X1 _49657_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3005]),
    .B(_10531_),
    .S(_21436_),
    .Z(_03050_));
 MUX2_X1 _49658_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3006]),
    .B(_10532_),
    .S(_21436_),
    .Z(_03051_));
 MUX2_X1 _49659_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3007]),
    .B(_10533_),
    .S(_21436_),
    .Z(_03052_));
 BUF_X8 _49660_ (.A(_21433_),
    .Z(_21437_));
 MUX2_X1 _49661_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3008]),
    .B(_10534_),
    .S(_21437_),
    .Z(_03053_));
 MUX2_X1 _49662_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3009]),
    .B(_10535_),
    .S(_21437_),
    .Z(_03054_));
 MUX2_X1 _49663_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3010]),
    .B(_10536_),
    .S(_21437_),
    .Z(_03056_));
 MUX2_X1 _49664_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3011]),
    .B(_10538_),
    .S(_21437_),
    .Z(_03057_));
 NAND4_X1 _49665_ (.A1(_10833_),
    .A2(_10580_),
    .A3(_21429_),
    .A4(_21404_),
    .ZN(_21438_));
 INV_X1 _49666_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3012]),
    .ZN(_21439_));
 OAI21_X1 _49667_ (.A(_21438_),
    .B1(_21435_),
    .B2(_21439_),
    .ZN(_03058_));
 MUX2_X1 _49668_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3013]),
    .B(_10540_),
    .S(_21437_),
    .Z(_03059_));
 MUX2_X1 _49669_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3014]),
    .B(_10541_),
    .S(_21437_),
    .Z(_03060_));
 MUX2_X1 _49670_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3015]),
    .B(_10542_),
    .S(_21437_),
    .Z(_03061_));
 MUX2_X1 _49671_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3016]),
    .B(_10543_),
    .S(_21437_),
    .Z(_03062_));
 MUX2_X1 _49672_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3017]),
    .B(_10544_),
    .S(_21437_),
    .Z(_03063_));
 MUX2_X1 _49673_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3018]),
    .B(_10545_),
    .S(_21437_),
    .Z(_03064_));
 BUF_X8 _49674_ (.A(_21433_),
    .Z(_21440_));
 MUX2_X1 _49675_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3019]),
    .B(_10546_),
    .S(_21440_),
    .Z(_03065_));
 MUX2_X1 _49676_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3020]),
    .B(_10547_),
    .S(_21440_),
    .Z(_03067_));
 MUX2_X1 _49677_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3021]),
    .B(_10548_),
    .S(_21440_),
    .Z(_03068_));
 MUX2_X1 _49678_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3022]),
    .B(_10549_),
    .S(_21440_),
    .Z(_03069_));
 MUX2_X1 _49679_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3023]),
    .B(_10550_),
    .S(_21440_),
    .Z(_03070_));
 MUX2_X1 _49680_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3024]),
    .B(_10551_),
    .S(_21440_),
    .Z(_03071_));
 MUX2_X1 _49681_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3025]),
    .B(_10552_),
    .S(_21440_),
    .Z(_03072_));
 MUX2_X1 _49682_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3026]),
    .B(_10553_),
    .S(_21440_),
    .Z(_03073_));
 MUX2_X1 _49683_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3027]),
    .B(_10554_),
    .S(_21440_),
    .Z(_03074_));
 MUX2_X1 _49684_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3028]),
    .B(_21340_),
    .S(_21440_),
    .Z(_03075_));
 MUX2_X1 _49685_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3029]),
    .B(_21344_),
    .S(_21434_),
    .Z(_03076_));
 MUX2_X1 _49686_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3030]),
    .B(_21348_),
    .S(_21434_),
    .Z(_03078_));
 MUX2_X1 _49687_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3031]),
    .B(_21352_),
    .S(_21434_),
    .Z(_03079_));
 MUX2_X1 _49688_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3032]),
    .B(_21356_),
    .S(_21434_),
    .Z(_03080_));
 MUX2_X1 _49689_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3033]),
    .B(_21410_),
    .S(_21434_),
    .Z(_03081_));
 MUX2_X1 _49690_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3034]),
    .B(_21366_),
    .S(_21434_),
    .Z(_03082_));
 MUX2_X1 _49691_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3035]),
    .B(_21370_),
    .S(_21434_),
    .Z(_03083_));
 MUX2_X1 _49692_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3036]),
    .B(_21374_),
    .S(_21434_),
    .Z(_03084_));
 MUX2_X1 _49693_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3037]),
    .B(_21411_),
    .S(_21434_),
    .Z(_03085_));
 BUF_X32 _49694_ (.A(_10762_),
    .Z(_21441_));
 AND2_X4 _49695_ (.A1(_10838_),
    .A2(_21441_),
    .ZN(_21442_));
 BUF_X8 _49696_ (.A(_21442_),
    .Z(_21443_));
 BUF_X8 _49697_ (.A(_21443_),
    .Z(_21444_));
 MUX2_X1 _49698_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2940]),
    .B(_08524_),
    .S(_21444_),
    .Z(_02977_));
 MUX2_X1 _49699_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2941]),
    .B(_08529_),
    .S(_21444_),
    .Z(_02978_));
 MUX2_X1 _49700_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2942]),
    .B(_21295_),
    .S(_21444_),
    .Z(_02979_));
 BUF_X8 _49701_ (.A(_21442_),
    .Z(_21445_));
 MUX2_X1 _49702_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2943]),
    .B(_08537_),
    .S(_21445_),
    .Z(_02980_));
 MUX2_X1 _49703_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2944]),
    .B(_21298_),
    .S(_21445_),
    .Z(_02981_));
 MUX2_X1 _49704_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2945]),
    .B(_21300_),
    .S(_21445_),
    .Z(_02982_));
 MUX2_X1 _49705_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2946]),
    .B(_21302_),
    .S(_21445_),
    .Z(_02983_));
 MUX2_X1 _49706_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2947]),
    .B(_21304_),
    .S(_21445_),
    .Z(_02984_));
 MUX2_X1 _49707_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2948]),
    .B(_21306_),
    .S(_21445_),
    .Z(_02985_));
 MUX2_X1 _49708_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2949]),
    .B(_21308_),
    .S(_21445_),
    .Z(_02986_));
 BUF_X16 _49709_ (.A(_21309_),
    .Z(_21446_));
 NAND4_X1 _49710_ (.A1(_10846_),
    .A2(_21446_),
    .A3(_21429_),
    .A4(_21404_),
    .ZN(_21447_));
 INV_X2 _49711_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2950]),
    .ZN(_21448_));
 OAI21_X1 _49712_ (.A(_21447_),
    .B1(_21444_),
    .B2(_21448_),
    .ZN(_02988_));
 MUX2_X1 _49713_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2951]),
    .B(_21312_),
    .S(_21445_),
    .Z(_02989_));
 MUX2_X1 _49714_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2952]),
    .B(_10515_),
    .S(_21445_),
    .Z(_02990_));
 NAND4_X1 _49715_ (.A1(_10846_),
    .A2(_10569_),
    .A3(_21429_),
    .A4(_21404_),
    .ZN(_21449_));
 INV_X1 _49716_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2953]),
    .ZN(_21450_));
 OAI21_X1 _49717_ (.A(_21449_),
    .B1(_21444_),
    .B2(_21450_),
    .ZN(_02991_));
 MUX2_X1 _49718_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2954]),
    .B(_10529_),
    .S(_21445_),
    .Z(_02992_));
 BUF_X8 _49719_ (.A(_21442_),
    .Z(_21451_));
 MUX2_X1 _49720_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2955]),
    .B(_10530_),
    .S(_21451_),
    .Z(_02993_));
 MUX2_X1 _49721_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2956]),
    .B(_10531_),
    .S(_21451_),
    .Z(_02994_));
 BUF_X8 _49722_ (.A(_10845_),
    .Z(_21452_));
 NAND4_X1 _49723_ (.A1(_21452_),
    .A2(_10599_),
    .A3(_21429_),
    .A4(_21404_),
    .ZN(_21453_));
 INV_X1 _49724_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2957]),
    .ZN(_21454_));
 OAI21_X1 _49725_ (.A(_21453_),
    .B1(_21444_),
    .B2(_21454_),
    .ZN(_02995_));
 MUX2_X1 _49726_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2958]),
    .B(_10533_),
    .S(_21451_),
    .Z(_02996_));
 MUX2_X1 _49727_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2959]),
    .B(_10534_),
    .S(_21451_),
    .Z(_02997_));
 MUX2_X1 _49728_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2960]),
    .B(_10535_),
    .S(_21451_),
    .Z(_02999_));
 MUX2_X1 _49729_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2961]),
    .B(_10536_),
    .S(_21451_),
    .Z(_03000_));
 MUX2_X1 _49730_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2962]),
    .B(_10538_),
    .S(_21451_),
    .Z(_03001_));
 MUX2_X1 _49731_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2963]),
    .B(_10539_),
    .S(_21451_),
    .Z(_03002_));
 MUX2_X1 _49732_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2964]),
    .B(_10540_),
    .S(_21451_),
    .Z(_03003_));
 MUX2_X1 _49733_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2965]),
    .B(_10541_),
    .S(_21451_),
    .Z(_03004_));
 BUF_X8 _49734_ (.A(_21442_),
    .Z(_21455_));
 MUX2_X1 _49735_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2966]),
    .B(_10542_),
    .S(_21455_),
    .Z(_03005_));
 MUX2_X1 _49736_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2967]),
    .B(_10543_),
    .S(_21455_),
    .Z(_03006_));
 BUF_X4 _49737_ (.A(_10791_),
    .Z(_21456_));
 NAND4_X1 _49738_ (.A1(_21452_),
    .A2(_10585_),
    .A3(_21429_),
    .A4(_21456_),
    .ZN(_21457_));
 INV_X1 _49739_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2968]),
    .ZN(_21458_));
 OAI21_X1 _49740_ (.A(_21457_),
    .B1(_21444_),
    .B2(_21458_),
    .ZN(_03007_));
 MUX2_X1 _49741_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2969]),
    .B(_10545_),
    .S(_21455_),
    .Z(_03008_));
 MUX2_X1 _49742_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2970]),
    .B(_10546_),
    .S(_21455_),
    .Z(_03010_));
 MUX2_X1 _49743_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2971]),
    .B(_10547_),
    .S(_21455_),
    .Z(_03011_));
 MUX2_X1 _49744_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2972]),
    .B(_10548_),
    .S(_21455_),
    .Z(_03012_));
 MUX2_X1 _49745_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2973]),
    .B(_10549_),
    .S(_21455_),
    .Z(_03013_));
 MUX2_X1 _49746_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2974]),
    .B(_10550_),
    .S(_21455_),
    .Z(_03014_));
 MUX2_X1 _49747_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2975]),
    .B(_10551_),
    .S(_21455_),
    .Z(_03015_));
 MUX2_X1 _49748_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2976]),
    .B(_10552_),
    .S(_21455_),
    .Z(_03016_));
 NAND4_X1 _49749_ (.A1(_21452_),
    .A2(_21330_),
    .A3(_21429_),
    .A4(_21456_),
    .ZN(_21459_));
 INV_X1 _49750_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2977]),
    .ZN(_21460_));
 OAI21_X1 _49751_ (.A(_21459_),
    .B1(_21444_),
    .B2(_21460_),
    .ZN(_03017_));
 MUX2_X1 _49752_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2978]),
    .B(_10554_),
    .S(_21443_),
    .Z(_03018_));
 MUX2_X1 _49753_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2979]),
    .B(_21340_),
    .S(_21443_),
    .Z(_03019_));
 MUX2_X1 _49754_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2980]),
    .B(_21344_),
    .S(_21443_),
    .Z(_03021_));
 MUX2_X1 _49755_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2981]),
    .B(_21348_),
    .S(_21443_),
    .Z(_03022_));
 BUF_X8 _49756_ (.A(_21351_),
    .Z(_21461_));
 NAND4_X1 _49757_ (.A1(_21452_),
    .A2(_11193_),
    .A3(_21316_),
    .A4(_21461_),
    .ZN(_21462_));
 INV_X2 _49758_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2982]),
    .ZN(_21463_));
 OAI21_X1 _49759_ (.A(_21462_),
    .B1(_21444_),
    .B2(_21463_),
    .ZN(_03023_));
 MUX2_X1 _49760_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2983]),
    .B(_21356_),
    .S(_21443_),
    .Z(_03024_));
 NAND4_X1 _49761_ (.A1(_21452_),
    .A2(_11193_),
    .A3(_21316_),
    .A4(_21360_),
    .ZN(_21464_));
 INV_X1 _49762_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2984]),
    .ZN(_21465_));
 OAI21_X1 _49763_ (.A(_21464_),
    .B1(_21444_),
    .B2(_21465_),
    .ZN(_03025_));
 MUX2_X1 _49764_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2985]),
    .B(_21366_),
    .S(_21443_),
    .Z(_03026_));
 MUX2_X1 _49765_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2986]),
    .B(_21370_),
    .S(_21443_),
    .Z(_03027_));
 MUX2_X1 _49766_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2987]),
    .B(_21374_),
    .S(_21443_),
    .Z(_03028_));
 MUX2_X1 _49767_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2988]),
    .B(_21411_),
    .S(_21443_),
    .Z(_03029_));
 BUF_X8 _49768_ (.A(_10773_),
    .Z(_21466_));
 AND2_X4 _49769_ (.A1(_21466_),
    .A2(_21412_),
    .ZN(_21467_));
 BUF_X8 _49770_ (.A(_21467_),
    .Z(_21468_));
 BUF_X8 _49771_ (.A(_21468_),
    .Z(_21469_));
 MUX2_X1 _49772_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2891]),
    .B(_08524_),
    .S(_21469_),
    .Z(_02922_));
 MUX2_X1 _49773_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2892]),
    .B(_08529_),
    .S(_21469_),
    .Z(_02923_));
 MUX2_X1 _49774_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2893]),
    .B(_21295_),
    .S(_21469_),
    .Z(_02924_));
 MUX2_X1 _49775_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2894]),
    .B(_08537_),
    .S(_21469_),
    .Z(_02925_));
 MUX2_X1 _49776_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2895]),
    .B(_21298_),
    .S(_21469_),
    .Z(_02926_));
 BUF_X8 _49777_ (.A(_21467_),
    .Z(_21470_));
 MUX2_X1 _49778_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2896]),
    .B(_21300_),
    .S(_21470_),
    .Z(_02927_));
 MUX2_X1 _49779_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2897]),
    .B(_21302_),
    .S(_21470_),
    .Z(_02928_));
 MUX2_X1 _49780_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2898]),
    .B(_21304_),
    .S(_21470_),
    .Z(_02929_));
 MUX2_X1 _49781_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2899]),
    .B(_21306_),
    .S(_21470_),
    .Z(_02930_));
 NAND4_X2 _49782_ (.A1(_10782_),
    .A2(_21307_),
    .A3(_21429_),
    .A4(_21456_),
    .ZN(_21471_));
 INV_X4 _49783_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2900]),
    .ZN(_21472_));
 OAI21_X1 _49784_ (.A(_21471_),
    .B1(_21469_),
    .B2(_21472_),
    .ZN(_02933_));
 MUX2_X1 _49785_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2901]),
    .B(_21310_),
    .S(_21470_),
    .Z(_02934_));
 MUX2_X1 _49786_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2902]),
    .B(_21312_),
    .S(_21470_),
    .Z(_02935_));
 BUF_X8 _49787_ (.A(_08551_),
    .Z(_21473_));
 MUX2_X1 _49788_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2903]),
    .B(_21473_),
    .S(_21470_),
    .Z(_02936_));
 MUX2_X1 _49789_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2904]),
    .B(_10528_),
    .S(_21470_),
    .Z(_02937_));
 NAND4_X1 _49790_ (.A1(_10782_),
    .A2(_10570_),
    .A3(_21429_),
    .A4(_21456_),
    .ZN(_21474_));
 INV_X2 _49791_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2905]),
    .ZN(_21475_));
 OAI21_X1 _49792_ (.A(_21474_),
    .B1(_21469_),
    .B2(_21475_),
    .ZN(_02938_));
 BUF_X4 _49793_ (.A(_08561_),
    .Z(_21476_));
 MUX2_X1 _49794_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2906]),
    .B(_21476_),
    .S(_21470_),
    .Z(_02939_));
 BUF_X8 _49795_ (.A(_08564_),
    .Z(_21477_));
 MUX2_X1 _49796_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2907]),
    .B(_21477_),
    .S(_21470_),
    .Z(_02940_));
 BUF_X8 _49797_ (.A(_21467_),
    .Z(_21478_));
 MUX2_X1 _49798_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2908]),
    .B(_10532_),
    .S(_21478_),
    .Z(_02941_));
 BUF_X8 _49799_ (.A(_08571_),
    .Z(_21479_));
 MUX2_X1 _49800_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2909]),
    .B(_21479_),
    .S(_21478_),
    .Z(_02942_));
 BUF_X4 _49801_ (.A(_08575_),
    .Z(_21480_));
 MUX2_X1 _49802_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2910]),
    .B(_21480_),
    .S(_21478_),
    .Z(_02944_));
 BUF_X8 _49803_ (.A(_08578_),
    .Z(_21481_));
 MUX2_X1 _49804_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2911]),
    .B(_21481_),
    .S(_21478_),
    .Z(_02945_));
 BUF_X4 _49805_ (.A(_08581_),
    .Z(_21482_));
 MUX2_X1 _49806_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2912]),
    .B(_21482_),
    .S(_21478_),
    .Z(_02946_));
 BUF_X4 _49807_ (.A(_08584_),
    .Z(_21483_));
 MUX2_X1 _49808_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2913]),
    .B(_21483_),
    .S(_21478_),
    .Z(_02947_));
 MUX2_X1 _49809_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2914]),
    .B(_10539_),
    .S(_21478_),
    .Z(_02948_));
 BUF_X8 _49810_ (.A(_08591_),
    .Z(_21484_));
 MUX2_X1 _49811_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2915]),
    .B(_21484_),
    .S(_21478_),
    .Z(_02949_));
 MUX2_X1 _49812_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2916]),
    .B(_10541_),
    .S(_21478_),
    .Z(_02950_));
 BUF_X4 _49813_ (.A(_08597_),
    .Z(_21485_));
 MUX2_X1 _49814_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2917]),
    .B(_21485_),
    .S(_21478_),
    .Z(_02951_));
 BUF_X8 _49815_ (.A(_10781_),
    .Z(_21486_));
 NAND4_X1 _49816_ (.A1(_21486_),
    .A2(_10584_),
    .A3(_21429_),
    .A4(_21456_),
    .ZN(_21487_));
 INV_X1 _49817_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2918]),
    .ZN(_21488_));
 OAI21_X1 _49818_ (.A(_21487_),
    .B1(_21469_),
    .B2(_21488_),
    .ZN(_02952_));
 BUF_X16 _49819_ (.A(_21467_),
    .Z(_21489_));
 MUX2_X1 _49820_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2919]),
    .B(_10544_),
    .S(_21489_),
    .Z(_02953_));
 MUX2_X1 _49821_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2920]),
    .B(_10545_),
    .S(_21489_),
    .Z(_02955_));
 BUF_X8 _49822_ (.A(_08611_),
    .Z(_21490_));
 MUX2_X1 _49823_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2921]),
    .B(_21490_),
    .S(_21489_),
    .Z(_02956_));
 MUX2_X1 _49824_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2922]),
    .B(_10547_),
    .S(_21489_),
    .Z(_02957_));
 BUF_X8 _49825_ (.A(_08617_),
    .Z(_21491_));
 MUX2_X1 _49826_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2923]),
    .B(_21491_),
    .S(_21489_),
    .Z(_02958_));
 BUF_X4 _49827_ (.A(_08620_),
    .Z(_21492_));
 MUX2_X1 _49828_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2924]),
    .B(_21492_),
    .S(_21489_),
    .Z(_02959_));
 BUF_X4 _49829_ (.A(_21314_),
    .Z(_21493_));
 NAND4_X2 _49830_ (.A1(_21486_),
    .A2(_10591_),
    .A3(_21493_),
    .A4(_21456_),
    .ZN(_21494_));
 INV_X1 _49831_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2925]),
    .ZN(_21495_));
 OAI21_X1 _49832_ (.A(_21494_),
    .B1(_21469_),
    .B2(_21495_),
    .ZN(_02960_));
 BUF_X4 _49833_ (.A(_08626_),
    .Z(_21496_));
 MUX2_X1 _49834_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2926]),
    .B(_21496_),
    .S(_21489_),
    .Z(_02961_));
 BUF_X2 _49835_ (.A(_08629_),
    .Z(_21497_));
 MUX2_X1 _49836_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2927]),
    .B(_21497_),
    .S(_21489_),
    .Z(_02962_));
 MUX2_X1 _49837_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2928]),
    .B(_10553_),
    .S(_21489_),
    .Z(_02963_));
 BUF_X16 _49838_ (.A(_08635_),
    .Z(_21498_));
 MUX2_X1 _49839_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2929]),
    .B(_21498_),
    .S(_21489_),
    .Z(_02964_));
 MUX2_X1 _49840_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2930]),
    .B(_21340_),
    .S(_21468_),
    .Z(_02966_));
 MUX2_X1 _49841_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2931]),
    .B(_21344_),
    .S(_21468_),
    .Z(_02967_));
 BUF_X8 _49842_ (.A(_11015_),
    .Z(_21499_));
 NAND4_X1 _49843_ (.A1(_21486_),
    .A2(_21499_),
    .A3(_21316_),
    .A4(_21347_),
    .ZN(_21500_));
 INV_X4 _49844_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2932]),
    .ZN(_21501_));
 OAI21_X1 _49845_ (.A(_21500_),
    .B1(_21469_),
    .B2(_21501_),
    .ZN(_02968_));
 MUX2_X1 _49846_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2933]),
    .B(_21352_),
    .S(_21468_),
    .Z(_02969_));
 MUX2_X1 _49847_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2934]),
    .B(_21356_),
    .S(_21468_),
    .Z(_02970_));
 MUX2_X1 _49848_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2935]),
    .B(_21410_),
    .S(_21468_),
    .Z(_02971_));
 MUX2_X1 _49849_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2936]),
    .B(_21366_),
    .S(_21468_),
    .Z(_02972_));
 MUX2_X1 _49850_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2937]),
    .B(_21370_),
    .S(_21468_),
    .Z(_02973_));
 MUX2_X1 _49851_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2938]),
    .B(_21374_),
    .S(_21468_),
    .Z(_02974_));
 MUX2_X1 _49852_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2939]),
    .B(_21411_),
    .S(_21468_),
    .Z(_02975_));
 BUF_X8 _49853_ (.A(_10851_),
    .Z(_21502_));
 AND2_X4 _49854_ (.A1(_21502_),
    .A2(_21290_),
    .ZN(_21503_));
 BUF_X8 _49855_ (.A(_21503_),
    .Z(_21504_));
 MUX2_X1 _49856_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2842]),
    .B(_08524_),
    .S(_21504_),
    .Z(_02868_));
 MUX2_X1 _49857_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2843]),
    .B(_08529_),
    .S(_21504_),
    .Z(_02869_));
 MUX2_X1 _49858_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2844]),
    .B(_21295_),
    .S(_21504_),
    .Z(_02870_));
 MUX2_X1 _49859_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2845]),
    .B(_08537_),
    .S(_21504_),
    .Z(_02871_));
 MUX2_X1 _49860_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2846]),
    .B(_21298_),
    .S(_21504_),
    .Z(_02872_));
 MUX2_X1 _49861_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2847]),
    .B(_21300_),
    .S(_21504_),
    .Z(_02873_));
 MUX2_X1 _49862_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2848]),
    .B(_21302_),
    .S(_21504_),
    .Z(_02874_));
 MUX2_X1 _49863_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2849]),
    .B(_21304_),
    .S(_21504_),
    .Z(_02875_));
 MUX2_X1 _49864_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2850]),
    .B(_21306_),
    .S(_21504_),
    .Z(_02877_));
 BUF_X8 _49865_ (.A(_21503_),
    .Z(_21505_));
 MUX2_X1 _49866_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2851]),
    .B(_21308_),
    .S(_21505_),
    .Z(_02878_));
 MUX2_X1 _49867_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2852]),
    .B(_21310_),
    .S(_21505_),
    .Z(_02879_));
 BUF_X16 _49868_ (.A(_21311_),
    .Z(_21506_));
 NAND4_X1 _49869_ (.A1(_10860_),
    .A2(_21506_),
    .A3(_21493_),
    .A4(_21456_),
    .ZN(_21507_));
 BUF_X4 _49870_ (.A(_21504_),
    .Z(_21508_));
 INV_X1 _49871_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2853]),
    .ZN(_21509_));
 OAI21_X1 _49872_ (.A(_21507_),
    .B1(_21508_),
    .B2(_21509_),
    .ZN(_02880_));
 NAND4_X1 _49873_ (.A1(_10860_),
    .A2(_10563_),
    .A3(_21493_),
    .A4(_21456_),
    .ZN(_21510_));
 INV_X1 _49874_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2854]),
    .ZN(_21511_));
 OAI21_X1 _49875_ (.A(_21510_),
    .B1(_21508_),
    .B2(_21511_),
    .ZN(_02881_));
 MUX2_X1 _49876_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2855]),
    .B(_10528_),
    .S(_21505_),
    .Z(_02882_));
 BUF_X8 _49877_ (.A(_08558_),
    .Z(_21512_));
 MUX2_X1 _49878_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2856]),
    .B(_21512_),
    .S(_21505_),
    .Z(_02883_));
 MUX2_X1 _49879_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2857]),
    .B(_21476_),
    .S(_21505_),
    .Z(_02884_));
 BUF_X4 _49880_ (.A(_10859_),
    .Z(_21513_));
 NAND4_X2 _49881_ (.A1(_21513_),
    .A2(_10572_),
    .A3(_21493_),
    .A4(_21456_),
    .ZN(_21514_));
 INV_X1 _49882_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2858]),
    .ZN(_21515_));
 OAI21_X1 _49883_ (.A(_21514_),
    .B1(_21508_),
    .B2(_21515_),
    .ZN(_02885_));
 BUF_X8 _49884_ (.A(_08567_),
    .Z(_21516_));
 MUX2_X1 _49885_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2859]),
    .B(_21516_),
    .S(_21505_),
    .Z(_02886_));
 NAND4_X1 _49886_ (.A1(_21513_),
    .A2(_10600_),
    .A3(_21493_),
    .A4(_21456_),
    .ZN(_21517_));
 INV_X1 _49887_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2860]),
    .ZN(_21518_));
 OAI21_X1 _49888_ (.A(_21517_),
    .B1(_21508_),
    .B2(_21518_),
    .ZN(_02888_));
 MUX2_X1 _49889_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2861]),
    .B(_21480_),
    .S(_21505_),
    .Z(_02889_));
 MUX2_X1 _49890_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2862]),
    .B(_21481_),
    .S(_21505_),
    .Z(_02890_));
 MUX2_X1 _49891_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2863]),
    .B(_21482_),
    .S(_21505_),
    .Z(_02891_));
 MUX2_X1 _49892_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2864]),
    .B(_21483_),
    .S(_21505_),
    .Z(_02892_));
 BUF_X8 _49893_ (.A(_21503_),
    .Z(_21519_));
 MUX2_X1 _49894_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2865]),
    .B(_10539_),
    .S(_21519_),
    .Z(_02893_));
 MUX2_X1 _49895_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2866]),
    .B(_21484_),
    .S(_21519_),
    .Z(_02894_));
 MUX2_X1 _49896_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2867]),
    .B(_10541_),
    .S(_21519_),
    .Z(_02895_));
 MUX2_X1 _49897_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2868]),
    .B(_21485_),
    .S(_21519_),
    .Z(_02896_));
 BUF_X16 _49898_ (.A(_08600_),
    .Z(_21520_));
 BUF_X4 _49899_ (.A(_10791_),
    .Z(_21521_));
 NAND4_X1 _49900_ (.A1(_21513_),
    .A2(_21520_),
    .A3(_21493_),
    .A4(_21521_),
    .ZN(_21522_));
 INV_X1 _49901_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2869]),
    .ZN(_21523_));
 OAI21_X1 _49902_ (.A(_21522_),
    .B1(_21508_),
    .B2(_21523_),
    .ZN(_02897_));
 MUX2_X1 _49903_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2870]),
    .B(_10544_),
    .S(_21519_),
    .Z(_02899_));
 NAND4_X1 _49904_ (.A1(_21513_),
    .A2(_10616_),
    .A3(_21493_),
    .A4(_21521_),
    .ZN(_21524_));
 INV_X1 _49905_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2871]),
    .ZN(_21525_));
 OAI21_X1 _49906_ (.A(_21524_),
    .B1(_21508_),
    .B2(_21525_),
    .ZN(_02900_));
 NAND4_X1 _49907_ (.A1(_21513_),
    .A2(_10587_),
    .A3(_21493_),
    .A4(_21521_),
    .ZN(_21526_));
 INV_X1 _49908_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2872]),
    .ZN(_21527_));
 OAI21_X1 _49909_ (.A(_21526_),
    .B1(_21508_),
    .B2(_21527_),
    .ZN(_02901_));
 NAND4_X1 _49910_ (.A1(_21513_),
    .A2(_10588_),
    .A3(_21493_),
    .A4(_21521_),
    .ZN(_21528_));
 INV_X1 _49911_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2873]),
    .ZN(_21529_));
 OAI21_X1 _49912_ (.A(_21528_),
    .B1(_21508_),
    .B2(_21529_),
    .ZN(_02902_));
 MUX2_X1 _49913_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2874]),
    .B(_21491_),
    .S(_21519_),
    .Z(_02903_));
 MUX2_X1 _49914_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2875]),
    .B(_21492_),
    .S(_21519_),
    .Z(_02904_));
 MUX2_X1 _49915_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2876]),
    .B(_10550_),
    .S(_21519_),
    .Z(_02905_));
 MUX2_X1 _49916_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2877]),
    .B(_21496_),
    .S(_21519_),
    .Z(_02906_));
 MUX2_X1 _49917_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2878]),
    .B(_21497_),
    .S(_21519_),
    .Z(_02907_));
 BUF_X8 _49918_ (.A(_21503_),
    .Z(_21530_));
 MUX2_X1 _49919_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2879]),
    .B(_10553_),
    .S(_21530_),
    .Z(_02908_));
 NAND4_X1 _49920_ (.A1(_21513_),
    .A2(_10595_),
    .A3(_21493_),
    .A4(_21521_),
    .ZN(_21531_));
 INV_X2 _49921_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2880]),
    .ZN(_21532_));
 OAI21_X1 _49922_ (.A(_21531_),
    .B1(_21508_),
    .B2(_21532_),
    .ZN(_02910_));
 MUX2_X1 _49923_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2881]),
    .B(_21340_),
    .S(_21530_),
    .Z(_02911_));
 MUX2_X1 _49924_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2882]),
    .B(_21344_),
    .S(_21530_),
    .Z(_02912_));
 MUX2_X1 _49925_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2883]),
    .B(_21348_),
    .S(_21530_),
    .Z(_02913_));
 MUX2_X1 _49926_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2884]),
    .B(_21352_),
    .S(_21530_),
    .Z(_02914_));
 BUF_X16 _49927_ (.A(_21355_),
    .Z(_21533_));
 NAND4_X1 _49928_ (.A1(_21513_),
    .A2(_21499_),
    .A3(_21316_),
    .A4(_21533_),
    .ZN(_21534_));
 INV_X1 _49929_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2885]),
    .ZN(_21535_));
 OAI21_X1 _49930_ (.A(_21534_),
    .B1(_21508_),
    .B2(_21535_),
    .ZN(_02915_));
 MUX2_X1 _49931_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2886]),
    .B(_21410_),
    .S(_21530_),
    .Z(_02916_));
 MUX2_X1 _49932_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2887]),
    .B(_21366_),
    .S(_21530_),
    .Z(_02917_));
 MUX2_X1 _49933_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2888]),
    .B(_21370_),
    .S(_21530_),
    .Z(_02918_));
 MUX2_X1 _49934_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2889]),
    .B(_21374_),
    .S(_21530_),
    .Z(_02919_));
 MUX2_X1 _49935_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2890]),
    .B(_21411_),
    .S(_21530_),
    .Z(_02921_));
 BUF_X8 _49936_ (.A(_10863_),
    .Z(_21536_));
 AND2_X4 _49937_ (.A1(_21536_),
    .A2(_10784_),
    .ZN(_21537_));
 BUF_X8 _49938_ (.A(_21537_),
    .Z(_21538_));
 MUX2_X1 _49939_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2793]),
    .B(_08524_),
    .S(_21538_),
    .Z(_02813_));
 MUX2_X1 _49940_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2794]),
    .B(_08529_),
    .S(_21538_),
    .Z(_02814_));
 MUX2_X1 _49941_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2795]),
    .B(_21295_),
    .S(_21538_),
    .Z(_02815_));
 MUX2_X1 _49942_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2796]),
    .B(_08537_),
    .S(_21538_),
    .Z(_02816_));
 MUX2_X1 _49943_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2797]),
    .B(_21298_),
    .S(_21538_),
    .Z(_02817_));
 MUX2_X1 _49944_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2798]),
    .B(_21300_),
    .S(_21538_),
    .Z(_02818_));
 MUX2_X1 _49945_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2799]),
    .B(_21302_),
    .S(_21538_),
    .Z(_02819_));
 MUX2_X1 _49946_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2800]),
    .B(_21304_),
    .S(_21538_),
    .Z(_02822_));
 BUF_X8 _49947_ (.A(_21537_),
    .Z(_21539_));
 MUX2_X1 _49948_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2801]),
    .B(_21306_),
    .S(_21539_),
    .Z(_02823_));
 MUX2_X1 _49949_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2802]),
    .B(_21308_),
    .S(_21539_),
    .Z(_02824_));
 MUX2_X1 _49950_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2803]),
    .B(_21310_),
    .S(_21539_),
    .Z(_02825_));
 BUF_X4 _49951_ (.A(_21314_),
    .Z(_21540_));
 NAND4_X1 _49952_ (.A1(_10870_),
    .A2(_21506_),
    .A3(_21540_),
    .A4(_21521_),
    .ZN(_21541_));
 BUF_X4 _49953_ (.A(_21538_),
    .Z(_21542_));
 INV_X1 _49954_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2804]),
    .ZN(_21543_));
 OAI21_X1 _49955_ (.A(_21541_),
    .B1(_21542_),
    .B2(_21543_),
    .ZN(_02826_));
 NAND4_X1 _49956_ (.A1(_10870_),
    .A2(_10563_),
    .A3(_21540_),
    .A4(_21521_),
    .ZN(_21544_));
 INV_X1 _49957_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2805]),
    .ZN(_21545_));
 OAI21_X1 _49958_ (.A(_21544_),
    .B1(_21542_),
    .B2(_21545_),
    .ZN(_02827_));
 BUF_X8 _49959_ (.A(_10869_),
    .Z(_21546_));
 NAND4_X1 _49960_ (.A1(_21546_),
    .A2(_10569_),
    .A3(_21540_),
    .A4(_21521_),
    .ZN(_21547_));
 INV_X1 _49961_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2806]),
    .ZN(_21548_));
 OAI21_X1 _49962_ (.A(_21547_),
    .B1(_21542_),
    .B2(_21548_),
    .ZN(_02828_));
 MUX2_X1 _49963_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2807]),
    .B(_21512_),
    .S(_21539_),
    .Z(_02829_));
 MUX2_X1 _49964_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2808]),
    .B(_21476_),
    .S(_21539_),
    .Z(_02830_));
 MUX2_X1 _49965_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2809]),
    .B(_21477_),
    .S(_21539_),
    .Z(_02831_));
 MUX2_X1 _49966_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2810]),
    .B(_21516_),
    .S(_21539_),
    .Z(_02833_));
 MUX2_X1 _49967_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2811]),
    .B(_21479_),
    .S(_21539_),
    .Z(_02834_));
 MUX2_X1 _49968_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2812]),
    .B(_21480_),
    .S(_21539_),
    .Z(_02835_));
 MUX2_X1 _49969_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2813]),
    .B(_21481_),
    .S(_21539_),
    .Z(_02836_));
 BUF_X16 _49970_ (.A(_21537_),
    .Z(_21549_));
 MUX2_X1 _49971_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2814]),
    .B(_21482_),
    .S(_21549_),
    .Z(_02837_));
 MUX2_X1 _49972_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2815]),
    .B(_21483_),
    .S(_21549_),
    .Z(_02838_));
 NAND4_X1 _49973_ (.A1(_21546_),
    .A2(_10580_),
    .A3(_21540_),
    .A4(_21521_),
    .ZN(_21550_));
 INV_X1 _49974_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2816]),
    .ZN(_21551_));
 OAI21_X1 _49975_ (.A(_21550_),
    .B1(_21542_),
    .B2(_21551_),
    .ZN(_02839_));
 MUX2_X1 _49976_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2817]),
    .B(_21484_),
    .S(_21549_),
    .Z(_02840_));
 NAND4_X1 _49977_ (.A1(_21546_),
    .A2(_10582_),
    .A3(_21540_),
    .A4(_21521_),
    .ZN(_21552_));
 INV_X1 _49978_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2818]),
    .ZN(_21553_));
 OAI21_X1 _49979_ (.A(_21552_),
    .B1(_21542_),
    .B2(_21553_),
    .ZN(_02841_));
 MUX2_X1 _49980_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2819]),
    .B(_21485_),
    .S(_21549_),
    .Z(_02842_));
 BUF_X8 _49981_ (.A(_08600_),
    .Z(_21554_));
 MUX2_X1 _49982_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2820]),
    .B(_21554_),
    .S(_21549_),
    .Z(_02844_));
 BUF_X8 _49983_ (.A(_08604_),
    .Z(_21555_));
 MUX2_X1 _49984_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2821]),
    .B(_21555_),
    .S(_21549_),
    .Z(_02845_));
 NAND4_X1 _49985_ (.A1(_21546_),
    .A2(_10616_),
    .A3(_21540_),
    .A4(_10791_),
    .ZN(_21556_));
 INV_X1 _49986_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2822]),
    .ZN(_21557_));
 OAI21_X1 _49987_ (.A(_21556_),
    .B1(_21542_),
    .B2(_21557_),
    .ZN(_02846_));
 BUF_X16 _49988_ (.A(_08611_),
    .Z(_21558_));
 NAND4_X1 _49989_ (.A1(_21546_),
    .A2(_21558_),
    .A3(_21540_),
    .A4(_10791_),
    .ZN(_21559_));
 INV_X1 _49990_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2823]),
    .ZN(_21560_));
 OAI21_X1 _49991_ (.A(_21559_),
    .B1(_21542_),
    .B2(_21560_),
    .ZN(_02847_));
 BUF_X8 _49992_ (.A(_08614_),
    .Z(_21561_));
 MUX2_X1 _49993_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2824]),
    .B(_21561_),
    .S(_21549_),
    .Z(_02848_));
 MUX2_X1 _49994_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2825]),
    .B(_21491_),
    .S(_21549_),
    .Z(_02849_));
 MUX2_X1 _49995_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2826]),
    .B(_21492_),
    .S(_21549_),
    .Z(_02850_));
 BUF_X32 _49996_ (.A(_08623_),
    .Z(_21562_));
 NAND4_X1 _49997_ (.A1(_21546_),
    .A2(_21562_),
    .A3(_21540_),
    .A4(_10791_),
    .ZN(_21563_));
 INV_X1 _49998_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2827]),
    .ZN(_21564_));
 OAI21_X1 _49999_ (.A(_21563_),
    .B1(_21542_),
    .B2(_21564_),
    .ZN(_02851_));
 MUX2_X1 _50000_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2828]),
    .B(_21496_),
    .S(_21549_),
    .Z(_02852_));
 BUF_X8 _50001_ (.A(_21537_),
    .Z(_21565_));
 MUX2_X1 _50002_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2829]),
    .B(_21497_),
    .S(_21565_),
    .Z(_02853_));
 BUF_X8 _50003_ (.A(_08632_),
    .Z(_21566_));
 MUX2_X1 _50004_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2830]),
    .B(_21566_),
    .S(_21565_),
    .Z(_02855_));
 MUX2_X1 _50005_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2831]),
    .B(_21498_),
    .S(_21565_),
    .Z(_02856_));
 MUX2_X1 _50006_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2832]),
    .B(_21340_),
    .S(_21565_),
    .Z(_02857_));
 MUX2_X1 _50007_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2833]),
    .B(_21344_),
    .S(_21565_),
    .Z(_02858_));
 MUX2_X1 _50008_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2834]),
    .B(_21348_),
    .S(_21565_),
    .Z(_02859_));
 MUX2_X1 _50009_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2835]),
    .B(_21352_),
    .S(_21565_),
    .Z(_02860_));
 NAND4_X1 _50010_ (.A1(_21546_),
    .A2(_21499_),
    .A3(_21316_),
    .A4(_21533_),
    .ZN(_21567_));
 INV_X1 _50011_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2836]),
    .ZN(_21568_));
 OAI21_X1 _50012_ (.A(_21567_),
    .B1(_21542_),
    .B2(_21568_),
    .ZN(_02861_));
 MUX2_X1 _50013_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2837]),
    .B(_21410_),
    .S(_21565_),
    .Z(_02862_));
 MUX2_X1 _50014_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2838]),
    .B(_21366_),
    .S(_21565_),
    .Z(_02863_));
 NAND4_X1 _50015_ (.A1(_21546_),
    .A2(_21499_),
    .A3(_21316_),
    .A4(_21369_),
    .ZN(_21569_));
 INV_X1 _50016_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2839]),
    .ZN(_21570_));
 OAI21_X1 _50017_ (.A(_21569_),
    .B1(_21542_),
    .B2(_21570_),
    .ZN(_02864_));
 MUX2_X1 _50018_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2840]),
    .B(_21374_),
    .S(_21565_),
    .Z(_02866_));
 NAND4_X2 _50019_ (.A1(_21546_),
    .A2(_21499_),
    .A3(_21316_),
    .A4(_21377_),
    .ZN(_21571_));
 INV_X1 _50020_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2841]),
    .ZN(_21572_));
 OAI21_X1 _50021_ (.A(_21571_),
    .B1(_21538_),
    .B2(_21572_),
    .ZN(_02867_));
 BUF_X8 _50022_ (.A(_10887_),
    .Z(_21573_));
 BUF_X32 _50023_ (.A(_10762_),
    .Z(_21574_));
 AND2_X4 _50024_ (.A1(_21573_),
    .A2(_21574_),
    .ZN(_21575_));
 BUF_X16 _50025_ (.A(_21575_),
    .Z(_21576_));
 BUF_X8 _50026_ (.A(_21576_),
    .Z(_21577_));
 MUX2_X1 _50027_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2695]),
    .B(_08524_),
    .S(_21577_),
    .Z(_02704_));
 MUX2_X1 _50028_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2696]),
    .B(_08529_),
    .S(_21577_),
    .Z(_02705_));
 MUX2_X1 _50029_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2697]),
    .B(_21295_),
    .S(_21577_),
    .Z(_02706_));
 MUX2_X1 _50030_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2698]),
    .B(_08537_),
    .S(_21577_),
    .Z(_02707_));
 MUX2_X1 _50031_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2699]),
    .B(_21298_),
    .S(_21577_),
    .Z(_02708_));
 MUX2_X1 _50032_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2700]),
    .B(_21300_),
    .S(_21577_),
    .Z(_02711_));
 BUF_X16 _50033_ (.A(_21301_),
    .Z(_21578_));
 BUF_X8 _50034_ (.A(_10893_),
    .Z(_21579_));
 NAND4_X1 _50035_ (.A1(_21391_),
    .A2(_21578_),
    .A3(_21540_),
    .A4(_21579_),
    .ZN(_21580_));
 INV_X1 _50036_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2701]),
    .ZN(_21581_));
 OAI21_X1 _50037_ (.A(_21580_),
    .B1(_21577_),
    .B2(_21581_),
    .ZN(_02712_));
 BUF_X32 _50038_ (.A(_21303_),
    .Z(_21582_));
 NAND4_X2 _50039_ (.A1(_21391_),
    .A2(_21582_),
    .A3(_21540_),
    .A4(_21579_),
    .ZN(_21583_));
 INV_X1 _50040_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2702]),
    .ZN(_21584_));
 OAI21_X1 _50041_ (.A(_21583_),
    .B1(_21577_),
    .B2(_21584_),
    .ZN(_02713_));
 BUF_X8 _50042_ (.A(_21575_),
    .Z(_21585_));
 MUX2_X1 _50043_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2703]),
    .B(_21306_),
    .S(_21585_),
    .Z(_02714_));
 MUX2_X1 _50044_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2704]),
    .B(_21308_),
    .S(_21585_),
    .Z(_02715_));
 MUX2_X1 _50045_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2705]),
    .B(_21310_),
    .S(_21585_),
    .Z(_02716_));
 MUX2_X1 _50046_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2706]),
    .B(_21312_),
    .S(_21585_),
    .Z(_02717_));
 MUX2_X1 _50047_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2707]),
    .B(_21473_),
    .S(_21585_),
    .Z(_02718_));
 BUF_X4 _50048_ (.A(_08555_),
    .Z(_21586_));
 MUX2_X1 _50049_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2708]),
    .B(_21586_),
    .S(_21585_),
    .Z(_02719_));
 MUX2_X1 _50050_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2709]),
    .B(_21512_),
    .S(_21585_),
    .Z(_02720_));
 MUX2_X1 _50051_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2710]),
    .B(_21476_),
    .S(_21585_),
    .Z(_02722_));
 MUX2_X1 _50052_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2711]),
    .B(_21477_),
    .S(_21585_),
    .Z(_02723_));
 MUX2_X1 _50053_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2712]),
    .B(_21516_),
    .S(_21585_),
    .Z(_02724_));
 BUF_X16 _50054_ (.A(_21575_),
    .Z(_21587_));
 MUX2_X1 _50055_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2713]),
    .B(_21479_),
    .S(_21587_),
    .Z(_02725_));
 MUX2_X1 _50056_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2714]),
    .B(_21480_),
    .S(_21587_),
    .Z(_02726_));
 MUX2_X1 _50057_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2715]),
    .B(_21481_),
    .S(_21587_),
    .Z(_02727_));
 MUX2_X1 _50058_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2716]),
    .B(_21482_),
    .S(_21587_),
    .Z(_02728_));
 MUX2_X1 _50059_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2717]),
    .B(_21483_),
    .S(_21587_),
    .Z(_02729_));
 BUF_X8 _50060_ (.A(_08588_),
    .Z(_21588_));
 MUX2_X1 _50061_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2718]),
    .B(_21588_),
    .S(_21587_),
    .Z(_02730_));
 MUX2_X1 _50062_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2719]),
    .B(_21484_),
    .S(_21587_),
    .Z(_02731_));
 MUX2_X1 _50063_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2720]),
    .B(_10541_),
    .S(_21587_),
    .Z(_02733_));
 MUX2_X1 _50064_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2721]),
    .B(_21485_),
    .S(_21587_),
    .Z(_02734_));
 MUX2_X1 _50065_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2722]),
    .B(_21554_),
    .S(_21587_),
    .Z(_02735_));
 BUF_X8 _50066_ (.A(_21575_),
    .Z(_21589_));
 MUX2_X1 _50067_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2723]),
    .B(_21555_),
    .S(_21589_),
    .Z(_02736_));
 BUF_X4 _50068_ (.A(_08608_),
    .Z(_21590_));
 MUX2_X1 _50069_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2724]),
    .B(_21590_),
    .S(_21589_),
    .Z(_02737_));
 MUX2_X1 _50070_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2725]),
    .B(_21490_),
    .S(_21589_),
    .Z(_02738_));
 MUX2_X1 _50071_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2726]),
    .B(_21561_),
    .S(_21589_),
    .Z(_02739_));
 MUX2_X1 _50072_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2727]),
    .B(_21491_),
    .S(_21589_),
    .Z(_02740_));
 MUX2_X1 _50073_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2728]),
    .B(_21492_),
    .S(_21589_),
    .Z(_02741_));
 MUX2_X1 _50074_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2729]),
    .B(_10550_),
    .S(_21589_),
    .Z(_02742_));
 MUX2_X1 _50075_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2730]),
    .B(_21496_),
    .S(_21589_),
    .Z(_02744_));
 MUX2_X1 _50076_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2731]),
    .B(_21497_),
    .S(_21589_),
    .Z(_02745_));
 MUX2_X1 _50077_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2732]),
    .B(_21566_),
    .S(_21589_),
    .Z(_02746_));
 BUF_X32 _50078_ (.A(_08635_),
    .Z(_21591_));
 BUF_X8 _50079_ (.A(_21314_),
    .Z(_21592_));
 NAND4_X1 _50080_ (.A1(_21391_),
    .A2(_21591_),
    .A3(_21592_),
    .A4(_21579_),
    .ZN(_21593_));
 INV_X2 _50081_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2733]),
    .ZN(_21594_));
 OAI21_X1 _50082_ (.A(_21593_),
    .B1(_21577_),
    .B2(_21594_),
    .ZN(_02747_));
 BUF_X16 _50083_ (.A(_21339_),
    .Z(_21595_));
 NAND4_X1 _50084_ (.A1(_21391_),
    .A2(_21499_),
    .A3(_10894_),
    .A4(_21595_),
    .ZN(_21596_));
 INV_X1 _50085_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2734]),
    .ZN(_21597_));
 OAI21_X1 _50086_ (.A(_21596_),
    .B1(_21577_),
    .B2(_21597_),
    .ZN(_02748_));
 MUX2_X1 _50087_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2735]),
    .B(_21344_),
    .S(_21576_),
    .Z(_02749_));
 MUX2_X1 _50088_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2736]),
    .B(_21348_),
    .S(_21576_),
    .Z(_02750_));
 MUX2_X1 _50089_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2737]),
    .B(_21352_),
    .S(_21576_),
    .Z(_02751_));
 MUX2_X1 _50090_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2738]),
    .B(_21356_),
    .S(_21576_),
    .Z(_02752_));
 MUX2_X1 _50091_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2739]),
    .B(_21410_),
    .S(_21576_),
    .Z(_02753_));
 MUX2_X1 _50092_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2740]),
    .B(_21366_),
    .S(_21576_),
    .Z(_02755_));
 MUX2_X1 _50093_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2741]),
    .B(_21370_),
    .S(_21576_),
    .Z(_02756_));
 MUX2_X1 _50094_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2742]),
    .B(_21374_),
    .S(_21576_),
    .Z(_02757_));
 MUX2_X1 _50095_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2743]),
    .B(_21411_),
    .S(_21576_),
    .Z(_02758_));
 BUF_X32 _50096_ (.A(fe_cmd_i[34]),
    .Z(_21598_));
 BUF_X8 _50097_ (.A(_21598_),
    .Z(_21599_));
 BUF_X8 _50098_ (.A(_10896_),
    .Z(_21600_));
 BUF_X8 _50099_ (.A(_21600_),
    .Z(_21601_));
 AND2_X4 _50100_ (.A1(_21601_),
    .A2(_21290_),
    .ZN(_21602_));
 BUF_X16 _50101_ (.A(_21602_),
    .Z(_21603_));
 BUF_X8 _50102_ (.A(_21603_),
    .Z(_21604_));
 MUX2_X1 _50103_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2646]),
    .B(_21599_),
    .S(_21604_),
    .Z(_02650_));
 BUF_X32 _50104_ (.A(fe_cmd_i[35]),
    .Z(_21605_));
 BUF_X8 _50105_ (.A(_21605_),
    .Z(_21606_));
 MUX2_X1 _50106_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2647]),
    .B(_21606_),
    .S(_21604_),
    .Z(_02651_));
 BUF_X16 _50107_ (.A(_21602_),
    .Z(_21607_));
 MUX2_X1 _50108_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2648]),
    .B(_21295_),
    .S(_21607_),
    .Z(_02652_));
 BUF_X32 _50109_ (.A(fe_cmd_i[37]),
    .Z(_21608_));
 BUF_X8 _50110_ (.A(_21608_),
    .Z(_21609_));
 MUX2_X1 _50111_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2649]),
    .B(_21609_),
    .S(_21607_),
    .Z(_02653_));
 MUX2_X1 _50112_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2650]),
    .B(_21298_),
    .S(_21607_),
    .Z(_02655_));
 MUX2_X1 _50113_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2651]),
    .B(_21300_),
    .S(_21607_),
    .Z(_02656_));
 NAND4_X1 _50114_ (.A1(_21422_),
    .A2(_21578_),
    .A3(_21592_),
    .A4(_21579_),
    .ZN(_21610_));
 INV_X1 _50115_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2652]),
    .ZN(_21611_));
 OAI21_X1 _50116_ (.A(_21610_),
    .B1(_21604_),
    .B2(_21611_),
    .ZN(_02657_));
 NAND4_X1 _50117_ (.A1(_21422_),
    .A2(_21582_),
    .A3(_21592_),
    .A4(_21579_),
    .ZN(_21612_));
 INV_X1 _50118_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2653]),
    .ZN(_21613_));
 OAI21_X1 _50119_ (.A(_21612_),
    .B1(_21604_),
    .B2(_21613_),
    .ZN(_02658_));
 MUX2_X1 _50120_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2654]),
    .B(_21306_),
    .S(_21607_),
    .Z(_02659_));
 NAND4_X1 _50121_ (.A1(_21422_),
    .A2(_21307_),
    .A3(_21592_),
    .A4(_21579_),
    .ZN(_21614_));
 INV_X1 _50122_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2655]),
    .ZN(_21615_));
 OAI21_X1 _50123_ (.A(_21614_),
    .B1(_21604_),
    .B2(_21615_),
    .ZN(_02660_));
 MUX2_X1 _50124_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2656]),
    .B(_21310_),
    .S(_21607_),
    .Z(_02661_));
 MUX2_X1 _50125_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2657]),
    .B(_21312_),
    .S(_21607_),
    .Z(_02662_));
 MUX2_X1 _50126_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2658]),
    .B(_21473_),
    .S(_21607_),
    .Z(_02663_));
 MUX2_X1 _50127_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2659]),
    .B(_21586_),
    .S(_21607_),
    .Z(_02664_));
 MUX2_X1 _50128_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2660]),
    .B(_21512_),
    .S(_21607_),
    .Z(_02666_));
 BUF_X8 _50129_ (.A(_21602_),
    .Z(_21616_));
 MUX2_X1 _50130_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2661]),
    .B(_21476_),
    .S(_21616_),
    .Z(_02667_));
 MUX2_X1 _50131_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2662]),
    .B(_21477_),
    .S(_21616_),
    .Z(_02668_));
 MUX2_X1 _50132_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2663]),
    .B(_21516_),
    .S(_21616_),
    .Z(_02669_));
 MUX2_X1 _50133_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2664]),
    .B(_21479_),
    .S(_21616_),
    .Z(_02670_));
 MUX2_X1 _50134_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2665]),
    .B(_21480_),
    .S(_21616_),
    .Z(_02671_));
 MUX2_X1 _50135_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2666]),
    .B(_21481_),
    .S(_21616_),
    .Z(_02672_));
 MUX2_X1 _50136_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2667]),
    .B(_21482_),
    .S(_21616_),
    .Z(_02673_));
 MUX2_X1 _50137_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2668]),
    .B(_21483_),
    .S(_21616_),
    .Z(_02674_));
 MUX2_X1 _50138_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2669]),
    .B(_21588_),
    .S(_21616_),
    .Z(_02675_));
 MUX2_X1 _50139_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2670]),
    .B(_21484_),
    .S(_21616_),
    .Z(_02677_));
 BUF_X8 _50140_ (.A(_08594_),
    .Z(_21617_));
 BUF_X16 _50141_ (.A(_21602_),
    .Z(_21618_));
 MUX2_X1 _50142_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2671]),
    .B(_21617_),
    .S(_21618_),
    .Z(_02678_));
 MUX2_X1 _50143_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2672]),
    .B(_21485_),
    .S(_21618_),
    .Z(_02679_));
 MUX2_X1 _50144_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2673]),
    .B(_21554_),
    .S(_21618_),
    .Z(_02680_));
 MUX2_X1 _50145_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2674]),
    .B(_21555_),
    .S(_21618_),
    .Z(_02681_));
 MUX2_X1 _50146_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2675]),
    .B(_21590_),
    .S(_21618_),
    .Z(_02682_));
 NAND4_X1 _50147_ (.A1(_21422_),
    .A2(_21558_),
    .A3(_21592_),
    .A4(_21579_),
    .ZN(_21619_));
 INV_X1 _50148_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2676]),
    .ZN(_21620_));
 OAI21_X1 _50149_ (.A(_21619_),
    .B1(_21604_),
    .B2(_21620_),
    .ZN(_02683_));
 MUX2_X1 _50150_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2677]),
    .B(_21561_),
    .S(_21618_),
    .Z(_02684_));
 MUX2_X1 _50151_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2678]),
    .B(_21491_),
    .S(_21618_),
    .Z(_02685_));
 MUX2_X1 _50152_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2679]),
    .B(_21492_),
    .S(_21618_),
    .Z(_02686_));
 BUF_X8 _50153_ (.A(_08623_),
    .Z(_21621_));
 MUX2_X1 _50154_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2680]),
    .B(_21621_),
    .S(_21618_),
    .Z(_02688_));
 MUX2_X1 _50155_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2681]),
    .B(_21496_),
    .S(_21618_),
    .Z(_02689_));
 MUX2_X1 _50156_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2682]),
    .B(_21497_),
    .S(_21603_),
    .Z(_02690_));
 MUX2_X1 _50157_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2683]),
    .B(_21566_),
    .S(_21603_),
    .Z(_02691_));
 NAND4_X2 _50158_ (.A1(_21422_),
    .A2(_21591_),
    .A3(_21592_),
    .A4(_21579_),
    .ZN(_21622_));
 INV_X4 _50159_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2684]),
    .ZN(_21623_));
 OAI21_X1 _50160_ (.A(_21622_),
    .B1(_21604_),
    .B2(_21623_),
    .ZN(_02692_));
 NAND4_X1 _50161_ (.A1(_21422_),
    .A2(_21499_),
    .A3(_10894_),
    .A4(_21595_),
    .ZN(_21624_));
 INV_X1 _50162_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2685]),
    .ZN(_21625_));
 OAI21_X1 _50163_ (.A(_21624_),
    .B1(_21604_),
    .B2(_21625_),
    .ZN(_02693_));
 MUX2_X1 _50164_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2686]),
    .B(_21344_),
    .S(_21603_),
    .Z(_02694_));
 BUF_X4 _50165_ (.A(_10893_),
    .Z(_21626_));
 NAND4_X1 _50166_ (.A1(_21422_),
    .A2(_21499_),
    .A3(_21626_),
    .A4(_21347_),
    .ZN(_21627_));
 INV_X1 _50167_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2687]),
    .ZN(_21628_));
 OAI21_X1 _50168_ (.A(_21627_),
    .B1(_21604_),
    .B2(_21628_),
    .ZN(_02695_));
 MUX2_X1 _50169_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2688]),
    .B(_21352_),
    .S(_21603_),
    .Z(_02696_));
 BUF_X8 _50170_ (.A(_10819_),
    .Z(_21629_));
 NAND4_X1 _50171_ (.A1(_21629_),
    .A2(_21499_),
    .A3(_21626_),
    .A4(_21533_),
    .ZN(_21630_));
 INV_X1 _50172_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2689]),
    .ZN(_21631_));
 OAI21_X1 _50173_ (.A(_21630_),
    .B1(_21604_),
    .B2(_21631_),
    .ZN(_02697_));
 MUX2_X1 _50174_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2690]),
    .B(_21410_),
    .S(_21603_),
    .Z(_02699_));
 MUX2_X1 _50175_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2691]),
    .B(_21366_),
    .S(_21603_),
    .Z(_02700_));
 MUX2_X1 _50176_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2692]),
    .B(_21370_),
    .S(_21603_),
    .Z(_02701_));
 MUX2_X1 _50177_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2693]),
    .B(_21374_),
    .S(_21603_),
    .Z(_02702_));
 MUX2_X1 _50178_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2694]),
    .B(_21411_),
    .S(_21603_),
    .Z(_02703_));
 AND2_X4 _50179_ (.A1(_10902_),
    .A2(_21412_),
    .ZN(_21632_));
 BUF_X16 _50180_ (.A(_21632_),
    .Z(_21633_));
 BUF_X8 _50181_ (.A(_21633_),
    .Z(_21634_));
 MUX2_X1 _50182_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2597]),
    .B(_21599_),
    .S(_21634_),
    .Z(_02595_));
 MUX2_X1 _50183_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2598]),
    .B(_21606_),
    .S(_21634_),
    .Z(_02596_));
 MUX2_X1 _50184_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2599]),
    .B(_21295_),
    .S(_21634_),
    .Z(_02597_));
 MUX2_X1 _50185_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2600]),
    .B(_21609_),
    .S(_21634_),
    .Z(_02600_));
 MUX2_X1 _50186_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2601]),
    .B(_21298_),
    .S(_21634_),
    .Z(_02601_));
 BUF_X4 _50187_ (.A(_21299_),
    .Z(_21635_));
 BUF_X8 _50188_ (.A(_21632_),
    .Z(_21636_));
 MUX2_X1 _50189_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2602]),
    .B(_21635_),
    .S(_21636_),
    .Z(_02602_));
 MUX2_X1 _50190_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2603]),
    .B(_21302_),
    .S(_21636_),
    .Z(_02603_));
 MUX2_X1 _50191_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2604]),
    .B(_21304_),
    .S(_21636_),
    .Z(_02604_));
 MUX2_X1 _50192_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2605]),
    .B(_21306_),
    .S(_21636_),
    .Z(_02605_));
 MUX2_X1 _50193_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2606]),
    .B(_21308_),
    .S(_21636_),
    .Z(_02606_));
 NAND4_X1 _50194_ (.A1(_10833_),
    .A2(_21446_),
    .A3(_21592_),
    .A4(_21579_),
    .ZN(_21637_));
 INV_X1 _50195_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2607]),
    .ZN(_21638_));
 OAI21_X1 _50196_ (.A(_21637_),
    .B1(_21634_),
    .B2(_21638_),
    .ZN(_02607_));
 MUX2_X1 _50197_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2608]),
    .B(_21312_),
    .S(_21636_),
    .Z(_02608_));
 MUX2_X1 _50198_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2609]),
    .B(_21473_),
    .S(_21636_),
    .Z(_02609_));
 MUX2_X1 _50199_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2610]),
    .B(_21586_),
    .S(_21636_),
    .Z(_02611_));
 MUX2_X1 _50200_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2611]),
    .B(_21512_),
    .S(_21636_),
    .Z(_02612_));
 MUX2_X1 _50201_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2612]),
    .B(_21476_),
    .S(_21636_),
    .Z(_02613_));
 BUF_X16 _50202_ (.A(_21632_),
    .Z(_21639_));
 MUX2_X1 _50203_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2613]),
    .B(_21477_),
    .S(_21639_),
    .Z(_02614_));
 BUF_X16 _50204_ (.A(_10832_),
    .Z(_21640_));
 BUF_X4 _50205_ (.A(_10893_),
    .Z(_21641_));
 NAND4_X1 _50206_ (.A1(_21640_),
    .A2(_10599_),
    .A3(_21592_),
    .A4(_21641_),
    .ZN(_21642_));
 INV_X1 _50207_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2614]),
    .ZN(_21643_));
 OAI21_X1 _50208_ (.A(_21642_),
    .B1(_21634_),
    .B2(_21643_),
    .ZN(_02615_));
 MUX2_X1 _50209_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2615]),
    .B(_21479_),
    .S(_21639_),
    .Z(_02616_));
 MUX2_X1 _50210_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2616]),
    .B(_21480_),
    .S(_21639_),
    .Z(_02617_));
 MUX2_X1 _50211_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2617]),
    .B(_21481_),
    .S(_21639_),
    .Z(_02618_));
 MUX2_X1 _50212_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2618]),
    .B(_21482_),
    .S(_21639_),
    .Z(_02619_));
 MUX2_X1 _50213_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2619]),
    .B(_21483_),
    .S(_21639_),
    .Z(_02620_));
 MUX2_X1 _50214_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2620]),
    .B(_21588_),
    .S(_21639_),
    .Z(_02622_));
 MUX2_X1 _50215_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2621]),
    .B(_21484_),
    .S(_21639_),
    .Z(_02623_));
 MUX2_X1 _50216_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2622]),
    .B(_21617_),
    .S(_21639_),
    .Z(_02624_));
 MUX2_X1 _50217_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2623]),
    .B(_21485_),
    .S(_21639_),
    .Z(_02625_));
 BUF_X16 _50218_ (.A(_21632_),
    .Z(_21644_));
 MUX2_X1 _50219_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2624]),
    .B(_21554_),
    .S(_21644_),
    .Z(_02626_));
 NAND4_X1 _50220_ (.A1(_21640_),
    .A2(_10585_),
    .A3(_21592_),
    .A4(_21641_),
    .ZN(_21645_));
 INV_X1 _50221_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2625]),
    .ZN(_21646_));
 OAI21_X1 _50222_ (.A(_21645_),
    .B1(_21634_),
    .B2(_21646_),
    .ZN(_02627_));
 MUX2_X1 _50223_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2626]),
    .B(_21590_),
    .S(_21644_),
    .Z(_02628_));
 NAND4_X1 _50224_ (.A1(_21640_),
    .A2(_21558_),
    .A3(_21592_),
    .A4(_21641_),
    .ZN(_21647_));
 INV_X1 _50225_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2627]),
    .ZN(_21648_));
 OAI21_X1 _50226_ (.A(_21647_),
    .B1(_21634_),
    .B2(_21648_),
    .ZN(_02629_));
 MUX2_X1 _50227_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2628]),
    .B(_21561_),
    .S(_21644_),
    .Z(_02630_));
 MUX2_X1 _50228_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2629]),
    .B(_21491_),
    .S(_21644_),
    .Z(_02631_));
 MUX2_X1 _50229_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2630]),
    .B(_21492_),
    .S(_21644_),
    .Z(_02633_));
 MUX2_X1 _50230_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2631]),
    .B(_21621_),
    .S(_21644_),
    .Z(_02634_));
 MUX2_X1 _50231_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2632]),
    .B(_21496_),
    .S(_21644_),
    .Z(_02635_));
 MUX2_X1 _50232_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2633]),
    .B(_21497_),
    .S(_21644_),
    .Z(_02636_));
 MUX2_X1 _50233_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2634]),
    .B(_21566_),
    .S(_21644_),
    .Z(_02637_));
 MUX2_X1 _50234_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2635]),
    .B(_21498_),
    .S(_21644_),
    .Z(_02638_));
 MUX2_X1 _50235_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2636]),
    .B(_21340_),
    .S(_21633_),
    .Z(_02639_));
 BUF_X4 _50236_ (.A(_21343_),
    .Z(_21649_));
 MUX2_X1 _50237_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2637]),
    .B(_21649_),
    .S(_21633_),
    .Z(_02640_));
 MUX2_X1 _50238_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2638]),
    .B(_21348_),
    .S(_21633_),
    .Z(_02641_));
 NAND4_X1 _50239_ (.A1(_21640_),
    .A2(_21499_),
    .A3(_21626_),
    .A4(_21461_),
    .ZN(_21650_));
 INV_X1 _50240_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2639]),
    .ZN(_21651_));
 OAI21_X1 _50241_ (.A(_21650_),
    .B1(_21634_),
    .B2(_21651_),
    .ZN(_02642_));
 MUX2_X1 _50242_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2640]),
    .B(_21356_),
    .S(_21633_),
    .Z(_02644_));
 MUX2_X1 _50243_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2641]),
    .B(_21410_),
    .S(_21633_),
    .Z(_02645_));
 BUF_X4 _50244_ (.A(_21365_),
    .Z(_21652_));
 MUX2_X1 _50245_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2642]),
    .B(_21652_),
    .S(_21633_),
    .Z(_02646_));
 MUX2_X1 _50246_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2643]),
    .B(_21370_),
    .S(_21633_),
    .Z(_02647_));
 BUF_X8 _50247_ (.A(_21373_),
    .Z(_21653_));
 MUX2_X1 _50248_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2644]),
    .B(_21653_),
    .S(_21633_),
    .Z(_02648_));
 MUX2_X1 _50249_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2645]),
    .B(_21411_),
    .S(_21633_),
    .Z(_02649_));
 BUF_X8 _50250_ (.A(_10907_),
    .Z(_21654_));
 AND2_X4 _50251_ (.A1(_21654_),
    .A2(_21441_),
    .ZN(_21655_));
 BUF_X16 _50252_ (.A(_21655_),
    .Z(_21656_));
 BUF_X8 _50253_ (.A(_21656_),
    .Z(_21657_));
 MUX2_X1 _50254_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2548]),
    .B(_21599_),
    .S(_21657_),
    .Z(_02541_));
 MUX2_X1 _50255_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2549]),
    .B(_21606_),
    .S(_21657_),
    .Z(_02542_));
 MUX2_X1 _50256_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2550]),
    .B(_21295_),
    .S(_21657_),
    .Z(_02544_));
 BUF_X16 _50257_ (.A(_21655_),
    .Z(_21658_));
 MUX2_X1 _50258_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2551]),
    .B(_21609_),
    .S(_21658_),
    .Z(_02545_));
 MUX2_X1 _50259_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2552]),
    .B(_21298_),
    .S(_21658_),
    .Z(_02546_));
 MUX2_X1 _50260_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2553]),
    .B(_21635_),
    .S(_21658_),
    .Z(_02547_));
 MUX2_X1 _50261_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2554]),
    .B(_21302_),
    .S(_21658_),
    .Z(_02548_));
 MUX2_X1 _50262_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2555]),
    .B(_21304_),
    .S(_21658_),
    .Z(_02549_));
 MUX2_X1 _50263_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2556]),
    .B(_21306_),
    .S(_21658_),
    .Z(_02550_));
 MUX2_X1 _50264_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2557]),
    .B(_21308_),
    .S(_21658_),
    .Z(_02551_));
 BUF_X4 _50265_ (.A(_21314_),
    .Z(_21659_));
 NAND4_X1 _50266_ (.A1(_21452_),
    .A2(_21446_),
    .A3(_21659_),
    .A4(_21641_),
    .ZN(_21660_));
 INV_X2 _50267_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2558]),
    .ZN(_21661_));
 OAI21_X1 _50268_ (.A(_21660_),
    .B1(_21657_),
    .B2(_21661_),
    .ZN(_02552_));
 MUX2_X1 _50269_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2559]),
    .B(_21312_),
    .S(_21658_),
    .Z(_02553_));
 MUX2_X1 _50270_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2560]),
    .B(_21473_),
    .S(_21658_),
    .Z(_02555_));
 MUX2_X1 _50271_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2561]),
    .B(_21586_),
    .S(_21658_),
    .Z(_02556_));
 BUF_X8 _50272_ (.A(_21655_),
    .Z(_21662_));
 MUX2_X1 _50273_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2562]),
    .B(_21512_),
    .S(_21662_),
    .Z(_02557_));
 MUX2_X1 _50274_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2563]),
    .B(_21476_),
    .S(_21662_),
    .Z(_02558_));
 MUX2_X1 _50275_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2564]),
    .B(_21477_),
    .S(_21662_),
    .Z(_02559_));
 NAND4_X1 _50276_ (.A1(_21452_),
    .A2(_10599_),
    .A3(_21659_),
    .A4(_21641_),
    .ZN(_21663_));
 INV_X1 _50277_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2565]),
    .ZN(_21664_));
 OAI21_X1 _50278_ (.A(_21663_),
    .B1(_21657_),
    .B2(_21664_),
    .ZN(_02560_));
 MUX2_X1 _50279_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2566]),
    .B(_21479_),
    .S(_21662_),
    .Z(_02561_));
 MUX2_X1 _50280_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2567]),
    .B(_21480_),
    .S(_21662_),
    .Z(_02562_));
 MUX2_X1 _50281_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2568]),
    .B(_21481_),
    .S(_21662_),
    .Z(_02563_));
 MUX2_X1 _50282_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2569]),
    .B(_21482_),
    .S(_21662_),
    .Z(_02564_));
 MUX2_X1 _50283_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2570]),
    .B(_21483_),
    .S(_21662_),
    .Z(_02566_));
 MUX2_X1 _50284_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2571]),
    .B(_21588_),
    .S(_21662_),
    .Z(_02567_));
 MUX2_X1 _50285_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2572]),
    .B(_21484_),
    .S(_21662_),
    .Z(_02568_));
 BUF_X16 _50286_ (.A(_21655_),
    .Z(_21665_));
 MUX2_X1 _50287_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2573]),
    .B(_21617_),
    .S(_21665_),
    .Z(_02569_));
 MUX2_X1 _50288_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2574]),
    .B(_21485_),
    .S(_21665_),
    .Z(_02570_));
 MUX2_X1 _50289_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2575]),
    .B(_21554_),
    .S(_21665_),
    .Z(_02571_));
 NAND4_X1 _50290_ (.A1(_21452_),
    .A2(_10585_),
    .A3(_21659_),
    .A4(_21641_),
    .ZN(_21666_));
 INV_X1 _50291_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2576]),
    .ZN(_21667_));
 OAI21_X1 _50292_ (.A(_21666_),
    .B1(_21657_),
    .B2(_21667_),
    .ZN(_02572_));
 MUX2_X1 _50293_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2577]),
    .B(_21590_),
    .S(_21665_),
    .Z(_02573_));
 MUX2_X1 _50294_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2578]),
    .B(_21490_),
    .S(_21665_),
    .Z(_02574_));
 NAND4_X1 _50295_ (.A1(_21452_),
    .A2(_08614_),
    .A3(_21659_),
    .A4(_21641_),
    .ZN(_21668_));
 INV_X4 _50296_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2579]),
    .ZN(_21669_));
 OAI21_X1 _50297_ (.A(_21668_),
    .B1(_21657_),
    .B2(_21669_),
    .ZN(_02575_));
 MUX2_X1 _50298_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2580]),
    .B(_21491_),
    .S(_21665_),
    .Z(_02577_));
 MUX2_X1 _50299_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2581]),
    .B(_21492_),
    .S(_21665_),
    .Z(_02578_));
 MUX2_X1 _50300_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2582]),
    .B(_21621_),
    .S(_21665_),
    .Z(_02579_));
 MUX2_X1 _50301_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2583]),
    .B(_21496_),
    .S(_21665_),
    .Z(_02580_));
 MUX2_X1 _50302_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2584]),
    .B(_21497_),
    .S(_21665_),
    .Z(_02581_));
 MUX2_X1 _50303_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2585]),
    .B(_21566_),
    .S(_21656_),
    .Z(_02582_));
 NAND4_X1 _50304_ (.A1(_21452_),
    .A2(_21591_),
    .A3(_21659_),
    .A4(_21641_),
    .ZN(_21670_));
 INV_X4 _50305_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2586]),
    .ZN(_21671_));
 OAI21_X1 _50306_ (.A(_21670_),
    .B1(_21657_),
    .B2(_21671_),
    .ZN(_02583_));
 MUX2_X1 _50307_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2587]),
    .B(_21340_),
    .S(_21656_),
    .Z(_02584_));
 MUX2_X1 _50308_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2588]),
    .B(_21649_),
    .S(_21656_),
    .Z(_02585_));
 MUX2_X1 _50309_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2589]),
    .B(_21348_),
    .S(_21656_),
    .Z(_02586_));
 BUF_X16 _50310_ (.A(_10845_),
    .Z(_21672_));
 BUF_X8 _50311_ (.A(_11015_),
    .Z(_21673_));
 NAND4_X1 _50312_ (.A1(_21672_),
    .A2(_21673_),
    .A3(_21626_),
    .A4(_21461_),
    .ZN(_21674_));
 INV_X2 _50313_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2590]),
    .ZN(_21675_));
 OAI21_X1 _50314_ (.A(_21674_),
    .B1(_21657_),
    .B2(_21675_),
    .ZN(_02588_));
 NAND4_X2 _50315_ (.A1(_21672_),
    .A2(_21673_),
    .A3(_21626_),
    .A4(_21533_),
    .ZN(_21676_));
 INV_X1 _50316_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2591]),
    .ZN(_21677_));
 OAI21_X1 _50317_ (.A(_21676_),
    .B1(_21657_),
    .B2(_21677_),
    .ZN(_02589_));
 MUX2_X1 _50318_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2592]),
    .B(_21410_),
    .S(_21656_),
    .Z(_02590_));
 MUX2_X1 _50319_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2593]),
    .B(_21652_),
    .S(_21656_),
    .Z(_02591_));
 BUF_X4 _50320_ (.A(_21369_),
    .Z(_21678_));
 MUX2_X1 _50321_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2594]),
    .B(_21678_),
    .S(_21656_),
    .Z(_02592_));
 MUX2_X1 _50322_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2595]),
    .B(_21653_),
    .S(_21656_),
    .Z(_02593_));
 MUX2_X1 _50323_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2596]),
    .B(_21411_),
    .S(_21656_),
    .Z(_02594_));
 BUF_X32 _50324_ (.A(_10762_),
    .Z(_21679_));
 AND2_X4 _50325_ (.A1(_10912_),
    .A2(_21679_),
    .ZN(_21680_));
 BUF_X16 _50326_ (.A(_21680_),
    .Z(_21681_));
 BUF_X8 _50327_ (.A(_21681_),
    .Z(_21682_));
 MUX2_X1 _50328_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2499]),
    .B(_21599_),
    .S(_21682_),
    .Z(_02486_));
 MUX2_X1 _50329_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2500]),
    .B(_21606_),
    .S(_21682_),
    .Z(_02489_));
 BUF_X4 _50330_ (.A(_21294_),
    .Z(_21683_));
 MUX2_X1 _50331_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2501]),
    .B(_21683_),
    .S(_21682_),
    .Z(_02490_));
 MUX2_X1 _50332_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2502]),
    .B(_21609_),
    .S(_21682_),
    .Z(_02491_));
 BUF_X8 _50333_ (.A(_21297_),
    .Z(_21684_));
 BUF_X16 _50334_ (.A(_21680_),
    .Z(_21685_));
 MUX2_X1 _50335_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2503]),
    .B(_21684_),
    .S(_21685_),
    .Z(_02492_));
 MUX2_X1 _50336_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2504]),
    .B(_21635_),
    .S(_21685_),
    .Z(_02493_));
 NAND4_X1 _50337_ (.A1(_21486_),
    .A2(_21578_),
    .A3(_21659_),
    .A4(_21641_),
    .ZN(_21686_));
 INV_X1 _50338_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2505]),
    .ZN(_21687_));
 OAI21_X1 _50339_ (.A(_21686_),
    .B1(_21682_),
    .B2(_21687_),
    .ZN(_02494_));
 BUF_X8 _50340_ (.A(_21303_),
    .Z(_21688_));
 MUX2_X1 _50341_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2506]),
    .B(_21688_),
    .S(_21685_),
    .Z(_02495_));
 BUF_X8 _50342_ (.A(_21305_),
    .Z(_21689_));
 MUX2_X1 _50343_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2507]),
    .B(_21689_),
    .S(_21685_),
    .Z(_02496_));
 MUX2_X1 _50344_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2508]),
    .B(_21308_),
    .S(_21685_),
    .Z(_02497_));
 MUX2_X1 _50345_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2509]),
    .B(_21310_),
    .S(_21685_),
    .Z(_02498_));
 NAND4_X1 _50346_ (.A1(_21486_),
    .A2(_21506_),
    .A3(_21659_),
    .A4(_21641_),
    .ZN(_21690_));
 INV_X1 _50347_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2510]),
    .ZN(_21691_));
 OAI21_X1 _50348_ (.A(_21690_),
    .B1(_21682_),
    .B2(_21691_),
    .ZN(_02500_));
 MUX2_X1 _50349_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2511]),
    .B(_21473_),
    .S(_21685_),
    .Z(_02501_));
 MUX2_X1 _50350_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2512]),
    .B(_21586_),
    .S(_21685_),
    .Z(_02502_));
 MUX2_X1 _50351_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2513]),
    .B(_21512_),
    .S(_21685_),
    .Z(_02503_));
 MUX2_X1 _50352_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2514]),
    .B(_21476_),
    .S(_21685_),
    .Z(_02504_));
 BUF_X16 _50353_ (.A(_21680_),
    .Z(_21692_));
 MUX2_X1 _50354_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2515]),
    .B(_21477_),
    .S(_21692_),
    .Z(_02505_));
 MUX2_X1 _50355_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2516]),
    .B(_21516_),
    .S(_21692_),
    .Z(_02506_));
 MUX2_X1 _50356_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2517]),
    .B(_21479_),
    .S(_21692_),
    .Z(_02507_));
 MUX2_X1 _50357_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2518]),
    .B(_21480_),
    .S(_21692_),
    .Z(_02508_));
 MUX2_X1 _50358_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2519]),
    .B(_21481_),
    .S(_21692_),
    .Z(_02509_));
 MUX2_X1 _50359_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2520]),
    .B(_21482_),
    .S(_21692_),
    .Z(_02511_));
 MUX2_X1 _50360_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2521]),
    .B(_21483_),
    .S(_21692_),
    .Z(_02512_));
 MUX2_X1 _50361_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2522]),
    .B(_21588_),
    .S(_21692_),
    .Z(_02513_));
 BUF_X2 _50362_ (.A(_10893_),
    .Z(_21693_));
 NAND4_X1 _50363_ (.A1(_21486_),
    .A2(_10602_),
    .A3(_21659_),
    .A4(_21693_),
    .ZN(_21694_));
 INV_X1 _50364_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2523]),
    .ZN(_21695_));
 OAI21_X1 _50365_ (.A(_21694_),
    .B1(_21682_),
    .B2(_21695_),
    .ZN(_02514_));
 MUX2_X1 _50366_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2524]),
    .B(_21617_),
    .S(_21692_),
    .Z(_02515_));
 MUX2_X1 _50367_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2525]),
    .B(_21485_),
    .S(_21692_),
    .Z(_02516_));
 BUF_X16 _50368_ (.A(_21680_),
    .Z(_21696_));
 MUX2_X1 _50369_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2526]),
    .B(_21554_),
    .S(_21696_),
    .Z(_02517_));
 NAND4_X1 _50370_ (.A1(_21486_),
    .A2(_10585_),
    .A3(_21659_),
    .A4(_21693_),
    .ZN(_21697_));
 INV_X1 _50371_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2527]),
    .ZN(_21698_));
 OAI21_X1 _50372_ (.A(_21697_),
    .B1(_21682_),
    .B2(_21698_),
    .ZN(_02518_));
 MUX2_X1 _50373_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2528]),
    .B(_21590_),
    .S(_21696_),
    .Z(_02519_));
 MUX2_X1 _50374_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2529]),
    .B(_21490_),
    .S(_21696_),
    .Z(_02520_));
 MUX2_X1 _50375_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2530]),
    .B(_21561_),
    .S(_21696_),
    .Z(_02522_));
 MUX2_X1 _50376_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2531]),
    .B(_21491_),
    .S(_21696_),
    .Z(_02523_));
 MUX2_X1 _50377_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2532]),
    .B(_21492_),
    .S(_21696_),
    .Z(_02524_));
 MUX2_X1 _50378_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2533]),
    .B(_21621_),
    .S(_21696_),
    .Z(_02525_));
 MUX2_X1 _50379_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2534]),
    .B(_21496_),
    .S(_21696_),
    .Z(_02526_));
 MUX2_X1 _50380_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2535]),
    .B(_21497_),
    .S(_21696_),
    .Z(_02527_));
 MUX2_X1 _50381_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2536]),
    .B(_21566_),
    .S(_21696_),
    .Z(_02528_));
 MUX2_X1 _50382_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2537]),
    .B(_21498_),
    .S(_21681_),
    .Z(_02529_));
 NAND4_X1 _50383_ (.A1(_21486_),
    .A2(_21673_),
    .A3(_21626_),
    .A4(_21595_),
    .ZN(_21699_));
 INV_X1 _50384_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2538]),
    .ZN(_21700_));
 OAI21_X1 _50385_ (.A(_21699_),
    .B1(_21682_),
    .B2(_21700_),
    .ZN(_02530_));
 MUX2_X1 _50386_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2539]),
    .B(_21649_),
    .S(_21681_),
    .Z(_02531_));
 MUX2_X1 _50387_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2540]),
    .B(_21348_),
    .S(_21681_),
    .Z(_02533_));
 MUX2_X1 _50388_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2541]),
    .B(_21352_),
    .S(_21681_),
    .Z(_02534_));
 NAND4_X1 _50389_ (.A1(_21486_),
    .A2(_21673_),
    .A3(_21626_),
    .A4(_21533_),
    .ZN(_21701_));
 INV_X1 _50390_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2542]),
    .ZN(_21702_));
 OAI21_X1 _50391_ (.A(_21701_),
    .B1(_21682_),
    .B2(_21702_),
    .ZN(_02535_));
 BUF_X4 _50392_ (.A(_21359_),
    .Z(_21703_));
 MUX2_X1 _50393_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2543]),
    .B(_21703_),
    .S(_21681_),
    .Z(_02536_));
 MUX2_X1 _50394_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2544]),
    .B(_21652_),
    .S(_21681_),
    .Z(_02537_));
 MUX2_X1 _50395_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2545]),
    .B(_21678_),
    .S(_21681_),
    .Z(_02538_));
 MUX2_X1 _50396_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2546]),
    .B(_21653_),
    .S(_21681_),
    .Z(_02539_));
 BUF_X4 _50397_ (.A(_21377_),
    .Z(_21704_));
 MUX2_X1 _50398_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2547]),
    .B(_21704_),
    .S(_21681_),
    .Z(_02540_));
 BUF_X16 _50399_ (.A(_10916_),
    .Z(_21705_));
 AND2_X4 _50400_ (.A1(_21705_),
    .A2(_10784_),
    .ZN(_21706_));
 BUF_X8 _50401_ (.A(_21706_),
    .Z(_21707_));
 MUX2_X1 _50402_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2450]),
    .B(_21599_),
    .S(_21707_),
    .Z(_02433_));
 MUX2_X1 _50403_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2451]),
    .B(_21606_),
    .S(_21707_),
    .Z(_02434_));
 MUX2_X1 _50404_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2452]),
    .B(_21683_),
    .S(_21707_),
    .Z(_02435_));
 MUX2_X1 _50405_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2453]),
    .B(_21609_),
    .S(_21707_),
    .Z(_02436_));
 MUX2_X1 _50406_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2454]),
    .B(_21684_),
    .S(_21707_),
    .Z(_02437_));
 MUX2_X1 _50407_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2455]),
    .B(_21635_),
    .S(_21707_),
    .Z(_02438_));
 NAND4_X1 _50408_ (.A1(_21513_),
    .A2(_21578_),
    .A3(_21659_),
    .A4(_21693_),
    .ZN(_21708_));
 BUF_X4 _50409_ (.A(_21707_),
    .Z(_21709_));
 INV_X1 _50410_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2456]),
    .ZN(_21710_));
 OAI21_X1 _50411_ (.A(_21708_),
    .B1(_21709_),
    .B2(_21710_),
    .ZN(_02439_));
 MUX2_X1 _50412_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2457]),
    .B(_21688_),
    .S(_21707_),
    .Z(_02440_));
 MUX2_X1 _50413_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2458]),
    .B(_21689_),
    .S(_21707_),
    .Z(_02441_));
 BUF_X4 _50414_ (.A(_21314_),
    .Z(_21711_));
 NAND4_X1 _50415_ (.A1(_21513_),
    .A2(_21307_),
    .A3(_21711_),
    .A4(_21693_),
    .ZN(_21712_));
 INV_X2 _50416_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2459]),
    .ZN(_21713_));
 OAI21_X1 _50417_ (.A(_21712_),
    .B1(_21709_),
    .B2(_21713_),
    .ZN(_02442_));
 BUF_X4 _50418_ (.A(_21309_),
    .Z(_21714_));
 BUF_X16 _50419_ (.A(_21706_),
    .Z(_21715_));
 MUX2_X1 _50420_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2460]),
    .B(_21714_),
    .S(_21715_),
    .Z(_02444_));
 BUF_X4 _50421_ (.A(_10859_),
    .Z(_21716_));
 BUF_X16 _50422_ (.A(_21311_),
    .Z(_21717_));
 NAND4_X1 _50423_ (.A1(_21716_),
    .A2(_21717_),
    .A3(_21711_),
    .A4(_21693_),
    .ZN(_21718_));
 INV_X1 _50424_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2461]),
    .ZN(_21719_));
 OAI21_X1 _50425_ (.A(_21718_),
    .B1(_21709_),
    .B2(_21719_),
    .ZN(_02445_));
 MUX2_X1 _50426_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2462]),
    .B(_21473_),
    .S(_21715_),
    .Z(_02446_));
 MUX2_X1 _50427_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2463]),
    .B(_21586_),
    .S(_21715_),
    .Z(_02447_));
 MUX2_X1 _50428_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2464]),
    .B(_21512_),
    .S(_21715_),
    .Z(_02448_));
 MUX2_X1 _50429_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2465]),
    .B(_21476_),
    .S(_21715_),
    .Z(_02449_));
 MUX2_X1 _50430_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2466]),
    .B(_21477_),
    .S(_21715_),
    .Z(_02450_));
 MUX2_X1 _50431_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2467]),
    .B(_21516_),
    .S(_21715_),
    .Z(_02451_));
 MUX2_X1 _50432_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2468]),
    .B(_21479_),
    .S(_21715_),
    .Z(_02452_));
 MUX2_X1 _50433_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2469]),
    .B(_21480_),
    .S(_21715_),
    .Z(_02453_));
 MUX2_X1 _50434_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2470]),
    .B(_21481_),
    .S(_21715_),
    .Z(_02455_));
 BUF_X16 _50435_ (.A(_21706_),
    .Z(_21720_));
 MUX2_X1 _50436_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2471]),
    .B(_21482_),
    .S(_21720_),
    .Z(_02456_));
 MUX2_X1 _50437_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2472]),
    .B(_21483_),
    .S(_21720_),
    .Z(_02457_));
 NAND4_X1 _50438_ (.A1(_21716_),
    .A2(_10580_),
    .A3(_21711_),
    .A4(_21693_),
    .ZN(_21721_));
 INV_X1 _50439_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2473]),
    .ZN(_21722_));
 OAI21_X1 _50440_ (.A(_21721_),
    .B1(_21709_),
    .B2(_21722_),
    .ZN(_02458_));
 NAND4_X1 _50441_ (.A1(_21716_),
    .A2(_10602_),
    .A3(_21711_),
    .A4(_21693_),
    .ZN(_21723_));
 INV_X1 _50442_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2474]),
    .ZN(_21724_));
 OAI21_X1 _50443_ (.A(_21723_),
    .B1(_21709_),
    .B2(_21724_),
    .ZN(_02459_));
 MUX2_X1 _50444_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2475]),
    .B(_21617_),
    .S(_21720_),
    .Z(_02460_));
 MUX2_X1 _50445_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2476]),
    .B(_21485_),
    .S(_21720_),
    .Z(_02461_));
 MUX2_X1 _50446_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2477]),
    .B(_21554_),
    .S(_21720_),
    .Z(_02462_));
 BUF_X16 _50447_ (.A(_08604_),
    .Z(_21725_));
 NAND4_X1 _50448_ (.A1(_21716_),
    .A2(_21725_),
    .A3(_21711_),
    .A4(_21693_),
    .ZN(_21726_));
 INV_X1 _50449_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2478]),
    .ZN(_21727_));
 OAI21_X1 _50450_ (.A(_21726_),
    .B1(_21709_),
    .B2(_21727_),
    .ZN(_02463_));
 MUX2_X1 _50451_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2479]),
    .B(_21590_),
    .S(_21720_),
    .Z(_02464_));
 NAND4_X1 _50452_ (.A1(_21716_),
    .A2(_21558_),
    .A3(_21711_),
    .A4(_21693_),
    .ZN(_21728_));
 INV_X1 _50453_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2480]),
    .ZN(_21729_));
 OAI21_X1 _50454_ (.A(_21728_),
    .B1(_21709_),
    .B2(_21729_),
    .ZN(_02466_));
 MUX2_X1 _50455_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2481]),
    .B(_21561_),
    .S(_21720_),
    .Z(_02467_));
 MUX2_X1 _50456_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2482]),
    .B(_21491_),
    .S(_21720_),
    .Z(_02468_));
 MUX2_X1 _50457_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2483]),
    .B(_21492_),
    .S(_21720_),
    .Z(_02469_));
 MUX2_X1 _50458_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2484]),
    .B(_21621_),
    .S(_21720_),
    .Z(_02470_));
 BUF_X16 _50459_ (.A(_21706_),
    .Z(_21730_));
 MUX2_X1 _50460_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2485]),
    .B(_21496_),
    .S(_21730_),
    .Z(_02471_));
 MUX2_X1 _50461_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2486]),
    .B(_21497_),
    .S(_21730_),
    .Z(_02472_));
 MUX2_X1 _50462_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2487]),
    .B(_21566_),
    .S(_21730_),
    .Z(_02473_));
 NAND4_X1 _50463_ (.A1(_21716_),
    .A2(_21591_),
    .A3(_21711_),
    .A4(_21693_),
    .ZN(_21731_));
 INV_X1 _50464_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2488]),
    .ZN(_21732_));
 OAI21_X1 _50465_ (.A(_21731_),
    .B1(_21709_),
    .B2(_21732_),
    .ZN(_02474_));
 NAND4_X1 _50466_ (.A1(_21716_),
    .A2(_21673_),
    .A3(_21626_),
    .A4(_21595_),
    .ZN(_21733_));
 INV_X1 _50467_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2489]),
    .ZN(_21734_));
 OAI21_X1 _50468_ (.A(_21733_),
    .B1(_21709_),
    .B2(_21734_),
    .ZN(_02475_));
 MUX2_X1 _50469_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2490]),
    .B(_21649_),
    .S(_21730_),
    .Z(_02477_));
 NAND4_X1 _50470_ (.A1(_21716_),
    .A2(_21673_),
    .A3(_21626_),
    .A4(_21347_),
    .ZN(_21735_));
 INV_X2 _50471_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2491]),
    .ZN(_21736_));
 OAI21_X1 _50472_ (.A(_21735_),
    .B1(_21709_),
    .B2(_21736_),
    .ZN(_02478_));
 BUF_X8 _50473_ (.A(_21351_),
    .Z(_21737_));
 MUX2_X1 _50474_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2492]),
    .B(_21737_),
    .S(_21730_),
    .Z(_02479_));
 BUF_X32 _50475_ (.A(_21355_),
    .Z(_21738_));
 NAND4_X1 _50476_ (.A1(_21716_),
    .A2(_21673_),
    .A3(_21626_),
    .A4(_21738_),
    .ZN(_21739_));
 INV_X1 _50477_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2493]),
    .ZN(_21740_));
 OAI21_X1 _50478_ (.A(_21739_),
    .B1(_21707_),
    .B2(_21740_),
    .ZN(_02480_));
 MUX2_X1 _50479_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2494]),
    .B(_21703_),
    .S(_21730_),
    .Z(_02481_));
 MUX2_X1 _50480_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2495]),
    .B(_21652_),
    .S(_21730_),
    .Z(_02482_));
 MUX2_X1 _50481_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2496]),
    .B(_21678_),
    .S(_21730_),
    .Z(_02483_));
 MUX2_X1 _50482_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2497]),
    .B(_21653_),
    .S(_21730_),
    .Z(_02484_));
 MUX2_X1 _50483_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2498]),
    .B(_21704_),
    .S(_21730_),
    .Z(_02485_));
 AND2_X4 _50484_ (.A1(_10921_),
    .A2(_21412_),
    .ZN(_21741_));
 BUF_X16 _50485_ (.A(_21741_),
    .Z(_21742_));
 BUF_X8 _50486_ (.A(_21742_),
    .Z(_21743_));
 MUX2_X1 _50487_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2401]),
    .B(_21599_),
    .S(_21743_),
    .Z(_02379_));
 MUX2_X1 _50488_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2402]),
    .B(_21606_),
    .S(_21743_),
    .Z(_02380_));
 MUX2_X1 _50489_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2403]),
    .B(_21683_),
    .S(_21743_),
    .Z(_02381_));
 MUX2_X1 _50490_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2404]),
    .B(_21609_),
    .S(_21743_),
    .Z(_02382_));
 MUX2_X1 _50491_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2405]),
    .B(_21684_),
    .S(_21743_),
    .Z(_02383_));
 BUF_X16 _50492_ (.A(_21741_),
    .Z(_21744_));
 MUX2_X1 _50493_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2406]),
    .B(_21635_),
    .S(_21744_),
    .Z(_02384_));
 BUF_X8 _50494_ (.A(_21301_),
    .Z(_21745_));
 MUX2_X1 _50495_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2407]),
    .B(_21745_),
    .S(_21744_),
    .Z(_02385_));
 MUX2_X1 _50496_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2408]),
    .B(_21688_),
    .S(_21744_),
    .Z(_02386_));
 BUF_X4 _50497_ (.A(_10893_),
    .Z(_21746_));
 NAND4_X2 _50498_ (.A1(_21546_),
    .A2(_21392_),
    .A3(_21711_),
    .A4(_21746_),
    .ZN(_21747_));
 INV_X1 _50499_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2409]),
    .ZN(_21748_));
 OAI21_X1 _50500_ (.A(_21747_),
    .B1(_21743_),
    .B2(_21748_),
    .ZN(_02387_));
 BUF_X4 _50501_ (.A(_21307_),
    .Z(_21749_));
 MUX2_X1 _50502_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2410]),
    .B(_21749_),
    .S(_21744_),
    .Z(_02389_));
 MUX2_X1 _50503_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2411]),
    .B(_21714_),
    .S(_21744_),
    .Z(_02390_));
 BUF_X8 _50504_ (.A(_21311_),
    .Z(_21750_));
 MUX2_X1 _50505_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2412]),
    .B(_21750_),
    .S(_21744_),
    .Z(_02391_));
 MUX2_X1 _50506_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2413]),
    .B(_21473_),
    .S(_21744_),
    .Z(_02392_));
 MUX2_X1 _50507_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2414]),
    .B(_21586_),
    .S(_21744_),
    .Z(_02393_));
 MUX2_X1 _50508_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2415]),
    .B(_21512_),
    .S(_21744_),
    .Z(_02394_));
 MUX2_X1 _50509_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2416]),
    .B(_21476_),
    .S(_21744_),
    .Z(_02395_));
 BUF_X16 _50510_ (.A(_21741_),
    .Z(_21751_));
 MUX2_X1 _50511_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2417]),
    .B(_21477_),
    .S(_21751_),
    .Z(_02396_));
 BUF_X8 _50512_ (.A(_10869_),
    .Z(_21752_));
 NAND4_X1 _50513_ (.A1(_21752_),
    .A2(_10599_),
    .A3(_21711_),
    .A4(_21746_),
    .ZN(_21753_));
 INV_X1 _50514_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2418]),
    .ZN(_21754_));
 OAI21_X1 _50515_ (.A(_21753_),
    .B1(_21743_),
    .B2(_21754_),
    .ZN(_02397_));
 MUX2_X1 _50516_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2419]),
    .B(_21479_),
    .S(_21751_),
    .Z(_02398_));
 MUX2_X1 _50517_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2420]),
    .B(_21480_),
    .S(_21751_),
    .Z(_02400_));
 MUX2_X1 _50518_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2421]),
    .B(_21481_),
    .S(_21751_),
    .Z(_02401_));
 MUX2_X1 _50519_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2422]),
    .B(_21482_),
    .S(_21751_),
    .Z(_02402_));
 MUX2_X1 _50520_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2423]),
    .B(_21483_),
    .S(_21751_),
    .Z(_02403_));
 NAND4_X1 _50521_ (.A1(_21752_),
    .A2(_10580_),
    .A3(_21711_),
    .A4(_21746_),
    .ZN(_21755_));
 INV_X1 _50522_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2424]),
    .ZN(_21756_));
 OAI21_X1 _50523_ (.A(_21755_),
    .B1(_21743_),
    .B2(_21756_),
    .ZN(_02404_));
 MUX2_X1 _50524_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2425]),
    .B(_21484_),
    .S(_21751_),
    .Z(_02405_));
 BUF_X32 _50525_ (.A(_08594_),
    .Z(_21757_));
 BUF_X8 _50526_ (.A(_21314_),
    .Z(_21758_));
 NAND4_X1 _50527_ (.A1(_21752_),
    .A2(_21757_),
    .A3(_21758_),
    .A4(_21746_),
    .ZN(_21759_));
 INV_X1 _50528_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2426]),
    .ZN(_21760_));
 OAI21_X1 _50529_ (.A(_21759_),
    .B1(_21743_),
    .B2(_21760_),
    .ZN(_02406_));
 MUX2_X1 _50530_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2427]),
    .B(_21485_),
    .S(_21751_),
    .Z(_02407_));
 MUX2_X1 _50531_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2428]),
    .B(_21554_),
    .S(_21751_),
    .Z(_02408_));
 MUX2_X1 _50532_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2429]),
    .B(_21555_),
    .S(_21751_),
    .Z(_02409_));
 BUF_X16 _50533_ (.A(_21741_),
    .Z(_21761_));
 MUX2_X1 _50534_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2430]),
    .B(_21590_),
    .S(_21761_),
    .Z(_02411_));
 MUX2_X1 _50535_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2431]),
    .B(_21490_),
    .S(_21761_),
    .Z(_02412_));
 MUX2_X1 _50536_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2432]),
    .B(_21561_),
    .S(_21761_),
    .Z(_02413_));
 MUX2_X1 _50537_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2433]),
    .B(_21491_),
    .S(_21761_),
    .Z(_02414_));
 MUX2_X1 _50538_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2434]),
    .B(_21492_),
    .S(_21761_),
    .Z(_02415_));
 MUX2_X1 _50539_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2435]),
    .B(_21621_),
    .S(_21761_),
    .Z(_02416_));
 MUX2_X1 _50540_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2436]),
    .B(_21496_),
    .S(_21761_),
    .Z(_02417_));
 MUX2_X1 _50541_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2437]),
    .B(_21497_),
    .S(_21761_),
    .Z(_02418_));
 MUX2_X1 _50542_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2438]),
    .B(_21566_),
    .S(_21761_),
    .Z(_02419_));
 MUX2_X1 _50543_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2439]),
    .B(_21498_),
    .S(_21761_),
    .Z(_02420_));
 BUF_X8 _50544_ (.A(_21339_),
    .Z(_21762_));
 MUX2_X1 _50545_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2440]),
    .B(_21762_),
    .S(_21742_),
    .Z(_02422_));
 BUF_X16 _50546_ (.A(_21343_),
    .Z(_21763_));
 NAND4_X4 _50547_ (.A1(_21752_),
    .A2(_21673_),
    .A3(_21579_),
    .A4(_21763_),
    .ZN(_21764_));
 INV_X1 _50548_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2441]),
    .ZN(_21765_));
 OAI21_X1 _50549_ (.A(_21764_),
    .B1(_21743_),
    .B2(_21765_),
    .ZN(_02423_));
 BUF_X8 _50550_ (.A(_21347_),
    .Z(_21766_));
 MUX2_X1 _50551_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2442]),
    .B(_21766_),
    .S(_21742_),
    .Z(_02424_));
 MUX2_X1 _50552_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2443]),
    .B(_21737_),
    .S(_21742_),
    .Z(_02425_));
 MUX2_X1 _50553_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2444]),
    .B(_21356_),
    .S(_21742_),
    .Z(_02426_));
 MUX2_X1 _50554_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2445]),
    .B(_21703_),
    .S(_21742_),
    .Z(_02427_));
 MUX2_X1 _50555_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2446]),
    .B(_21652_),
    .S(_21742_),
    .Z(_02428_));
 MUX2_X1 _50556_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2447]),
    .B(_21678_),
    .S(_21742_),
    .Z(_02429_));
 MUX2_X1 _50557_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2448]),
    .B(_21653_),
    .S(_21742_),
    .Z(_02430_));
 MUX2_X1 _50558_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2449]),
    .B(_21704_),
    .S(_21742_),
    .Z(_02431_));
 AND2_X4 _50559_ (.A1(_10928_),
    .A2(_21679_),
    .ZN(_21767_));
 BUF_X16 _50560_ (.A(_21767_),
    .Z(_21768_));
 BUF_X8 _50561_ (.A(_21768_),
    .Z(_21769_));
 MUX2_X1 _50562_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2352]),
    .B(_21599_),
    .S(_21769_),
    .Z(_02324_));
 MUX2_X1 _50563_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2353]),
    .B(_21606_),
    .S(_21769_),
    .Z(_02325_));
 MUX2_X1 _50564_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2354]),
    .B(_21683_),
    .S(_21769_),
    .Z(_02326_));
 MUX2_X1 _50565_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2355]),
    .B(_21609_),
    .S(_21769_),
    .Z(_02327_));
 BUF_X16 _50566_ (.A(_21767_),
    .Z(_21770_));
 MUX2_X1 _50567_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2356]),
    .B(_21684_),
    .S(_21770_),
    .Z(_02328_));
 MUX2_X1 _50568_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2357]),
    .B(_21635_),
    .S(_21770_),
    .Z(_02329_));
 MUX2_X1 _50569_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2358]),
    .B(_21745_),
    .S(_21770_),
    .Z(_02330_));
 MUX2_X1 _50570_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2359]),
    .B(_21688_),
    .S(_21770_),
    .Z(_02331_));
 NAND4_X1 _50571_ (.A1(_21322_),
    .A2(_21392_),
    .A3(_21758_),
    .A4(_21746_),
    .ZN(_21771_));
 INV_X1 _50572_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2360]),
    .ZN(_21772_));
 OAI21_X1 _50573_ (.A(_21771_),
    .B1(_21769_),
    .B2(_21772_),
    .ZN(_02333_));
 MUX2_X1 _50574_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2361]),
    .B(_21749_),
    .S(_21770_),
    .Z(_02334_));
 MUX2_X1 _50575_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2362]),
    .B(_21714_),
    .S(_21770_),
    .Z(_02335_));
 MUX2_X1 _50576_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2363]),
    .B(_21750_),
    .S(_21770_),
    .Z(_02336_));
 MUX2_X1 _50577_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2364]),
    .B(_21473_),
    .S(_21770_),
    .Z(_02337_));
 MUX2_X1 _50578_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2365]),
    .B(_21586_),
    .S(_21770_),
    .Z(_02338_));
 MUX2_X1 _50579_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2366]),
    .B(_21512_),
    .S(_21770_),
    .Z(_02339_));
 BUF_X8 _50580_ (.A(_08561_),
    .Z(_21773_));
 BUF_X16 _50581_ (.A(_21767_),
    .Z(_21774_));
 MUX2_X1 _50582_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2367]),
    .B(_21773_),
    .S(_21774_),
    .Z(_02340_));
 MUX2_X1 _50583_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2368]),
    .B(_21477_),
    .S(_21774_),
    .Z(_02341_));
 NAND4_X1 _50584_ (.A1(_21322_),
    .A2(_10599_),
    .A3(_21758_),
    .A4(_21746_),
    .ZN(_21775_));
 INV_X1 _50585_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2369]),
    .ZN(_21776_));
 OAI21_X1 _50586_ (.A(_21775_),
    .B1(_21769_),
    .B2(_21776_),
    .ZN(_02342_));
 MUX2_X1 _50587_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2370]),
    .B(_21479_),
    .S(_21774_),
    .Z(_02344_));
 BUF_X4 _50588_ (.A(_08575_),
    .Z(_21777_));
 MUX2_X1 _50589_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2371]),
    .B(_21777_),
    .S(_21774_),
    .Z(_02345_));
 BUF_X8 _50590_ (.A(_08578_),
    .Z(_21778_));
 MUX2_X1 _50591_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2372]),
    .B(_21778_),
    .S(_21774_),
    .Z(_02346_));
 BUF_X8 _50592_ (.A(_08581_),
    .Z(_21779_));
 MUX2_X1 _50593_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2373]),
    .B(_21779_),
    .S(_21774_),
    .Z(_02347_));
 BUF_X8 _50594_ (.A(_08584_),
    .Z(_21780_));
 MUX2_X1 _50595_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2374]),
    .B(_21780_),
    .S(_21774_),
    .Z(_02348_));
 MUX2_X1 _50596_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2375]),
    .B(_21588_),
    .S(_21774_),
    .Z(_02349_));
 MUX2_X1 _50597_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2376]),
    .B(_21484_),
    .S(_21774_),
    .Z(_02350_));
 NAND4_X1 _50598_ (.A1(_21322_),
    .A2(_21757_),
    .A3(_21758_),
    .A4(_21746_),
    .ZN(_21781_));
 INV_X1 _50599_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2377]),
    .ZN(_21782_));
 OAI21_X1 _50600_ (.A(_21781_),
    .B1(_21769_),
    .B2(_21782_),
    .ZN(_02351_));
 BUF_X8 _50601_ (.A(_08597_),
    .Z(_21783_));
 MUX2_X1 _50602_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2378]),
    .B(_21783_),
    .S(_21774_),
    .Z(_02352_));
 NAND4_X1 _50603_ (.A1(_21322_),
    .A2(_21520_),
    .A3(_21758_),
    .A4(_21746_),
    .ZN(_21784_));
 INV_X1 _50604_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2379]),
    .ZN(_21785_));
 OAI21_X1 _50605_ (.A(_21784_),
    .B1(_21769_),
    .B2(_21785_),
    .ZN(_02353_));
 BUF_X8 _50606_ (.A(_10880_),
    .Z(_21786_));
 NAND4_X1 _50607_ (.A1(_21786_),
    .A2(_21725_),
    .A3(_21758_),
    .A4(_21746_),
    .ZN(_21787_));
 INV_X1 _50608_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2380]),
    .ZN(_21788_));
 OAI21_X1 _50609_ (.A(_21787_),
    .B1(_21769_),
    .B2(_21788_),
    .ZN(_02355_));
 BUF_X8 _50610_ (.A(_21767_),
    .Z(_21789_));
 MUX2_X1 _50611_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2381]),
    .B(_21590_),
    .S(_21789_),
    .Z(_02356_));
 NAND4_X2 _50612_ (.A1(_21786_),
    .A2(_21558_),
    .A3(_21758_),
    .A4(_21746_),
    .ZN(_21790_));
 INV_X1 _50613_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2382]),
    .ZN(_21791_));
 OAI21_X1 _50614_ (.A(_21790_),
    .B1(_21769_),
    .B2(_21791_),
    .ZN(_02357_));
 MUX2_X1 _50615_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2383]),
    .B(_21561_),
    .S(_21789_),
    .Z(_02358_));
 BUF_X8 _50616_ (.A(_08617_),
    .Z(_21792_));
 MUX2_X1 _50617_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2384]),
    .B(_21792_),
    .S(_21789_),
    .Z(_02359_));
 BUF_X8 _50618_ (.A(_08620_),
    .Z(_21793_));
 MUX2_X1 _50619_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2385]),
    .B(_21793_),
    .S(_21789_),
    .Z(_02360_));
 MUX2_X1 _50620_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2386]),
    .B(_21621_),
    .S(_21789_),
    .Z(_02361_));
 BUF_X8 _50621_ (.A(_08626_),
    .Z(_21794_));
 MUX2_X1 _50622_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2387]),
    .B(_21794_),
    .S(_21789_),
    .Z(_02362_));
 BUF_X8 _50623_ (.A(_08629_),
    .Z(_21795_));
 MUX2_X1 _50624_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2388]),
    .B(_21795_),
    .S(_21789_),
    .Z(_02363_));
 MUX2_X1 _50625_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2389]),
    .B(_21566_),
    .S(_21789_),
    .Z(_02364_));
 MUX2_X1 _50626_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2390]),
    .B(_21498_),
    .S(_21789_),
    .Z(_02366_));
 MUX2_X1 _50627_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2391]),
    .B(_21762_),
    .S(_21789_),
    .Z(_02367_));
 MUX2_X1 _50628_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2392]),
    .B(_21649_),
    .S(_21768_),
    .Z(_02368_));
 MUX2_X1 _50629_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2393]),
    .B(_21766_),
    .S(_21768_),
    .Z(_02369_));
 MUX2_X1 _50630_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2394]),
    .B(_21737_),
    .S(_21768_),
    .Z(_02370_));
 MUX2_X1 _50631_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2395]),
    .B(_21356_),
    .S(_21768_),
    .Z(_02371_));
 MUX2_X1 _50632_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2396]),
    .B(_21703_),
    .S(_21768_),
    .Z(_02372_));
 MUX2_X1 _50633_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2397]),
    .B(_21652_),
    .S(_21768_),
    .Z(_02373_));
 MUX2_X1 _50634_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2398]),
    .B(_21678_),
    .S(_21768_),
    .Z(_02374_));
 MUX2_X1 _50635_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2399]),
    .B(_21653_),
    .S(_21768_),
    .Z(_02375_));
 MUX2_X1 _50636_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2400]),
    .B(_21704_),
    .S(_21768_),
    .Z(_02378_));
 AND2_X4 _50637_ (.A1(_10936_),
    .A2(_21574_),
    .ZN(_21796_));
 BUF_X16 _50638_ (.A(_21796_),
    .Z(_21797_));
 BUF_X16 _50639_ (.A(_21797_),
    .Z(_21798_));
 MUX2_X1 _50640_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2303]),
    .B(_21599_),
    .S(_21798_),
    .Z(_02270_));
 MUX2_X1 _50641_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2304]),
    .B(_21606_),
    .S(_21798_),
    .Z(_02271_));
 MUX2_X1 _50642_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2305]),
    .B(_21683_),
    .S(_21798_),
    .Z(_02272_));
 MUX2_X1 _50643_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2306]),
    .B(_21609_),
    .S(_21798_),
    .Z(_02273_));
 MUX2_X1 _50644_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2307]),
    .B(_21684_),
    .S(_21798_),
    .Z(_02274_));
 MUX2_X1 _50645_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2308]),
    .B(_21635_),
    .S(_21798_),
    .Z(_02275_));
 BUF_X8 _50646_ (.A(_10805_),
    .Z(_21799_));
 BUF_X8 _50647_ (.A(_10942_),
    .Z(_21800_));
 NAND4_X2 _50648_ (.A1(_21799_),
    .A2(_21301_),
    .A3(_21758_),
    .A4(_21800_),
    .ZN(_21801_));
 INV_X1 _50649_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2309]),
    .ZN(_21802_));
 OAI21_X1 _50650_ (.A(_21801_),
    .B1(_21798_),
    .B2(_21802_),
    .ZN(_02276_));
 BUF_X8 _50651_ (.A(_21796_),
    .Z(_21803_));
 MUX2_X1 _50652_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2310]),
    .B(_21688_),
    .S(_21803_),
    .Z(_02278_));
 MUX2_X1 _50653_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2311]),
    .B(_21689_),
    .S(_21803_),
    .Z(_02279_));
 MUX2_X1 _50654_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2312]),
    .B(_21749_),
    .S(_21803_),
    .Z(_02280_));
 MUX2_X1 _50655_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2313]),
    .B(_21714_),
    .S(_21803_),
    .Z(_02281_));
 MUX2_X1 _50656_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2314]),
    .B(_21750_),
    .S(_21803_),
    .Z(_02282_));
 MUX2_X1 _50657_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2315]),
    .B(_21473_),
    .S(_21803_),
    .Z(_02283_));
 MUX2_X1 _50658_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2316]),
    .B(_21586_),
    .S(_21803_),
    .Z(_02284_));
 BUF_X8 _50659_ (.A(_08558_),
    .Z(_21804_));
 MUX2_X1 _50660_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2317]),
    .B(_21804_),
    .S(_21803_),
    .Z(_02285_));
 MUX2_X1 _50661_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2318]),
    .B(_21773_),
    .S(_21803_),
    .Z(_02286_));
 BUF_X2 _50662_ (.A(_08564_),
    .Z(_21805_));
 MUX2_X1 _50663_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2319]),
    .B(_21805_),
    .S(_21803_),
    .Z(_02287_));
 BUF_X16 _50664_ (.A(_21796_),
    .Z(_21806_));
 MUX2_X1 _50665_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2320]),
    .B(_21516_),
    .S(_21806_),
    .Z(_02289_));
 BUF_X8 _50666_ (.A(_08571_),
    .Z(_21807_));
 MUX2_X1 _50667_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2321]),
    .B(_21807_),
    .S(_21806_),
    .Z(_02290_));
 MUX2_X1 _50668_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2322]),
    .B(_21777_),
    .S(_21806_),
    .Z(_02291_));
 MUX2_X1 _50669_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2323]),
    .B(_21778_),
    .S(_21806_),
    .Z(_02292_));
 MUX2_X1 _50670_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2324]),
    .B(_21779_),
    .S(_21806_),
    .Z(_02293_));
 MUX2_X1 _50671_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2325]),
    .B(_21780_),
    .S(_21806_),
    .Z(_02294_));
 NAND4_X1 _50672_ (.A1(_21799_),
    .A2(_10580_),
    .A3(_21758_),
    .A4(_21800_),
    .ZN(_21808_));
 INV_X1 _50673_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2326]),
    .ZN(_21809_));
 OAI21_X1 _50674_ (.A(_21808_),
    .B1(_21798_),
    .B2(_21809_),
    .ZN(_02295_));
 MUX2_X1 _50675_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2327]),
    .B(_21484_),
    .S(_21806_),
    .Z(_02296_));
 MUX2_X1 _50676_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2328]),
    .B(_21617_),
    .S(_21806_),
    .Z(_02297_));
 MUX2_X1 _50677_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2329]),
    .B(_21783_),
    .S(_21806_),
    .Z(_02298_));
 MUX2_X1 _50678_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2330]),
    .B(_21554_),
    .S(_21806_),
    .Z(_02300_));
 BUF_X16 _50679_ (.A(_21796_),
    .Z(_21810_));
 MUX2_X1 _50680_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2331]),
    .B(_21555_),
    .S(_21810_),
    .Z(_02301_));
 MUX2_X1 _50681_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2332]),
    .B(_21590_),
    .S(_21810_),
    .Z(_02302_));
 MUX2_X1 _50682_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2333]),
    .B(_21490_),
    .S(_21810_),
    .Z(_02303_));
 MUX2_X1 _50683_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2334]),
    .B(_21561_),
    .S(_21810_),
    .Z(_02304_));
 MUX2_X1 _50684_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2335]),
    .B(_21792_),
    .S(_21810_),
    .Z(_02305_));
 MUX2_X1 _50685_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2336]),
    .B(_21793_),
    .S(_21810_),
    .Z(_02306_));
 MUX2_X1 _50686_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2337]),
    .B(_21621_),
    .S(_21810_),
    .Z(_02307_));
 MUX2_X1 _50687_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2338]),
    .B(_21794_),
    .S(_21810_),
    .Z(_02308_));
 MUX2_X1 _50688_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2339]),
    .B(_21795_),
    .S(_21810_),
    .Z(_02309_));
 MUX2_X1 _50689_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2340]),
    .B(_21566_),
    .S(_21810_),
    .Z(_02311_));
 NAND4_X1 _50690_ (.A1(_21799_),
    .A2(_21591_),
    .A3(_21758_),
    .A4(_21800_),
    .ZN(_21811_));
 INV_X1 _50691_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2341]),
    .ZN(_21812_));
 OAI21_X1 _50692_ (.A(_21811_),
    .B1(_21798_),
    .B2(_21812_),
    .ZN(_02312_));
 MUX2_X1 _50693_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2342]),
    .B(_21762_),
    .S(_21797_),
    .Z(_02313_));
 MUX2_X1 _50694_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2343]),
    .B(_21649_),
    .S(_21797_),
    .Z(_02314_));
 MUX2_X1 _50695_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2344]),
    .B(_21766_),
    .S(_21797_),
    .Z(_02315_));
 NAND4_X1 _50696_ (.A1(_21799_),
    .A2(_21673_),
    .A3(_10943_),
    .A4(_21351_),
    .ZN(_21813_));
 INV_X4 _50697_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2345]),
    .ZN(_21814_));
 OAI21_X1 _50698_ (.A(_21813_),
    .B1(_21798_),
    .B2(_21814_),
    .ZN(_02316_));
 BUF_X4 _50699_ (.A(_21355_),
    .Z(_21815_));
 MUX2_X1 _50700_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2346]),
    .B(_21815_),
    .S(_21797_),
    .Z(_02317_));
 MUX2_X1 _50701_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2347]),
    .B(_21703_),
    .S(_21797_),
    .Z(_02318_));
 MUX2_X1 _50702_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2348]),
    .B(_21652_),
    .S(_21797_),
    .Z(_02319_));
 MUX2_X1 _50703_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2349]),
    .B(_21678_),
    .S(_21797_),
    .Z(_02320_));
 MUX2_X1 _50704_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2350]),
    .B(_21653_),
    .S(_21797_),
    .Z(_02322_));
 MUX2_X1 _50705_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2351]),
    .B(_21704_),
    .S(_21797_),
    .Z(_02323_));
 BUF_X16 _50706_ (.A(_10945_),
    .Z(_21816_));
 AND2_X4 _50707_ (.A1(_21816_),
    .A2(_21290_),
    .ZN(_21817_));
 BUF_X16 _50708_ (.A(_21817_),
    .Z(_21818_));
 BUF_X8 _50709_ (.A(_21818_),
    .Z(_21819_));
 MUX2_X1 _50710_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2254]),
    .B(_21599_),
    .S(_21819_),
    .Z(_02215_));
 BUF_X8 _50711_ (.A(_21817_),
    .Z(_21820_));
 MUX2_X1 _50712_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2255]),
    .B(_21606_),
    .S(_21820_),
    .Z(_02216_));
 BUF_X4 _50713_ (.A(_21314_),
    .Z(_21821_));
 NAND4_X1 _50714_ (.A1(_21629_),
    .A2(_21383_),
    .A3(_21821_),
    .A4(_21800_),
    .ZN(_21822_));
 INV_X1 _50715_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2256]),
    .ZN(_21823_));
 OAI21_X1 _50716_ (.A(_21822_),
    .B1(_21819_),
    .B2(_21823_),
    .ZN(_02217_));
 MUX2_X1 _50717_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2257]),
    .B(_21609_),
    .S(_21820_),
    .Z(_02218_));
 NAND4_X1 _50718_ (.A1(_21629_),
    .A2(_21418_),
    .A3(_21821_),
    .A4(_21800_),
    .ZN(_21824_));
 INV_X1 _50719_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2258]),
    .ZN(_21825_));
 OAI21_X1 _50720_ (.A(_21824_),
    .B1(_21819_),
    .B2(_21825_),
    .ZN(_02219_));
 MUX2_X1 _50721_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2259]),
    .B(_21635_),
    .S(_21820_),
    .Z(_02220_));
 NAND4_X1 _50722_ (.A1(_21629_),
    .A2(_21301_),
    .A3(_21821_),
    .A4(_21800_),
    .ZN(_21826_));
 INV_X1 _50723_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2260]),
    .ZN(_21827_));
 OAI21_X1 _50724_ (.A(_21826_),
    .B1(_21819_),
    .B2(_21827_),
    .ZN(_02222_));
 MUX2_X1 _50725_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2261]),
    .B(_21688_),
    .S(_21820_),
    .Z(_02223_));
 BUF_X8 _50726_ (.A(_10942_),
    .Z(_21828_));
 NAND4_X2 _50727_ (.A1(_21629_),
    .A2(_21392_),
    .A3(_21821_),
    .A4(_21828_),
    .ZN(_21829_));
 INV_X1 _50728_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2262]),
    .ZN(_21830_));
 OAI21_X1 _50729_ (.A(_21829_),
    .B1(_21819_),
    .B2(_21830_),
    .ZN(_02224_));
 MUX2_X1 _50730_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2263]),
    .B(_21749_),
    .S(_21820_),
    .Z(_02225_));
 MUX2_X1 _50731_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2264]),
    .B(_21714_),
    .S(_21820_),
    .Z(_02226_));
 NAND4_X2 _50732_ (.A1(_21629_),
    .A2(_21717_),
    .A3(_21821_),
    .A4(_21828_),
    .ZN(_21831_));
 INV_X1 _50733_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2265]),
    .ZN(_21832_));
 OAI21_X1 _50734_ (.A(_21831_),
    .B1(_21819_),
    .B2(_21832_),
    .ZN(_02227_));
 BUF_X8 _50735_ (.A(_08551_),
    .Z(_21833_));
 MUX2_X1 _50736_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2266]),
    .B(_21833_),
    .S(_21820_),
    .Z(_02228_));
 MUX2_X1 _50737_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2267]),
    .B(_21586_),
    .S(_21820_),
    .Z(_02229_));
 MUX2_X1 _50738_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2268]),
    .B(_21804_),
    .S(_21820_),
    .Z(_02230_));
 MUX2_X1 _50739_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2269]),
    .B(_21773_),
    .S(_21820_),
    .Z(_02231_));
 BUF_X16 _50740_ (.A(_21817_),
    .Z(_21834_));
 MUX2_X1 _50741_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2270]),
    .B(_21805_),
    .S(_21834_),
    .Z(_02233_));
 MUX2_X1 _50742_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2271]),
    .B(_21516_),
    .S(_21834_),
    .Z(_02234_));
 MUX2_X1 _50743_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2272]),
    .B(_21807_),
    .S(_21834_),
    .Z(_02235_));
 MUX2_X1 _50744_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2273]),
    .B(_21777_),
    .S(_21834_),
    .Z(_02236_));
 MUX2_X1 _50745_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2274]),
    .B(_21778_),
    .S(_21834_),
    .Z(_02237_));
 MUX2_X1 _50746_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2275]),
    .B(_21779_),
    .S(_21834_),
    .Z(_02238_));
 MUX2_X1 _50747_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2276]),
    .B(_21780_),
    .S(_21834_),
    .Z(_02239_));
 NAND4_X1 _50748_ (.A1(_21629_),
    .A2(_10580_),
    .A3(_21821_),
    .A4(_21828_),
    .ZN(_21835_));
 INV_X1 _50749_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2277]),
    .ZN(_21836_));
 OAI21_X1 _50750_ (.A(_21835_),
    .B1(_21819_),
    .B2(_21836_),
    .ZN(_02240_));
 BUF_X8 _50751_ (.A(_08591_),
    .Z(_21837_));
 MUX2_X1 _50752_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2278]),
    .B(_21837_),
    .S(_21834_),
    .Z(_02241_));
 MUX2_X1 _50753_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2279]),
    .B(_21617_),
    .S(_21834_),
    .Z(_02242_));
 MUX2_X1 _50754_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2280]),
    .B(_21783_),
    .S(_21834_),
    .Z(_02244_));
 BUF_X16 _50755_ (.A(_21817_),
    .Z(_21838_));
 MUX2_X1 _50756_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2281]),
    .B(_21554_),
    .S(_21838_),
    .Z(_02245_));
 MUX2_X1 _50757_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2282]),
    .B(_21555_),
    .S(_21838_),
    .Z(_02246_));
 MUX2_X1 _50758_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2283]),
    .B(_21590_),
    .S(_21838_),
    .Z(_02247_));
 NAND4_X1 _50759_ (.A1(_21629_),
    .A2(_21558_),
    .A3(_21821_),
    .A4(_21828_),
    .ZN(_21839_));
 INV_X1 _50760_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2284]),
    .ZN(_21840_));
 OAI21_X1 _50761_ (.A(_21839_),
    .B1(_21819_),
    .B2(_21840_),
    .ZN(_02248_));
 MUX2_X1 _50762_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2285]),
    .B(_21561_),
    .S(_21838_),
    .Z(_02249_));
 MUX2_X1 _50763_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2286]),
    .B(_21792_),
    .S(_21838_),
    .Z(_02250_));
 MUX2_X1 _50764_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2287]),
    .B(_21793_),
    .S(_21838_),
    .Z(_02251_));
 MUX2_X1 _50765_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2288]),
    .B(_21621_),
    .S(_21838_),
    .Z(_02252_));
 MUX2_X1 _50766_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2289]),
    .B(_21794_),
    .S(_21838_),
    .Z(_02253_));
 NAND4_X2 _50767_ (.A1(_21629_),
    .A2(_10593_),
    .A3(_21821_),
    .A4(_21828_),
    .ZN(_21841_));
 INV_X1 _50768_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2290]),
    .ZN(_21842_));
 OAI21_X1 _50769_ (.A(_21841_),
    .B1(_21819_),
    .B2(_21842_),
    .ZN(_02255_));
 BUF_X8 _50770_ (.A(_08632_),
    .Z(_21843_));
 MUX2_X1 _50771_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2291]),
    .B(_21843_),
    .S(_21838_),
    .Z(_02256_));
 MUX2_X1 _50772_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2292]),
    .B(_21498_),
    .S(_21838_),
    .Z(_02257_));
 MUX2_X1 _50773_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2293]),
    .B(_21762_),
    .S(_21818_),
    .Z(_02258_));
 MUX2_X1 _50774_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2294]),
    .B(_21649_),
    .S(_21818_),
    .Z(_02259_));
 MUX2_X1 _50775_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2295]),
    .B(_21766_),
    .S(_21818_),
    .Z(_02260_));
 MUX2_X1 _50776_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2296]),
    .B(_21737_),
    .S(_21818_),
    .Z(_02261_));
 MUX2_X1 _50777_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2297]),
    .B(_21815_),
    .S(_21818_),
    .Z(_02262_));
 MUX2_X1 _50778_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2298]),
    .B(_21703_),
    .S(_21818_),
    .Z(_02263_));
 MUX2_X1 _50779_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2299]),
    .B(_21652_),
    .S(_21818_),
    .Z(_02264_));
 MUX2_X1 _50780_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2300]),
    .B(_21678_),
    .S(_21818_),
    .Z(_02267_));
 MUX2_X1 _50781_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2301]),
    .B(_21653_),
    .S(_21818_),
    .Z(_02268_));
 NAND4_X4 _50782_ (.A1(_21629_),
    .A2(_21673_),
    .A3(_10943_),
    .A4(_21377_),
    .ZN(_21844_));
 INV_X1 _50783_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2302]),
    .ZN(_21845_));
 OAI21_X1 _50784_ (.A(_21844_),
    .B1(_21819_),
    .B2(_21845_),
    .ZN(_02269_));
 AND2_X4 _50785_ (.A1(_10950_),
    .A2(_21574_),
    .ZN(_21846_));
 BUF_X16 _50786_ (.A(_21846_),
    .Z(_21847_));
 BUF_X16 _50787_ (.A(_21847_),
    .Z(_21848_));
 MUX2_X1 _50788_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2205]),
    .B(_21599_),
    .S(_21848_),
    .Z(_02161_));
 MUX2_X1 _50789_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2206]),
    .B(_21606_),
    .S(_21848_),
    .Z(_02162_));
 MUX2_X1 _50790_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2207]),
    .B(_21683_),
    .S(_21848_),
    .Z(_02163_));
 MUX2_X1 _50791_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2208]),
    .B(_21609_),
    .S(_21848_),
    .Z(_02164_));
 MUX2_X1 _50792_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2209]),
    .B(_21684_),
    .S(_21848_),
    .Z(_02165_));
 MUX2_X1 _50793_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2210]),
    .B(_21635_),
    .S(_21848_),
    .Z(_02167_));
 MUX2_X1 _50794_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2211]),
    .B(_21745_),
    .S(_21848_),
    .Z(_02168_));
 BUF_X8 _50795_ (.A(_21846_),
    .Z(_21849_));
 MUX2_X1 _50796_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2212]),
    .B(_21688_),
    .S(_21849_),
    .Z(_02169_));
 MUX2_X1 _50797_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2213]),
    .B(_21689_),
    .S(_21849_),
    .Z(_02170_));
 MUX2_X1 _50798_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2214]),
    .B(_21749_),
    .S(_21849_),
    .Z(_02171_));
 MUX2_X1 _50799_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2215]),
    .B(_21714_),
    .S(_21849_),
    .Z(_02172_));
 NAND4_X1 _50800_ (.A1(_21640_),
    .A2(_21717_),
    .A3(_21821_),
    .A4(_21828_),
    .ZN(_21850_));
 INV_X1 _50801_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2216]),
    .ZN(_21851_));
 OAI21_X1 _50802_ (.A(_21850_),
    .B1(_21848_),
    .B2(_21851_),
    .ZN(_02173_));
 MUX2_X1 _50803_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2217]),
    .B(_21833_),
    .S(_21849_),
    .Z(_02174_));
 BUF_X8 _50804_ (.A(_08555_),
    .Z(_21852_));
 MUX2_X1 _50805_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2218]),
    .B(_21852_),
    .S(_21849_),
    .Z(_02175_));
 MUX2_X1 _50806_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2219]),
    .B(_21804_),
    .S(_21849_),
    .Z(_02176_));
 MUX2_X1 _50807_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2220]),
    .B(_21773_),
    .S(_21849_),
    .Z(_02178_));
 MUX2_X1 _50808_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2221]),
    .B(_21805_),
    .S(_21849_),
    .Z(_02179_));
 MUX2_X1 _50809_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2222]),
    .B(_21516_),
    .S(_21849_),
    .Z(_02180_));
 BUF_X16 _50810_ (.A(_21846_),
    .Z(_21853_));
 MUX2_X1 _50811_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2223]),
    .B(_21807_),
    .S(_21853_),
    .Z(_02181_));
 MUX2_X1 _50812_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2224]),
    .B(_21777_),
    .S(_21853_),
    .Z(_02182_));
 NAND4_X1 _50813_ (.A1(_21640_),
    .A2(_10614_),
    .A3(_21821_),
    .A4(_21828_),
    .ZN(_21854_));
 INV_X1 _50814_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2225]),
    .ZN(_21855_));
 OAI21_X1 _50815_ (.A(_21854_),
    .B1(_21848_),
    .B2(_21855_),
    .ZN(_02183_));
 MUX2_X1 _50816_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2226]),
    .B(_21779_),
    .S(_21853_),
    .Z(_02184_));
 MUX2_X1 _50817_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2227]),
    .B(_21780_),
    .S(_21853_),
    .Z(_02185_));
 MUX2_X1 _50818_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2228]),
    .B(_21588_),
    .S(_21853_),
    .Z(_02186_));
 MUX2_X1 _50819_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2229]),
    .B(_21837_),
    .S(_21853_),
    .Z(_02187_));
 MUX2_X1 _50820_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2230]),
    .B(_21617_),
    .S(_21853_),
    .Z(_02189_));
 MUX2_X1 _50821_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2231]),
    .B(_21783_),
    .S(_21853_),
    .Z(_02190_));
 BUF_X16 _50822_ (.A(_10784_),
    .Z(_21856_));
 BUF_X4 _50823_ (.A(_21856_),
    .Z(_21857_));
 NAND4_X1 _50824_ (.A1(_21640_),
    .A2(_21520_),
    .A3(_21857_),
    .A4(_21828_),
    .ZN(_21858_));
 INV_X1 _50825_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2232]),
    .ZN(_21859_));
 OAI21_X1 _50826_ (.A(_21858_),
    .B1(_21848_),
    .B2(_21859_),
    .ZN(_02191_));
 MUX2_X1 _50827_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2233]),
    .B(_21555_),
    .S(_21853_),
    .Z(_02192_));
 BUF_X8 _50828_ (.A(_08608_),
    .Z(_21860_));
 MUX2_X1 _50829_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2234]),
    .B(_21860_),
    .S(_21853_),
    .Z(_02193_));
 BUF_X16 _50830_ (.A(_21846_),
    .Z(_21861_));
 MUX2_X1 _50831_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2235]),
    .B(_21490_),
    .S(_21861_),
    .Z(_02194_));
 BUF_X8 _50832_ (.A(_08614_),
    .Z(_21862_));
 MUX2_X1 _50833_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2236]),
    .B(_21862_),
    .S(_21861_),
    .Z(_02195_));
 MUX2_X1 _50834_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2237]),
    .B(_21792_),
    .S(_21861_),
    .Z(_02196_));
 MUX2_X1 _50835_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2238]),
    .B(_21793_),
    .S(_21861_),
    .Z(_02197_));
 MUX2_X1 _50836_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2239]),
    .B(_21621_),
    .S(_21861_),
    .Z(_02198_));
 MUX2_X1 _50837_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2240]),
    .B(_21794_),
    .S(_21861_),
    .Z(_02200_));
 MUX2_X1 _50838_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2241]),
    .B(_21795_),
    .S(_21861_),
    .Z(_02201_));
 MUX2_X1 _50839_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2242]),
    .B(_21843_),
    .S(_21861_),
    .Z(_02202_));
 MUX2_X1 _50840_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2243]),
    .B(_21498_),
    .S(_21861_),
    .Z(_02203_));
 MUX2_X1 _50841_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2244]),
    .B(_21762_),
    .S(_21861_),
    .Z(_02204_));
 MUX2_X1 _50842_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2245]),
    .B(_21649_),
    .S(_21847_),
    .Z(_02205_));
 MUX2_X1 _50843_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2246]),
    .B(_21766_),
    .S(_21847_),
    .Z(_02206_));
 MUX2_X1 _50844_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2247]),
    .B(_21737_),
    .S(_21847_),
    .Z(_02207_));
 MUX2_X1 _50845_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2248]),
    .B(_21815_),
    .S(_21847_),
    .Z(_02208_));
 MUX2_X1 _50846_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2249]),
    .B(_21703_),
    .S(_21847_),
    .Z(_02209_));
 MUX2_X1 _50847_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2250]),
    .B(_21652_),
    .S(_21847_),
    .Z(_02211_));
 MUX2_X1 _50848_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2251]),
    .B(_21678_),
    .S(_21847_),
    .Z(_02212_));
 MUX2_X1 _50849_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2252]),
    .B(_21653_),
    .S(_21847_),
    .Z(_02213_));
 MUX2_X1 _50850_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2253]),
    .B(_21704_),
    .S(_21847_),
    .Z(_02214_));
 BUF_X8 _50851_ (.A(_21598_),
    .Z(_21863_));
 AND2_X4 _50852_ (.A1(_10955_),
    .A2(_21574_),
    .ZN(_21864_));
 BUF_X16 _50853_ (.A(_21864_),
    .Z(_21865_));
 BUF_X8 _50854_ (.A(_21865_),
    .Z(_21866_));
 MUX2_X1 _50855_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2156]),
    .B(_21863_),
    .S(_21866_),
    .Z(_02106_));
 BUF_X8 _50856_ (.A(_21605_),
    .Z(_21867_));
 MUX2_X1 _50857_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2157]),
    .B(_21867_),
    .S(_21866_),
    .Z(_02107_));
 MUX2_X1 _50858_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2158]),
    .B(_21683_),
    .S(_21866_),
    .Z(_02108_));
 BUF_X4 _50859_ (.A(_21608_),
    .Z(_21868_));
 MUX2_X1 _50860_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2159]),
    .B(_21868_),
    .S(_21866_),
    .Z(_02109_));
 MUX2_X1 _50861_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2160]),
    .B(_21684_),
    .S(_21866_),
    .Z(_02111_));
 MUX2_X1 _50862_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2161]),
    .B(_21635_),
    .S(_21866_),
    .Z(_02112_));
 BUF_X8 _50863_ (.A(_21864_),
    .Z(_21869_));
 MUX2_X1 _50864_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2162]),
    .B(_21745_),
    .S(_21869_),
    .Z(_02113_));
 MUX2_X1 _50865_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2163]),
    .B(_21688_),
    .S(_21869_),
    .Z(_02114_));
 MUX2_X1 _50866_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2164]),
    .B(_21689_),
    .S(_21869_),
    .Z(_02115_));
 MUX2_X1 _50867_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2165]),
    .B(_21749_),
    .S(_21869_),
    .Z(_02116_));
 MUX2_X1 _50868_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2166]),
    .B(_21714_),
    .S(_21869_),
    .Z(_02117_));
 MUX2_X1 _50869_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2167]),
    .B(_21750_),
    .S(_21869_),
    .Z(_02118_));
 MUX2_X1 _50870_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2168]),
    .B(_21833_),
    .S(_21869_),
    .Z(_02119_));
 MUX2_X1 _50871_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2169]),
    .B(_21852_),
    .S(_21869_),
    .Z(_02120_));
 MUX2_X1 _50872_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2170]),
    .B(_21804_),
    .S(_21869_),
    .Z(_02122_));
 MUX2_X1 _50873_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2171]),
    .B(_21773_),
    .S(_21869_),
    .Z(_02123_));
 BUF_X16 _50874_ (.A(_21864_),
    .Z(_21870_));
 MUX2_X1 _50875_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2172]),
    .B(_21805_),
    .S(_21870_),
    .Z(_02124_));
 MUX2_X1 _50876_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2173]),
    .B(_21516_),
    .S(_21870_),
    .Z(_02125_));
 MUX2_X1 _50877_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2174]),
    .B(_21807_),
    .S(_21870_),
    .Z(_02126_));
 MUX2_X1 _50878_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2175]),
    .B(_21777_),
    .S(_21870_),
    .Z(_02127_));
 NAND4_X1 _50879_ (.A1(_21672_),
    .A2(_10614_),
    .A3(_21857_),
    .A4(_21828_),
    .ZN(_21871_));
 INV_X1 _50880_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2176]),
    .ZN(_21872_));
 OAI21_X1 _50881_ (.A(_21871_),
    .B1(_21866_),
    .B2(_21872_),
    .ZN(_02128_));
 MUX2_X1 _50882_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2177]),
    .B(_21779_),
    .S(_21870_),
    .Z(_02129_));
 MUX2_X1 _50883_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2178]),
    .B(_21780_),
    .S(_21870_),
    .Z(_02130_));
 MUX2_X1 _50884_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2179]),
    .B(_21588_),
    .S(_21870_),
    .Z(_02131_));
 MUX2_X1 _50885_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2180]),
    .B(_21837_),
    .S(_21870_),
    .Z(_02133_));
 MUX2_X1 _50886_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2181]),
    .B(_21617_),
    .S(_21870_),
    .Z(_02134_));
 MUX2_X1 _50887_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2182]),
    .B(_21783_),
    .S(_21870_),
    .Z(_02135_));
 NAND4_X1 _50888_ (.A1(_21672_),
    .A2(_21520_),
    .A3(_21857_),
    .A4(_21828_),
    .ZN(_21873_));
 INV_X1 _50889_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2183]),
    .ZN(_21874_));
 OAI21_X1 _50890_ (.A(_21873_),
    .B1(_21866_),
    .B2(_21874_),
    .ZN(_02136_));
 BUF_X16 _50891_ (.A(_21864_),
    .Z(_21875_));
 MUX2_X1 _50892_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2184]),
    .B(_21555_),
    .S(_21875_),
    .Z(_02137_));
 BUF_X8 _50893_ (.A(_10942_),
    .Z(_21876_));
 NAND4_X1 _50894_ (.A1(_21672_),
    .A2(_10616_),
    .A3(_21857_),
    .A4(_21876_),
    .ZN(_21877_));
 INV_X1 _50895_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2185]),
    .ZN(_21878_));
 OAI21_X1 _50896_ (.A(_21877_),
    .B1(_21866_),
    .B2(_21878_),
    .ZN(_02138_));
 MUX2_X1 _50897_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2186]),
    .B(_21490_),
    .S(_21875_),
    .Z(_02139_));
 MUX2_X1 _50898_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2187]),
    .B(_21862_),
    .S(_21875_),
    .Z(_02140_));
 MUX2_X1 _50899_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2188]),
    .B(_21792_),
    .S(_21875_),
    .Z(_02141_));
 MUX2_X1 _50900_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2189]),
    .B(_21793_),
    .S(_21875_),
    .Z(_02142_));
 BUF_X8 _50901_ (.A(_08623_),
    .Z(_21879_));
 MUX2_X1 _50902_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2190]),
    .B(_21879_),
    .S(_21875_),
    .Z(_02144_));
 MUX2_X1 _50903_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2191]),
    .B(_21794_),
    .S(_21875_),
    .Z(_02145_));
 NAND4_X4 _50904_ (.A1(_21672_),
    .A2(_10593_),
    .A3(_21857_),
    .A4(_21876_),
    .ZN(_21880_));
 INV_X1 _50905_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2192]),
    .ZN(_21881_));
 OAI21_X1 _50906_ (.A(_21880_),
    .B1(_21866_),
    .B2(_21881_),
    .ZN(_02146_));
 MUX2_X1 _50907_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2193]),
    .B(_21843_),
    .S(_21875_),
    .Z(_02147_));
 MUX2_X1 _50908_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2194]),
    .B(_21498_),
    .S(_21875_),
    .Z(_02148_));
 MUX2_X1 _50909_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2195]),
    .B(_21762_),
    .S(_21875_),
    .Z(_02149_));
 MUX2_X1 _50910_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2196]),
    .B(_21649_),
    .S(_21865_),
    .Z(_02150_));
 MUX2_X1 _50911_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2197]),
    .B(_21766_),
    .S(_21865_),
    .Z(_02151_));
 MUX2_X1 _50912_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2198]),
    .B(_21737_),
    .S(_21865_),
    .Z(_02152_));
 MUX2_X1 _50913_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2199]),
    .B(_21815_),
    .S(_21865_),
    .Z(_02153_));
 MUX2_X1 _50914_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2200]),
    .B(_21703_),
    .S(_21865_),
    .Z(_02156_));
 MUX2_X1 _50915_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2201]),
    .B(_21652_),
    .S(_21865_),
    .Z(_02157_));
 MUX2_X1 _50916_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2202]),
    .B(_21678_),
    .S(_21865_),
    .Z(_02158_));
 MUX2_X1 _50917_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2203]),
    .B(_21653_),
    .S(_21865_),
    .Z(_02159_));
 MUX2_X1 _50918_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2204]),
    .B(_21704_),
    .S(_21865_),
    .Z(_02160_));
 AND2_X4 _50919_ (.A1(_10961_),
    .A2(_21574_),
    .ZN(_21882_));
 BUF_X16 _50920_ (.A(_21882_),
    .Z(_21883_));
 BUF_X8 _50921_ (.A(_21883_),
    .Z(_21884_));
 MUX2_X1 _50922_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2107]),
    .B(_21863_),
    .S(_21884_),
    .Z(_02052_));
 MUX2_X1 _50923_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2108]),
    .B(_21867_),
    .S(_21884_),
    .Z(_02053_));
 MUX2_X1 _50924_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2109]),
    .B(_21683_),
    .S(_21884_),
    .Z(_02054_));
 MUX2_X1 _50925_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2110]),
    .B(_21868_),
    .S(_21884_),
    .Z(_02056_));
 MUX2_X1 _50926_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2111]),
    .B(_21684_),
    .S(_21884_),
    .Z(_02057_));
 BUF_X8 _50927_ (.A(_21299_),
    .Z(_21885_));
 MUX2_X1 _50928_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2112]),
    .B(_21885_),
    .S(_21884_),
    .Z(_02058_));
 BUF_X8 _50929_ (.A(_21882_),
    .Z(_21886_));
 MUX2_X1 _50930_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2113]),
    .B(_21745_),
    .S(_21886_),
    .Z(_02059_));
 MUX2_X1 _50931_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2114]),
    .B(_21688_),
    .S(_21886_),
    .Z(_02060_));
 MUX2_X1 _50932_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2115]),
    .B(_21689_),
    .S(_21886_),
    .Z(_02061_));
 MUX2_X1 _50933_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2116]),
    .B(_21749_),
    .S(_21886_),
    .Z(_02062_));
 MUX2_X1 _50934_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2117]),
    .B(_21714_),
    .S(_21886_),
    .Z(_02063_));
 MUX2_X1 _50935_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2118]),
    .B(_21750_),
    .S(_21886_),
    .Z(_02064_));
 MUX2_X1 _50936_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2119]),
    .B(_21833_),
    .S(_21886_),
    .Z(_02065_));
 MUX2_X1 _50937_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2120]),
    .B(_21852_),
    .S(_21886_),
    .Z(_02067_));
 MUX2_X1 _50938_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2121]),
    .B(_21804_),
    .S(_21886_),
    .Z(_02068_));
 MUX2_X1 _50939_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2122]),
    .B(_21773_),
    .S(_21886_),
    .Z(_02069_));
 BUF_X8 _50940_ (.A(_21882_),
    .Z(_21887_));
 MUX2_X1 _50941_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2123]),
    .B(_21805_),
    .S(_21887_),
    .Z(_02070_));
 NAND4_X1 _50942_ (.A1(_21486_),
    .A2(_10599_),
    .A3(_21857_),
    .A4(_21876_),
    .ZN(_21888_));
 INV_X1 _50943_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2124]),
    .ZN(_21889_));
 OAI21_X1 _50944_ (.A(_21888_),
    .B1(_21884_),
    .B2(_21889_),
    .ZN(_02071_));
 MUX2_X1 _50945_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2125]),
    .B(_21807_),
    .S(_21887_),
    .Z(_02072_));
 MUX2_X1 _50946_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2126]),
    .B(_21777_),
    .S(_21887_),
    .Z(_02073_));
 BUF_X8 _50947_ (.A(_10781_),
    .Z(_21890_));
 NAND4_X1 _50948_ (.A1(_21890_),
    .A2(_10614_),
    .A3(_21857_),
    .A4(_21876_),
    .ZN(_21891_));
 INV_X1 _50949_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2127]),
    .ZN(_21892_));
 OAI21_X1 _50950_ (.A(_21891_),
    .B1(_21884_),
    .B2(_21892_),
    .ZN(_02074_));
 MUX2_X1 _50951_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2128]),
    .B(_21779_),
    .S(_21887_),
    .Z(_02075_));
 MUX2_X1 _50952_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2129]),
    .B(_21780_),
    .S(_21887_),
    .Z(_02076_));
 MUX2_X1 _50953_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2130]),
    .B(_21588_),
    .S(_21887_),
    .Z(_02078_));
 MUX2_X1 _50954_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2131]),
    .B(_21837_),
    .S(_21887_),
    .Z(_02079_));
 MUX2_X1 _50955_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2132]),
    .B(_21617_),
    .S(_21887_),
    .Z(_02080_));
 MUX2_X1 _50956_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2133]),
    .B(_21783_),
    .S(_21887_),
    .Z(_02081_));
 NAND4_X1 _50957_ (.A1(_21890_),
    .A2(_21520_),
    .A3(_21857_),
    .A4(_21876_),
    .ZN(_21893_));
 INV_X1 _50958_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2134]),
    .ZN(_21894_));
 OAI21_X1 _50959_ (.A(_21893_),
    .B1(_21884_),
    .B2(_21894_),
    .ZN(_02082_));
 MUX2_X1 _50960_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2135]),
    .B(_21555_),
    .S(_21887_),
    .Z(_02083_));
 NAND4_X1 _50961_ (.A1(_21890_),
    .A2(_10616_),
    .A3(_21857_),
    .A4(_21876_),
    .ZN(_21895_));
 INV_X1 _50962_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2136]),
    .ZN(_21896_));
 OAI21_X1 _50963_ (.A(_21895_),
    .B1(_21884_),
    .B2(_21896_),
    .ZN(_02084_));
 BUF_X16 _50964_ (.A(_21882_),
    .Z(_21897_));
 MUX2_X1 _50965_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2137]),
    .B(_21490_),
    .S(_21897_),
    .Z(_02085_));
 MUX2_X1 _50966_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2138]),
    .B(_21862_),
    .S(_21897_),
    .Z(_02086_));
 MUX2_X1 _50967_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2139]),
    .B(_21792_),
    .S(_21897_),
    .Z(_02087_));
 MUX2_X1 _50968_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2140]),
    .B(_21793_),
    .S(_21897_),
    .Z(_02089_));
 MUX2_X1 _50969_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2141]),
    .B(_21879_),
    .S(_21897_),
    .Z(_02090_));
 MUX2_X1 _50970_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2142]),
    .B(_21794_),
    .S(_21897_),
    .Z(_02091_));
 MUX2_X1 _50971_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2143]),
    .B(_21795_),
    .S(_21897_),
    .Z(_02092_));
 MUX2_X1 _50972_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2144]),
    .B(_21843_),
    .S(_21897_),
    .Z(_02093_));
 MUX2_X1 _50973_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2145]),
    .B(_21498_),
    .S(_21897_),
    .Z(_02094_));
 MUX2_X1 _50974_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2146]),
    .B(_21762_),
    .S(_21897_),
    .Z(_02095_));
 MUX2_X1 _50975_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2147]),
    .B(_21649_),
    .S(_21883_),
    .Z(_02096_));
 MUX2_X1 _50976_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2148]),
    .B(_21766_),
    .S(_21883_),
    .Z(_02097_));
 MUX2_X1 _50977_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2149]),
    .B(_21737_),
    .S(_21883_),
    .Z(_02098_));
 MUX2_X1 _50978_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2150]),
    .B(_21815_),
    .S(_21883_),
    .Z(_02100_));
 MUX2_X1 _50979_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2151]),
    .B(_21703_),
    .S(_21883_),
    .Z(_02101_));
 BUF_X8 _50980_ (.A(_21365_),
    .Z(_21898_));
 MUX2_X1 _50981_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2152]),
    .B(_21898_),
    .S(_21883_),
    .Z(_02102_));
 MUX2_X1 _50982_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2153]),
    .B(_21678_),
    .S(_21883_),
    .Z(_02103_));
 BUF_X16 _50983_ (.A(_21373_),
    .Z(_21899_));
 MUX2_X1 _50984_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2154]),
    .B(_21899_),
    .S(_21883_),
    .Z(_02104_));
 MUX2_X1 _50985_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2155]),
    .B(_21704_),
    .S(_21883_),
    .Z(_02105_));
 BUF_X16 _50986_ (.A(_10968_),
    .Z(_21900_));
 AND2_X4 _50987_ (.A1(_21900_),
    .A2(_10784_),
    .ZN(_21901_));
 BUF_X16 _50988_ (.A(_21901_),
    .Z(_21902_));
 MUX2_X1 _50989_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2058]),
    .B(_21863_),
    .S(_21902_),
    .Z(_01997_));
 MUX2_X1 _50990_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2059]),
    .B(_21867_),
    .S(_21902_),
    .Z(_01998_));
 MUX2_X1 _50991_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2060]),
    .B(_21683_),
    .S(_21902_),
    .Z(_02000_));
 MUX2_X1 _50992_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2061]),
    .B(_21868_),
    .S(_21902_),
    .Z(_02001_));
 MUX2_X1 _50993_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2062]),
    .B(_21684_),
    .S(_21902_),
    .Z(_02002_));
 MUX2_X1 _50994_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2063]),
    .B(_21885_),
    .S(_21902_),
    .Z(_02003_));
 MUX2_X1 _50995_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2064]),
    .B(_21745_),
    .S(_21902_),
    .Z(_02004_));
 MUX2_X1 _50996_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2065]),
    .B(_21688_),
    .S(_21902_),
    .Z(_02005_));
 BUF_X16 _50997_ (.A(_21901_),
    .Z(_21903_));
 MUX2_X1 _50998_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2066]),
    .B(_21689_),
    .S(_21903_),
    .Z(_02006_));
 MUX2_X1 _50999_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2067]),
    .B(_21749_),
    .S(_21903_),
    .Z(_02007_));
 MUX2_X1 _51000_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2068]),
    .B(_21714_),
    .S(_21903_),
    .Z(_02008_));
 MUX2_X1 _51001_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2069]),
    .B(_21750_),
    .S(_21903_),
    .Z(_02009_));
 NAND4_X2 _51002_ (.A1(_21716_),
    .A2(_10563_),
    .A3(_21857_),
    .A4(_21876_),
    .ZN(_21904_));
 BUF_X4 _51003_ (.A(_21902_),
    .Z(_21905_));
 INV_X1 _51004_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2070]),
    .ZN(_21906_));
 OAI21_X1 _51005_ (.A(_21904_),
    .B1(_21905_),
    .B2(_21906_),
    .ZN(_02011_));
 BUF_X4 _51006_ (.A(_10859_),
    .Z(_21907_));
 BUF_X4 _51007_ (.A(_21856_),
    .Z(_21908_));
 NAND4_X1 _51008_ (.A1(_21907_),
    .A2(_08555_),
    .A3(_21908_),
    .A4(_21876_),
    .ZN(_21909_));
 INV_X1 _51009_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2071]),
    .ZN(_21910_));
 OAI21_X1 _51010_ (.A(_21909_),
    .B1(_21905_),
    .B2(_21910_),
    .ZN(_02012_));
 MUX2_X1 _51011_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2072]),
    .B(_21804_),
    .S(_21903_),
    .Z(_02013_));
 NAND4_X1 _51012_ (.A1(_21907_),
    .A2(_10571_),
    .A3(_21908_),
    .A4(_21876_),
    .ZN(_21911_));
 INV_X1 _51013_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2073]),
    .ZN(_21912_));
 OAI21_X1 _51014_ (.A(_21911_),
    .B1(_21905_),
    .B2(_21912_),
    .ZN(_02014_));
 MUX2_X1 _51015_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2074]),
    .B(_21805_),
    .S(_21903_),
    .Z(_02015_));
 NAND4_X1 _51016_ (.A1(_21907_),
    .A2(_10599_),
    .A3(_21908_),
    .A4(_21876_),
    .ZN(_21913_));
 INV_X1 _51017_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2075]),
    .ZN(_21914_));
 OAI21_X1 _51018_ (.A(_21913_),
    .B1(_21905_),
    .B2(_21914_),
    .ZN(_02016_));
 MUX2_X1 _51019_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2076]),
    .B(_21807_),
    .S(_21903_),
    .Z(_02017_));
 MUX2_X1 _51020_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2077]),
    .B(_21777_),
    .S(_21903_),
    .Z(_02018_));
 MUX2_X1 _51021_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2078]),
    .B(_21778_),
    .S(_21903_),
    .Z(_02019_));
 MUX2_X1 _51022_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2079]),
    .B(_21779_),
    .S(_21903_),
    .Z(_02020_));
 BUF_X16 _51023_ (.A(_21901_),
    .Z(_21915_));
 MUX2_X1 _51024_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2080]),
    .B(_21780_),
    .S(_21915_),
    .Z(_02022_));
 BUF_X4 _51025_ (.A(_10942_),
    .Z(_21916_));
 NAND4_X1 _51026_ (.A1(_21907_),
    .A2(_08588_),
    .A3(_21908_),
    .A4(_21916_),
    .ZN(_21917_));
 INV_X1 _51027_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2081]),
    .ZN(_21918_));
 OAI21_X1 _51028_ (.A(_21917_),
    .B1(_21905_),
    .B2(_21918_),
    .ZN(_02023_));
 MUX2_X1 _51029_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2082]),
    .B(_21837_),
    .S(_21915_),
    .Z(_02024_));
 BUF_X16 _51030_ (.A(_08594_),
    .Z(_21919_));
 MUX2_X1 _51031_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2083]),
    .B(_21919_),
    .S(_21915_),
    .Z(_02025_));
 MUX2_X1 _51032_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2084]),
    .B(_21783_),
    .S(_21915_),
    .Z(_02026_));
 NAND4_X1 _51033_ (.A1(_21907_),
    .A2(_21520_),
    .A3(_21908_),
    .A4(_21916_),
    .ZN(_21920_));
 INV_X1 _51034_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2085]),
    .ZN(_21921_));
 OAI21_X1 _51035_ (.A(_21920_),
    .B1(_21905_),
    .B2(_21921_),
    .ZN(_02027_));
 NAND4_X1 _51036_ (.A1(_21907_),
    .A2(_21725_),
    .A3(_21908_),
    .A4(_21916_),
    .ZN(_21922_));
 INV_X1 _51037_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2086]),
    .ZN(_21923_));
 OAI21_X1 _51038_ (.A(_21922_),
    .B1(_21905_),
    .B2(_21923_),
    .ZN(_02028_));
 NAND4_X1 _51039_ (.A1(_21907_),
    .A2(_10616_),
    .A3(_21908_),
    .A4(_21916_),
    .ZN(_21924_));
 INV_X1 _51040_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2087]),
    .ZN(_21925_));
 OAI21_X1 _51041_ (.A(_21924_),
    .B1(_21905_),
    .B2(_21925_),
    .ZN(_02029_));
 MUX2_X1 _51042_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2088]),
    .B(_21490_),
    .S(_21915_),
    .Z(_02030_));
 MUX2_X1 _51043_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2089]),
    .B(_21862_),
    .S(_21915_),
    .Z(_02031_));
 MUX2_X1 _51044_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2090]),
    .B(_21792_),
    .S(_21915_),
    .Z(_02033_));
 MUX2_X1 _51045_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2091]),
    .B(_21793_),
    .S(_21915_),
    .Z(_02034_));
 NAND4_X1 _51046_ (.A1(_21907_),
    .A2(_21562_),
    .A3(_21908_),
    .A4(_21916_),
    .ZN(_21926_));
 INV_X1 _51047_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2092]),
    .ZN(_21927_));
 OAI21_X1 _51048_ (.A(_21926_),
    .B1(_21905_),
    .B2(_21927_),
    .ZN(_02035_));
 MUX2_X1 _51049_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2093]),
    .B(_21794_),
    .S(_21915_),
    .Z(_02036_));
 MUX2_X1 _51050_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2094]),
    .B(_21795_),
    .S(_21915_),
    .Z(_02037_));
 NAND4_X1 _51051_ (.A1(_21907_),
    .A2(_21330_),
    .A3(_21908_),
    .A4(_21916_),
    .ZN(_21928_));
 INV_X1 _51052_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2095]),
    .ZN(_21929_));
 OAI21_X1 _51053_ (.A(_21928_),
    .B1(_21905_),
    .B2(_21929_),
    .ZN(_02038_));
 BUF_X8 _51054_ (.A(_08635_),
    .Z(_21930_));
 BUF_X16 _51055_ (.A(_21901_),
    .Z(_21931_));
 MUX2_X1 _51056_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2096]),
    .B(_21930_),
    .S(_21931_),
    .Z(_02039_));
 MUX2_X1 _51057_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2097]),
    .B(_21762_),
    .S(_21931_),
    .Z(_02040_));
 BUF_X8 _51058_ (.A(_21343_),
    .Z(_21932_));
 MUX2_X1 _51059_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2098]),
    .B(_21932_),
    .S(_21931_),
    .Z(_02041_));
 MUX2_X1 _51060_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2099]),
    .B(_21766_),
    .S(_21931_),
    .Z(_02042_));
 MUX2_X1 _51061_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2100]),
    .B(_21737_),
    .S(_21931_),
    .Z(_02045_));
 MUX2_X1 _51062_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2101]),
    .B(_21815_),
    .S(_21931_),
    .Z(_02046_));
 MUX2_X1 _51063_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2102]),
    .B(_21703_),
    .S(_21931_),
    .Z(_02047_));
 MUX2_X1 _51064_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2103]),
    .B(_21898_),
    .S(_21931_),
    .Z(_02048_));
 BUF_X8 _51065_ (.A(_21369_),
    .Z(_21933_));
 MUX2_X1 _51066_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2104]),
    .B(_21933_),
    .S(_21931_),
    .Z(_02049_));
 BUF_X8 _51067_ (.A(_11015_),
    .Z(_21934_));
 NAND4_X1 _51068_ (.A1(_21907_),
    .A2(_21934_),
    .A3(_21800_),
    .A4(_21373_),
    .ZN(_21935_));
 INV_X1 _51069_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2105]),
    .ZN(_21936_));
 OAI21_X1 _51070_ (.A(_21935_),
    .B1(_21902_),
    .B2(_21936_),
    .ZN(_02050_));
 MUX2_X1 _51071_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2106]),
    .B(_21704_),
    .S(_21931_),
    .Z(_02051_));
 BUF_X16 _51072_ (.A(_10972_),
    .Z(_21937_));
 AND2_X4 _51073_ (.A1(_21937_),
    .A2(_21441_),
    .ZN(_21938_));
 BUF_X16 _51074_ (.A(_21938_),
    .Z(_21939_));
 BUF_X8 _51075_ (.A(_21939_),
    .Z(_21940_));
 MUX2_X1 _51076_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2009]),
    .B(_21863_),
    .S(_21940_),
    .Z(_01943_));
 MUX2_X1 _51077_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2010]),
    .B(_21867_),
    .S(_21940_),
    .Z(_01945_));
 MUX2_X1 _51078_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2011]),
    .B(_21683_),
    .S(_21940_),
    .Z(_01946_));
 BUF_X16 _51079_ (.A(_21938_),
    .Z(_21941_));
 MUX2_X1 _51080_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2012]),
    .B(_21868_),
    .S(_21941_),
    .Z(_01947_));
 MUX2_X1 _51081_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2013]),
    .B(_21684_),
    .S(_21941_),
    .Z(_01948_));
 MUX2_X1 _51082_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2014]),
    .B(_21885_),
    .S(_21941_),
    .Z(_01949_));
 MUX2_X1 _51083_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2015]),
    .B(_21745_),
    .S(_21941_),
    .Z(_01950_));
 NAND4_X4 _51084_ (.A1(_21752_),
    .A2(_21582_),
    .A3(_21908_),
    .A4(_21916_),
    .ZN(_21942_));
 INV_X1 _51085_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2016]),
    .ZN(_21943_));
 OAI21_X1 _51086_ (.A(_21942_),
    .B1(_21940_),
    .B2(_21943_),
    .ZN(_01951_));
 MUX2_X1 _51087_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2017]),
    .B(_21689_),
    .S(_21941_),
    .Z(_01952_));
 MUX2_X1 _51088_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2018]),
    .B(_21749_),
    .S(_21941_),
    .Z(_01953_));
 MUX2_X1 _51089_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2019]),
    .B(_21714_),
    .S(_21941_),
    .Z(_01954_));
 MUX2_X1 _51090_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2020]),
    .B(_21750_),
    .S(_21941_),
    .Z(_01956_));
 MUX2_X1 _51091_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2021]),
    .B(_21833_),
    .S(_21941_),
    .Z(_01957_));
 MUX2_X1 _51092_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2022]),
    .B(_21852_),
    .S(_21941_),
    .Z(_01958_));
 BUF_X16 _51093_ (.A(_21938_),
    .Z(_21944_));
 MUX2_X1 _51094_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2023]),
    .B(_21804_),
    .S(_21944_),
    .Z(_01959_));
 BUF_X8 _51095_ (.A(_21856_),
    .Z(_21945_));
 NAND4_X1 _51096_ (.A1(_21752_),
    .A2(_10571_),
    .A3(_21945_),
    .A4(_21916_),
    .ZN(_21946_));
 INV_X1 _51097_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2024]),
    .ZN(_21947_));
 OAI21_X1 _51098_ (.A(_21946_),
    .B1(_21940_),
    .B2(_21947_),
    .ZN(_01960_));
 MUX2_X1 _51099_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2025]),
    .B(_21805_),
    .S(_21944_),
    .Z(_01961_));
 BUF_X8 _51100_ (.A(_08567_),
    .Z(_21948_));
 MUX2_X1 _51101_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2026]),
    .B(_21948_),
    .S(_21944_),
    .Z(_01962_));
 MUX2_X1 _51102_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2027]),
    .B(_21807_),
    .S(_21944_),
    .Z(_01963_));
 MUX2_X1 _51103_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2028]),
    .B(_21777_),
    .S(_21944_),
    .Z(_01964_));
 MUX2_X1 _51104_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2029]),
    .B(_21778_),
    .S(_21944_),
    .Z(_01965_));
 MUX2_X1 _51105_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2030]),
    .B(_21779_),
    .S(_21944_),
    .Z(_01967_));
 MUX2_X1 _51106_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2031]),
    .B(_21780_),
    .S(_21944_),
    .Z(_01968_));
 MUX2_X1 _51107_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2032]),
    .B(_21588_),
    .S(_21944_),
    .Z(_01969_));
 MUX2_X1 _51108_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2033]),
    .B(_21837_),
    .S(_21944_),
    .Z(_01970_));
 NAND4_X2 _51109_ (.A1(_21752_),
    .A2(_21757_),
    .A3(_21945_),
    .A4(_21916_),
    .ZN(_21949_));
 INV_X1 _51110_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2034]),
    .ZN(_21950_));
 OAI21_X1 _51111_ (.A(_21949_),
    .B1(_21940_),
    .B2(_21950_),
    .ZN(_01971_));
 BUF_X16 _51112_ (.A(_21938_),
    .Z(_21951_));
 MUX2_X1 _51113_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2035]),
    .B(_21783_),
    .S(_21951_),
    .Z(_01972_));
 BUF_X16 _51114_ (.A(_08600_),
    .Z(_21952_));
 MUX2_X1 _51115_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2036]),
    .B(_21952_),
    .S(_21951_),
    .Z(_01973_));
 NAND4_X1 _51116_ (.A1(_21752_),
    .A2(_21725_),
    .A3(_21945_),
    .A4(_21916_),
    .ZN(_21953_));
 INV_X1 _51117_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2037]),
    .ZN(_21954_));
 OAI21_X1 _51118_ (.A(_21953_),
    .B1(_21940_),
    .B2(_21954_),
    .ZN(_01974_));
 MUX2_X1 _51119_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2038]),
    .B(_21860_),
    .S(_21951_),
    .Z(_01975_));
 BUF_X16 _51120_ (.A(_08611_),
    .Z(_21955_));
 MUX2_X1 _51121_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2039]),
    .B(_21955_),
    .S(_21951_),
    .Z(_01976_));
 MUX2_X1 _51122_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2040]),
    .B(_21862_),
    .S(_21951_),
    .Z(_01978_));
 MUX2_X1 _51123_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2041]),
    .B(_21792_),
    .S(_21951_),
    .Z(_01979_));
 MUX2_X1 _51124_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2042]),
    .B(_21793_),
    .S(_21951_),
    .Z(_01980_));
 MUX2_X1 _51125_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2043]),
    .B(_21879_),
    .S(_21951_),
    .Z(_01981_));
 MUX2_X1 _51126_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2044]),
    .B(_21794_),
    .S(_21951_),
    .Z(_01982_));
 MUX2_X1 _51127_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2045]),
    .B(_21795_),
    .S(_21951_),
    .Z(_01983_));
 MUX2_X1 _51128_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2046]),
    .B(_21843_),
    .S(_21939_),
    .Z(_01984_));
 MUX2_X1 _51129_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2047]),
    .B(_21930_),
    .S(_21939_),
    .Z(_01985_));
 NAND4_X4 _51130_ (.A1(_21752_),
    .A2(_21934_),
    .A3(_21800_),
    .A4(_21595_),
    .ZN(_21956_));
 INV_X1 _51131_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2048]),
    .ZN(_21957_));
 OAI21_X1 _51132_ (.A(_21956_),
    .B1(_21940_),
    .B2(_21957_),
    .ZN(_01986_));
 MUX2_X1 _51133_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2049]),
    .B(_21932_),
    .S(_21939_),
    .Z(_01987_));
 MUX2_X1 _51134_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2050]),
    .B(_21766_),
    .S(_21939_),
    .Z(_01989_));
 MUX2_X1 _51135_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2051]),
    .B(_21737_),
    .S(_21939_),
    .Z(_01990_));
 MUX2_X1 _51136_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2052]),
    .B(_21815_),
    .S(_21939_),
    .Z(_01991_));
 BUF_X8 _51137_ (.A(_21359_),
    .Z(_21958_));
 MUX2_X1 _51138_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2053]),
    .B(_21958_),
    .S(_21939_),
    .Z(_01992_));
 MUX2_X1 _51139_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2054]),
    .B(_21898_),
    .S(_21939_),
    .Z(_01993_));
 NAND4_X1 _51140_ (.A1(_21752_),
    .A2(_21934_),
    .A3(_21800_),
    .A4(_21369_),
    .ZN(_21959_));
 INV_X4 _51141_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2055]),
    .ZN(_21960_));
 OAI21_X1 _51142_ (.A(_21959_),
    .B1(_21940_),
    .B2(_21960_),
    .ZN(_01994_));
 BUF_X16 _51143_ (.A(_10869_),
    .Z(_21961_));
 NAND4_X1 _51144_ (.A1(_21961_),
    .A2(_21934_),
    .A3(_21800_),
    .A4(_21373_),
    .ZN(_21962_));
 INV_X1 _51145_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2056]),
    .ZN(_21963_));
 OAI21_X1 _51146_ (.A(_21962_),
    .B1(_21940_),
    .B2(_21963_),
    .ZN(_01995_));
 MUX2_X1 _51147_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2057]),
    .B(_21704_),
    .S(_21939_),
    .Z(_01996_));
 AND2_X4 _51148_ (.A1(_10976_),
    .A2(_21432_),
    .ZN(_21964_));
 BUF_X16 _51149_ (.A(_21964_),
    .Z(_21965_));
 BUF_X8 _51150_ (.A(_21965_),
    .Z(_21966_));
 MUX2_X1 _51151_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1960]),
    .B(_21863_),
    .S(_21966_),
    .Z(_01888_));
 MUX2_X1 _51152_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1961]),
    .B(_21867_),
    .S(_21966_),
    .Z(_01889_));
 BUF_X16 _51153_ (.A(_21294_),
    .Z(_21967_));
 MUX2_X1 _51154_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1962]),
    .B(_21967_),
    .S(_21966_),
    .Z(_01890_));
 MUX2_X1 _51155_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1963]),
    .B(_21868_),
    .S(_21966_),
    .Z(_01891_));
 BUF_X16 _51156_ (.A(_21297_),
    .Z(_21968_));
 MUX2_X1 _51157_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1964]),
    .B(_21968_),
    .S(_21966_),
    .Z(_01892_));
 MUX2_X1 _51158_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1965]),
    .B(_21885_),
    .S(_21966_),
    .Z(_01893_));
 MUX2_X1 _51159_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1966]),
    .B(_21745_),
    .S(_21966_),
    .Z(_01894_));
 BUF_X16 _51160_ (.A(_21303_),
    .Z(_21969_));
 MUX2_X1 _51161_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1967]),
    .B(_21969_),
    .S(_21966_),
    .Z(_01895_));
 MUX2_X1 _51162_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1968]),
    .B(_21689_),
    .S(_21966_),
    .Z(_01896_));
 BUF_X8 _51163_ (.A(_21964_),
    .Z(_21970_));
 MUX2_X1 _51164_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1969]),
    .B(_21749_),
    .S(_21970_),
    .Z(_01897_));
 BUF_X16 _51165_ (.A(_21309_),
    .Z(_21971_));
 MUX2_X1 _51166_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1970]),
    .B(_21971_),
    .S(_21970_),
    .Z(_01899_));
 MUX2_X1 _51167_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1971]),
    .B(_21750_),
    .S(_21970_),
    .Z(_01900_));
 MUX2_X1 _51168_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1972]),
    .B(_21833_),
    .S(_21970_),
    .Z(_01901_));
 MUX2_X1 _51169_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1973]),
    .B(_21852_),
    .S(_21970_),
    .Z(_01902_));
 MUX2_X1 _51170_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1974]),
    .B(_21804_),
    .S(_21970_),
    .Z(_01903_));
 MUX2_X1 _51171_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1975]),
    .B(_21773_),
    .S(_21970_),
    .Z(_01904_));
 MUX2_X1 _51172_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1976]),
    .B(_21805_),
    .S(_21970_),
    .Z(_01905_));
 MUX2_X1 _51173_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1977]),
    .B(_21948_),
    .S(_21970_),
    .Z(_01906_));
 MUX2_X1 _51174_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1978]),
    .B(_21807_),
    .S(_21970_),
    .Z(_01907_));
 BUF_X8 _51175_ (.A(_21964_),
    .Z(_21972_));
 MUX2_X1 _51176_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1979]),
    .B(_21777_),
    .S(_21972_),
    .Z(_01908_));
 MUX2_X1 _51177_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1980]),
    .B(_21778_),
    .S(_21972_),
    .Z(_01910_));
 MUX2_X1 _51178_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1981]),
    .B(_21779_),
    .S(_21972_),
    .Z(_01911_));
 MUX2_X1 _51179_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1982]),
    .B(_21780_),
    .S(_21972_),
    .Z(_01912_));
 BUF_X16 _51180_ (.A(_08588_),
    .Z(_21973_));
 MUX2_X1 _51181_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1983]),
    .B(_21973_),
    .S(_21972_),
    .Z(_01913_));
 MUX2_X1 _51182_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1984]),
    .B(_21837_),
    .S(_21972_),
    .Z(_01914_));
 NAND4_X1 _51183_ (.A1(_21786_),
    .A2(_21757_),
    .A3(_21945_),
    .A4(_10942_),
    .ZN(_21974_));
 INV_X1 _51184_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1985]),
    .ZN(_21975_));
 OAI21_X1 _51185_ (.A(_21974_),
    .B1(_21966_),
    .B2(_21975_),
    .ZN(_01915_));
 MUX2_X1 _51186_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1986]),
    .B(_21783_),
    .S(_21972_),
    .Z(_01916_));
 MUX2_X1 _51187_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1987]),
    .B(_21952_),
    .S(_21972_),
    .Z(_01917_));
 MUX2_X1 _51188_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1988]),
    .B(_21555_),
    .S(_21972_),
    .Z(_01918_));
 MUX2_X1 _51189_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1989]),
    .B(_21860_),
    .S(_21972_),
    .Z(_01919_));
 BUF_X16 _51190_ (.A(_21964_),
    .Z(_21976_));
 MUX2_X1 _51191_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1990]),
    .B(_21955_),
    .S(_21976_),
    .Z(_01921_));
 MUX2_X1 _51192_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1991]),
    .B(_21862_),
    .S(_21976_),
    .Z(_01922_));
 MUX2_X1 _51193_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1992]),
    .B(_21792_),
    .S(_21976_),
    .Z(_01923_));
 MUX2_X1 _51194_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1993]),
    .B(_21793_),
    .S(_21976_),
    .Z(_01924_));
 MUX2_X1 _51195_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1994]),
    .B(_21879_),
    .S(_21976_),
    .Z(_01925_));
 MUX2_X1 _51196_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1995]),
    .B(_21794_),
    .S(_21976_),
    .Z(_01926_));
 MUX2_X1 _51197_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1996]),
    .B(_21795_),
    .S(_21976_),
    .Z(_01927_));
 MUX2_X1 _51198_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1997]),
    .B(_21843_),
    .S(_21976_),
    .Z(_01928_));
 MUX2_X1 _51199_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1998]),
    .B(_21930_),
    .S(_21976_),
    .Z(_01929_));
 MUX2_X1 _51200_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1999]),
    .B(_21762_),
    .S(_21976_),
    .Z(_01930_));
 MUX2_X1 _51201_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2000]),
    .B(_21932_),
    .S(_21965_),
    .Z(_01934_));
 MUX2_X1 _51202_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2001]),
    .B(_21766_),
    .S(_21965_),
    .Z(_01935_));
 MUX2_X1 _51203_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2002]),
    .B(_21737_),
    .S(_21965_),
    .Z(_01936_));
 MUX2_X1 _51204_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2003]),
    .B(_21815_),
    .S(_21965_),
    .Z(_01937_));
 MUX2_X1 _51205_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2004]),
    .B(_21958_),
    .S(_21965_),
    .Z(_01938_));
 MUX2_X1 _51206_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2005]),
    .B(_21898_),
    .S(_21965_),
    .Z(_01939_));
 MUX2_X1 _51207_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2006]),
    .B(_21933_),
    .S(_21965_),
    .Z(_01940_));
 MUX2_X1 _51208_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2007]),
    .B(_21899_),
    .S(_21965_),
    .Z(_01941_));
 BUF_X16 _51209_ (.A(_21377_),
    .Z(_21977_));
 MUX2_X1 _51210_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2008]),
    .B(_21977_),
    .S(_21965_),
    .Z(_01942_));
 BUF_X8 _51211_ (.A(_10983_),
    .Z(_21978_));
 AND2_X4 _51212_ (.A1(_21978_),
    .A2(_21679_),
    .ZN(_21979_));
 BUF_X16 _51213_ (.A(_21979_),
    .Z(_21980_));
 BUF_X8 _51214_ (.A(_21980_),
    .Z(_21981_));
 MUX2_X1 _51215_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1911]),
    .B(_21863_),
    .S(_21981_),
    .Z(_01834_));
 MUX2_X1 _51216_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1912]),
    .B(_21867_),
    .S(_21981_),
    .Z(_01835_));
 MUX2_X1 _51217_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1913]),
    .B(_21967_),
    .S(_21981_),
    .Z(_01836_));
 MUX2_X1 _51218_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1914]),
    .B(_21868_),
    .S(_21981_),
    .Z(_01837_));
 BUF_X16 _51219_ (.A(_21979_),
    .Z(_21982_));
 MUX2_X1 _51220_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1915]),
    .B(_21968_),
    .S(_21982_),
    .Z(_01838_));
 MUX2_X1 _51221_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1916]),
    .B(_21885_),
    .S(_21982_),
    .Z(_01839_));
 BUF_X8 _51222_ (.A(_10990_),
    .Z(_21983_));
 NAND4_X1 _51223_ (.A1(_21799_),
    .A2(_21301_),
    .A3(_21945_),
    .A4(_21983_),
    .ZN(_21984_));
 INV_X1 _51224_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1917]),
    .ZN(_21985_));
 OAI21_X1 _51225_ (.A(_21984_),
    .B1(_21981_),
    .B2(_21985_),
    .ZN(_01840_));
 NAND4_X4 _51226_ (.A1(_21799_),
    .A2(_21303_),
    .A3(_21945_),
    .A4(_21983_),
    .ZN(_21986_));
 INV_X1 _51227_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1918]),
    .ZN(_21987_));
 OAI21_X1 _51228_ (.A(_21986_),
    .B1(_21981_),
    .B2(_21987_),
    .ZN(_01841_));
 MUX2_X1 _51229_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1919]),
    .B(_21689_),
    .S(_21982_),
    .Z(_01842_));
 BUF_X8 _51230_ (.A(_21307_),
    .Z(_21988_));
 MUX2_X1 _51231_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1920]),
    .B(_21988_),
    .S(_21982_),
    .Z(_01844_));
 MUX2_X1 _51232_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1921]),
    .B(_21971_),
    .S(_21982_),
    .Z(_01845_));
 MUX2_X1 _51233_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1922]),
    .B(_21750_),
    .S(_21982_),
    .Z(_01846_));
 MUX2_X1 _51234_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1923]),
    .B(_21833_),
    .S(_21982_),
    .Z(_01847_));
 MUX2_X1 _51235_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1924]),
    .B(_21852_),
    .S(_21982_),
    .Z(_01848_));
 MUX2_X1 _51236_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1925]),
    .B(_21804_),
    .S(_21982_),
    .Z(_01849_));
 MUX2_X1 _51237_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1926]),
    .B(_21773_),
    .S(_21982_),
    .Z(_01850_));
 BUF_X8 _51238_ (.A(_21979_),
    .Z(_21989_));
 MUX2_X1 _51239_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1927]),
    .B(_21805_),
    .S(_21989_),
    .Z(_01851_));
 MUX2_X1 _51240_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1928]),
    .B(_21948_),
    .S(_21989_),
    .Z(_01852_));
 MUX2_X1 _51241_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1929]),
    .B(_21807_),
    .S(_21989_),
    .Z(_01853_));
 MUX2_X1 _51242_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1930]),
    .B(_21777_),
    .S(_21989_),
    .Z(_01855_));
 MUX2_X1 _51243_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1931]),
    .B(_21778_),
    .S(_21989_),
    .Z(_01856_));
 MUX2_X1 _51244_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1932]),
    .B(_21779_),
    .S(_21989_),
    .Z(_01857_));
 MUX2_X1 _51245_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1933]),
    .B(_21780_),
    .S(_21989_),
    .Z(_01858_));
 MUX2_X1 _51246_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1934]),
    .B(_21973_),
    .S(_21989_),
    .Z(_01859_));
 MUX2_X1 _51247_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1935]),
    .B(_21837_),
    .S(_21989_),
    .Z(_01860_));
 MUX2_X1 _51248_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1936]),
    .B(_21919_),
    .S(_21989_),
    .Z(_01861_));
 BUF_X8 _51249_ (.A(_21979_),
    .Z(_21990_));
 MUX2_X1 _51250_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1937]),
    .B(_21783_),
    .S(_21990_),
    .Z(_01862_));
 MUX2_X1 _51251_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1938]),
    .B(_21952_),
    .S(_21990_),
    .Z(_01863_));
 BUF_X8 _51252_ (.A(_08604_),
    .Z(_21991_));
 MUX2_X1 _51253_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1939]),
    .B(_21991_),
    .S(_21990_),
    .Z(_01864_));
 MUX2_X1 _51254_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1940]),
    .B(_21860_),
    .S(_21990_),
    .Z(_01866_));
 MUX2_X1 _51255_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1941]),
    .B(_21955_),
    .S(_21990_),
    .Z(_01867_));
 MUX2_X1 _51256_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1942]),
    .B(_21862_),
    .S(_21990_),
    .Z(_01868_));
 MUX2_X1 _51257_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1943]),
    .B(_21792_),
    .S(_21990_),
    .Z(_01869_));
 MUX2_X1 _51258_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1944]),
    .B(_21793_),
    .S(_21990_),
    .Z(_01870_));
 MUX2_X1 _51259_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1945]),
    .B(_21879_),
    .S(_21990_),
    .Z(_01871_));
 MUX2_X1 _51260_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1946]),
    .B(_21794_),
    .S(_21990_),
    .Z(_01872_));
 MUX2_X1 _51261_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1947]),
    .B(_21795_),
    .S(_21980_),
    .Z(_01873_));
 NAND4_X1 _51262_ (.A1(_21799_),
    .A2(_21330_),
    .A3(_21945_),
    .A4(_21983_),
    .ZN(_21992_));
 INV_X1 _51263_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1948]),
    .ZN(_21993_));
 OAI21_X1 _51264_ (.A(_21992_),
    .B1(_21981_),
    .B2(_21993_),
    .ZN(_01874_));
 BUF_X4 _51265_ (.A(_10990_),
    .Z(_21994_));
 NAND4_X1 _51266_ (.A1(_21799_),
    .A2(_21591_),
    .A3(_21945_),
    .A4(_21994_),
    .ZN(_21995_));
 INV_X2 _51267_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1949]),
    .ZN(_21996_));
 OAI21_X1 _51268_ (.A(_21995_),
    .B1(_21981_),
    .B2(_21996_),
    .ZN(_01875_));
 NAND4_X4 _51269_ (.A1(_21799_),
    .A2(_21934_),
    .A3(_10991_),
    .A4(_21339_),
    .ZN(_21997_));
 INV_X1 _51270_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1950]),
    .ZN(_21998_));
 OAI21_X1 _51271_ (.A(_21997_),
    .B1(_21981_),
    .B2(_21998_),
    .ZN(_01877_));
 MUX2_X1 _51272_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1951]),
    .B(_21932_),
    .S(_21980_),
    .Z(_01878_));
 BUF_X8 _51273_ (.A(_21347_),
    .Z(_21999_));
 MUX2_X1 _51274_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1952]),
    .B(_21999_),
    .S(_21980_),
    .Z(_01879_));
 BUF_X16 _51275_ (.A(_21351_),
    .Z(_22000_));
 MUX2_X1 _51276_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1953]),
    .B(_22000_),
    .S(_21980_),
    .Z(_01880_));
 MUX2_X1 _51277_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1954]),
    .B(_21815_),
    .S(_21980_),
    .Z(_01881_));
 MUX2_X1 _51278_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1955]),
    .B(_21958_),
    .S(_21980_),
    .Z(_01882_));
 MUX2_X1 _51279_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1956]),
    .B(_21898_),
    .S(_21980_),
    .Z(_01883_));
 MUX2_X1 _51280_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1957]),
    .B(_21933_),
    .S(_21980_),
    .Z(_01884_));
 NAND4_X1 _51281_ (.A1(_21799_),
    .A2(_21934_),
    .A3(_10991_),
    .A4(_21373_),
    .ZN(_22001_));
 INV_X1 _51282_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1958]),
    .ZN(_22002_));
 OAI21_X1 _51283_ (.A(_22001_),
    .B1(_21981_),
    .B2(_22002_),
    .ZN(_01885_));
 MUX2_X1 _51284_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1959]),
    .B(_21977_),
    .S(_21980_),
    .Z(_01886_));
 BUF_X16 _51285_ (.A(_10993_),
    .Z(_22003_));
 AND2_X4 _51286_ (.A1(_22003_),
    .A2(_21290_),
    .ZN(_22004_));
 BUF_X8 _51287_ (.A(_22004_),
    .Z(_22005_));
 MUX2_X1 _51288_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1862]),
    .B(_21863_),
    .S(_22005_),
    .Z(_01779_));
 MUX2_X1 _51289_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1863]),
    .B(_21867_),
    .S(_22005_),
    .Z(_01780_));
 MUX2_X1 _51290_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1864]),
    .B(_21967_),
    .S(_22005_),
    .Z(_01781_));
 MUX2_X1 _51291_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1865]),
    .B(_21868_),
    .S(_22005_),
    .Z(_01782_));
 MUX2_X1 _51292_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1866]),
    .B(_21968_),
    .S(_22005_),
    .Z(_01783_));
 MUX2_X1 _51293_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1867]),
    .B(_21885_),
    .S(_22005_),
    .Z(_01784_));
 BUF_X4 _51294_ (.A(_10819_),
    .Z(_22006_));
 NAND4_X1 _51295_ (.A1(_22006_),
    .A2(_21301_),
    .A3(_21945_),
    .A4(_21994_),
    .ZN(_22007_));
 BUF_X4 _51296_ (.A(_22005_),
    .Z(_22008_));
 INV_X1 _51297_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1868]),
    .ZN(_22009_));
 OAI21_X1 _51298_ (.A(_22007_),
    .B1(_22008_),
    .B2(_22009_),
    .ZN(_01785_));
 NAND4_X2 _51299_ (.A1(_22006_),
    .A2(_21303_),
    .A3(_21945_),
    .A4(_21994_),
    .ZN(_22010_));
 INV_X1 _51300_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1869]),
    .ZN(_22011_));
 OAI21_X1 _51301_ (.A(_22010_),
    .B1(_22008_),
    .B2(_22011_),
    .ZN(_01786_));
 BUF_X16 _51302_ (.A(_21305_),
    .Z(_22012_));
 MUX2_X1 _51303_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1870]),
    .B(_22012_),
    .S(_22005_),
    .Z(_01788_));
 MUX2_X1 _51304_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1871]),
    .B(_21988_),
    .S(_22005_),
    .Z(_01789_));
 BUF_X4 _51305_ (.A(_21856_),
    .Z(_22013_));
 NAND4_X1 _51306_ (.A1(_22006_),
    .A2(_21446_),
    .A3(_22013_),
    .A4(_21994_),
    .ZN(_22014_));
 INV_X2 _51307_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1872]),
    .ZN(_22015_));
 OAI21_X1 _51308_ (.A(_22014_),
    .B1(_22008_),
    .B2(_22015_),
    .ZN(_01790_));
 BUF_X16 _51309_ (.A(_22004_),
    .Z(_22016_));
 MUX2_X1 _51310_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1873]),
    .B(_21750_),
    .S(_22016_),
    .Z(_01791_));
 MUX2_X1 _51311_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1874]),
    .B(_21833_),
    .S(_22016_),
    .Z(_01792_));
 MUX2_X1 _51312_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1875]),
    .B(_21852_),
    .S(_22016_),
    .Z(_01793_));
 MUX2_X1 _51313_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1876]),
    .B(_21804_),
    .S(_22016_),
    .Z(_01794_));
 MUX2_X1 _51314_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1877]),
    .B(_21773_),
    .S(_22016_),
    .Z(_01795_));
 NAND4_X1 _51315_ (.A1(_22006_),
    .A2(_10572_),
    .A3(_22013_),
    .A4(_21994_),
    .ZN(_22017_));
 INV_X1 _51316_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1878]),
    .ZN(_22018_));
 OAI21_X1 _51317_ (.A(_22017_),
    .B1(_22008_),
    .B2(_22018_),
    .ZN(_01796_));
 MUX2_X1 _51318_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1879]),
    .B(_21948_),
    .S(_22016_),
    .Z(_01797_));
 MUX2_X1 _51319_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1880]),
    .B(_21807_),
    .S(_22016_),
    .Z(_01799_));
 BUF_X8 _51320_ (.A(_08575_),
    .Z(_22019_));
 MUX2_X1 _51321_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1881]),
    .B(_22019_),
    .S(_22016_),
    .Z(_01800_));
 NAND4_X1 _51322_ (.A1(_22006_),
    .A2(_10614_),
    .A3(_22013_),
    .A4(_21994_),
    .ZN(_22020_));
 INV_X1 _51323_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1882]),
    .ZN(_22021_));
 OAI21_X1 _51324_ (.A(_22020_),
    .B1(_22008_),
    .B2(_22021_),
    .ZN(_01801_));
 BUF_X8 _51325_ (.A(_08581_),
    .Z(_22022_));
 MUX2_X1 _51326_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1883]),
    .B(_22022_),
    .S(_22016_),
    .Z(_01802_));
 BUF_X8 _51327_ (.A(_08584_),
    .Z(_22023_));
 MUX2_X1 _51328_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1884]),
    .B(_22023_),
    .S(_22016_),
    .Z(_01803_));
 BUF_X8 _51329_ (.A(_22004_),
    .Z(_22024_));
 MUX2_X1 _51330_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1885]),
    .B(_21973_),
    .S(_22024_),
    .Z(_01804_));
 BUF_X32 _51331_ (.A(_08591_),
    .Z(_22025_));
 NAND4_X1 _51332_ (.A1(_22006_),
    .A2(_22025_),
    .A3(_22013_),
    .A4(_21994_),
    .ZN(_22026_));
 INV_X1 _51333_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1886]),
    .ZN(_22027_));
 OAI21_X1 _51334_ (.A(_22026_),
    .B1(_22008_),
    .B2(_22027_),
    .ZN(_01805_));
 MUX2_X1 _51335_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1887]),
    .B(_21919_),
    .S(_22024_),
    .Z(_01806_));
 BUF_X16 _51336_ (.A(_08597_),
    .Z(_22028_));
 MUX2_X1 _51337_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1888]),
    .B(_22028_),
    .S(_22024_),
    .Z(_01807_));
 NAND4_X1 _51338_ (.A1(_22006_),
    .A2(_21520_),
    .A3(_22013_),
    .A4(_21994_),
    .ZN(_22029_));
 INV_X1 _51339_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1889]),
    .ZN(_22030_));
 OAI21_X1 _51340_ (.A(_22029_),
    .B1(_22008_),
    .B2(_22030_),
    .ZN(_01808_));
 MUX2_X1 _51341_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1890]),
    .B(_21991_),
    .S(_22024_),
    .Z(_01810_));
 MUX2_X1 _51342_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1891]),
    .B(_21860_),
    .S(_22024_),
    .Z(_01811_));
 NAND4_X2 _51343_ (.A1(_22006_),
    .A2(_21558_),
    .A3(_22013_),
    .A4(_21994_),
    .ZN(_22031_));
 INV_X1 _51344_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1892]),
    .ZN(_22032_));
 OAI21_X1 _51345_ (.A(_22031_),
    .B1(_22008_),
    .B2(_22032_),
    .ZN(_01812_));
 MUX2_X1 _51346_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1893]),
    .B(_21862_),
    .S(_22024_),
    .Z(_01813_));
 BUF_X8 _51347_ (.A(_08617_),
    .Z(_22033_));
 MUX2_X1 _51348_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1894]),
    .B(_22033_),
    .S(_22024_),
    .Z(_01814_));
 BUF_X8 _51349_ (.A(_08620_),
    .Z(_22034_));
 MUX2_X1 _51350_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1895]),
    .B(_22034_),
    .S(_22024_),
    .Z(_01815_));
 MUX2_X1 _51351_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1896]),
    .B(_21879_),
    .S(_22024_),
    .Z(_01816_));
 BUF_X16 _51352_ (.A(_08626_),
    .Z(_22035_));
 MUX2_X1 _51353_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1897]),
    .B(_22035_),
    .S(_22024_),
    .Z(_01817_));
 BUF_X16 _51354_ (.A(_22004_),
    .Z(_22036_));
 MUX2_X1 _51355_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1898]),
    .B(_21795_),
    .S(_22036_),
    .Z(_01818_));
 NAND4_X1 _51356_ (.A1(_22006_),
    .A2(_21330_),
    .A3(_22013_),
    .A4(_21994_),
    .ZN(_22037_));
 INV_X1 _51357_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1899]),
    .ZN(_22038_));
 OAI21_X1 _51358_ (.A(_22037_),
    .B1(_22008_),
    .B2(_22038_),
    .ZN(_01819_));
 MUX2_X1 _51359_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1900]),
    .B(_21930_),
    .S(_22036_),
    .Z(_01822_));
 NAND4_X4 _51360_ (.A1(_22006_),
    .A2(_21934_),
    .A3(_21983_),
    .A4(_21339_),
    .ZN(_22039_));
 INV_X1 _51361_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1901]),
    .ZN(_22040_));
 OAI21_X1 _51362_ (.A(_22039_),
    .B1(_22008_),
    .B2(_22040_),
    .ZN(_01823_));
 MUX2_X1 _51363_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1902]),
    .B(_21932_),
    .S(_22036_),
    .Z(_01824_));
 MUX2_X1 _51364_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1903]),
    .B(_21999_),
    .S(_22036_),
    .Z(_01825_));
 BUF_X16 _51365_ (.A(_10819_),
    .Z(_22041_));
 NAND4_X2 _51366_ (.A1(_22041_),
    .A2(_21934_),
    .A3(_21983_),
    .A4(_21351_),
    .ZN(_22042_));
 INV_X1 _51367_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1904]),
    .ZN(_22043_));
 OAI21_X1 _51368_ (.A(_22042_),
    .B1(_22005_),
    .B2(_22043_),
    .ZN(_01826_));
 MUX2_X1 _51369_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1905]),
    .B(_21815_),
    .S(_22036_),
    .Z(_01827_));
 MUX2_X1 _51370_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1906]),
    .B(_21958_),
    .S(_22036_),
    .Z(_01828_));
 MUX2_X1 _51371_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1907]),
    .B(_21898_),
    .S(_22036_),
    .Z(_01829_));
 MUX2_X1 _51372_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1908]),
    .B(_21933_),
    .S(_22036_),
    .Z(_01830_));
 MUX2_X1 _51373_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1909]),
    .B(_21899_),
    .S(_22036_),
    .Z(_01831_));
 MUX2_X1 _51374_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1910]),
    .B(_21977_),
    .S(_22036_),
    .Z(_01833_));
 BUF_X16 _51375_ (.A(_10997_),
    .Z(_22044_));
 AND2_X4 _51376_ (.A1(_22044_),
    .A2(_21432_),
    .ZN(_22045_));
 BUF_X16 _51377_ (.A(_22045_),
    .Z(_22046_));
 BUF_X8 _51378_ (.A(_22046_),
    .Z(_22047_));
 MUX2_X1 _51379_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1813]),
    .B(_21863_),
    .S(_22047_),
    .Z(_01725_));
 MUX2_X1 _51380_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1814]),
    .B(_21867_),
    .S(_22047_),
    .Z(_01726_));
 MUX2_X1 _51381_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1815]),
    .B(_21967_),
    .S(_22047_),
    .Z(_01727_));
 MUX2_X1 _51382_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1816]),
    .B(_21868_),
    .S(_22047_),
    .Z(_01728_));
 MUX2_X1 _51383_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1817]),
    .B(_21968_),
    .S(_22047_),
    .Z(_01729_));
 MUX2_X1 _51384_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1818]),
    .B(_21885_),
    .S(_22047_),
    .Z(_01730_));
 MUX2_X1 _51385_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1819]),
    .B(_21745_),
    .S(_22047_),
    .Z(_01731_));
 BUF_X16 _51386_ (.A(_22045_),
    .Z(_22048_));
 MUX2_X1 _51387_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1820]),
    .B(_21969_),
    .S(_22048_),
    .Z(_01733_));
 MUX2_X1 _51388_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1821]),
    .B(_22012_),
    .S(_22048_),
    .Z(_01734_));
 MUX2_X1 _51389_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1822]),
    .B(_21988_),
    .S(_22048_),
    .Z(_01735_));
 MUX2_X1 _51390_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1823]),
    .B(_21971_),
    .S(_22048_),
    .Z(_01736_));
 BUF_X16 _51391_ (.A(_21311_),
    .Z(_22049_));
 MUX2_X1 _51392_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1824]),
    .B(_22049_),
    .S(_22048_),
    .Z(_01737_));
 MUX2_X1 _51393_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1825]),
    .B(_21833_),
    .S(_22048_),
    .Z(_01738_));
 MUX2_X1 _51394_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1826]),
    .B(_21852_),
    .S(_22048_),
    .Z(_01739_));
 BUF_X8 _51395_ (.A(_08558_),
    .Z(_22050_));
 MUX2_X1 _51396_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1827]),
    .B(_22050_),
    .S(_22048_),
    .Z(_01740_));
 MUX2_X1 _51397_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1828]),
    .B(_21773_),
    .S(_22048_),
    .Z(_01741_));
 MUX2_X1 _51398_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1829]),
    .B(_21805_),
    .S(_22048_),
    .Z(_01742_));
 BUF_X16 _51399_ (.A(_22045_),
    .Z(_22051_));
 MUX2_X1 _51400_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1830]),
    .B(_21948_),
    .S(_22051_),
    .Z(_01744_));
 BUF_X8 _51401_ (.A(_08571_),
    .Z(_22052_));
 MUX2_X1 _51402_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1831]),
    .B(_22052_),
    .S(_22051_),
    .Z(_01745_));
 MUX2_X1 _51403_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1832]),
    .B(_22019_),
    .S(_22051_),
    .Z(_01746_));
 BUF_X4 _51404_ (.A(_10990_),
    .Z(_22053_));
 NAND4_X1 _51405_ (.A1(_21640_),
    .A2(_10614_),
    .A3(_22013_),
    .A4(_22053_),
    .ZN(_22054_));
 INV_X1 _51406_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1833]),
    .ZN(_22055_));
 OAI21_X1 _51407_ (.A(_22054_),
    .B1(_22047_),
    .B2(_22055_),
    .ZN(_01747_));
 MUX2_X1 _51408_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1834]),
    .B(_22022_),
    .S(_22051_),
    .Z(_01748_));
 MUX2_X1 _51409_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1835]),
    .B(_22023_),
    .S(_22051_),
    .Z(_01749_));
 MUX2_X1 _51410_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1836]),
    .B(_21973_),
    .S(_22051_),
    .Z(_01750_));
 NAND4_X1 _51411_ (.A1(_21640_),
    .A2(_22025_),
    .A3(_22013_),
    .A4(_22053_),
    .ZN(_22056_));
 INV_X1 _51412_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1837]),
    .ZN(_22057_));
 OAI21_X1 _51413_ (.A(_22056_),
    .B1(_22047_),
    .B2(_22057_),
    .ZN(_01751_));
 MUX2_X1 _51414_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1838]),
    .B(_21919_),
    .S(_22051_),
    .Z(_01752_));
 MUX2_X1 _51415_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1839]),
    .B(_22028_),
    .S(_22051_),
    .Z(_01753_));
 MUX2_X1 _51416_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1840]),
    .B(_21952_),
    .S(_22051_),
    .Z(_01755_));
 MUX2_X1 _51417_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1841]),
    .B(_21991_),
    .S(_22051_),
    .Z(_01756_));
 BUF_X16 _51418_ (.A(_22045_),
    .Z(_22058_));
 MUX2_X1 _51419_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1842]),
    .B(_21860_),
    .S(_22058_),
    .Z(_01757_));
 NAND4_X2 _51420_ (.A1(_21640_),
    .A2(_21558_),
    .A3(_22013_),
    .A4(_22053_),
    .ZN(_22059_));
 INV_X1 _51421_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1843]),
    .ZN(_22060_));
 OAI21_X1 _51422_ (.A(_22059_),
    .B1(_22047_),
    .B2(_22060_),
    .ZN(_01758_));
 MUX2_X1 _51423_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1844]),
    .B(_21862_),
    .S(_22058_),
    .Z(_01759_));
 MUX2_X1 _51424_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1845]),
    .B(_22033_),
    .S(_22058_),
    .Z(_01760_));
 MUX2_X1 _51425_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1846]),
    .B(_22034_),
    .S(_22058_),
    .Z(_01761_));
 MUX2_X1 _51426_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1847]),
    .B(_21879_),
    .S(_22058_),
    .Z(_01762_));
 MUX2_X1 _51427_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1848]),
    .B(_22035_),
    .S(_22058_),
    .Z(_01763_));
 MUX2_X1 _51428_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1849]),
    .B(_21795_),
    .S(_22058_),
    .Z(_01764_));
 MUX2_X1 _51429_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1850]),
    .B(_21843_),
    .S(_22058_),
    .Z(_01766_));
 MUX2_X1 _51430_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1851]),
    .B(_21930_),
    .S(_22058_),
    .Z(_01767_));
 MUX2_X1 _51431_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1852]),
    .B(_21762_),
    .S(_22058_),
    .Z(_01768_));
 MUX2_X1 _51432_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1853]),
    .B(_21932_),
    .S(_22046_),
    .Z(_01769_));
 MUX2_X1 _51433_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1854]),
    .B(_21999_),
    .S(_22046_),
    .Z(_01770_));
 MUX2_X1 _51434_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1855]),
    .B(_22000_),
    .S(_22046_),
    .Z(_01771_));
 BUF_X16 _51435_ (.A(_21355_),
    .Z(_22061_));
 MUX2_X1 _51436_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1856]),
    .B(_22061_),
    .S(_22046_),
    .Z(_01772_));
 MUX2_X1 _51437_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1857]),
    .B(_21958_),
    .S(_22046_),
    .Z(_01773_));
 MUX2_X1 _51438_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1858]),
    .B(_21898_),
    .S(_22046_),
    .Z(_01774_));
 MUX2_X1 _51439_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1859]),
    .B(_21933_),
    .S(_22046_),
    .Z(_01775_));
 MUX2_X1 _51440_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1860]),
    .B(_21899_),
    .S(_22046_),
    .Z(_01777_));
 MUX2_X1 _51441_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1861]),
    .B(_21977_),
    .S(_22046_),
    .Z(_01778_));
 AND2_X4 _51442_ (.A1(_11002_),
    .A2(_21432_),
    .ZN(_22062_));
 BUF_X16 _51443_ (.A(_22062_),
    .Z(_22063_));
 BUF_X8 _51444_ (.A(_22063_),
    .Z(_22064_));
 MUX2_X1 _51445_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1764]),
    .B(_21863_),
    .S(_22064_),
    .Z(_01670_));
 MUX2_X1 _51446_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1765]),
    .B(_21867_),
    .S(_22064_),
    .Z(_01671_));
 MUX2_X1 _51447_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1766]),
    .B(_21967_),
    .S(_22064_),
    .Z(_01672_));
 MUX2_X1 _51448_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1767]),
    .B(_21868_),
    .S(_22064_),
    .Z(_01673_));
 MUX2_X1 _51449_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1768]),
    .B(_21968_),
    .S(_22064_),
    .Z(_01674_));
 MUX2_X1 _51450_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1769]),
    .B(_21885_),
    .S(_22064_),
    .Z(_01675_));
 MUX2_X1 _51451_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1770]),
    .B(_21745_),
    .S(_22064_),
    .Z(_01677_));
 BUF_X16 _51452_ (.A(_22062_),
    .Z(_22065_));
 MUX2_X1 _51453_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1771]),
    .B(_21969_),
    .S(_22065_),
    .Z(_01678_));
 MUX2_X1 _51454_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1772]),
    .B(_22012_),
    .S(_22065_),
    .Z(_01679_));
 MUX2_X1 _51455_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1773]),
    .B(_21988_),
    .S(_22065_),
    .Z(_01680_));
 MUX2_X1 _51456_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1774]),
    .B(_21971_),
    .S(_22065_),
    .Z(_01681_));
 MUX2_X1 _51457_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1775]),
    .B(_22049_),
    .S(_22065_),
    .Z(_01682_));
 MUX2_X1 _51458_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1776]),
    .B(_21833_),
    .S(_22065_),
    .Z(_01683_));
 MUX2_X1 _51459_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1777]),
    .B(_21852_),
    .S(_22065_),
    .Z(_01684_));
 MUX2_X1 _51460_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1778]),
    .B(_22050_),
    .S(_22065_),
    .Z(_01685_));
 BUF_X8 _51461_ (.A(_08561_),
    .Z(_22066_));
 MUX2_X1 _51462_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1779]),
    .B(_22066_),
    .S(_22065_),
    .Z(_01686_));
 BUF_X4 _51463_ (.A(_21856_),
    .Z(_22067_));
 NAND4_X1 _51464_ (.A1(_21672_),
    .A2(_10572_),
    .A3(_22067_),
    .A4(_22053_),
    .ZN(_22068_));
 INV_X1 _51465_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1780]),
    .ZN(_22069_));
 OAI21_X1 _51466_ (.A(_22068_),
    .B1(_22064_),
    .B2(_22069_),
    .ZN(_01688_));
 NAND4_X1 _51467_ (.A1(_21672_),
    .A2(_10599_),
    .A3(_22067_),
    .A4(_22053_),
    .ZN(_22070_));
 INV_X1 _51468_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1781]),
    .ZN(_22071_));
 OAI21_X1 _51469_ (.A(_22070_),
    .B1(_22064_),
    .B2(_22071_),
    .ZN(_01689_));
 MUX2_X1 _51470_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1782]),
    .B(_22052_),
    .S(_22065_),
    .Z(_01690_));
 BUF_X8 _51471_ (.A(_22062_),
    .Z(_22072_));
 MUX2_X1 _51472_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1783]),
    .B(_22019_),
    .S(_22072_),
    .Z(_01691_));
 MUX2_X1 _51473_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1784]),
    .B(_21778_),
    .S(_22072_),
    .Z(_01692_));
 MUX2_X1 _51474_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1785]),
    .B(_22022_),
    .S(_22072_),
    .Z(_01693_));
 MUX2_X1 _51475_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1786]),
    .B(_22023_),
    .S(_22072_),
    .Z(_01694_));
 MUX2_X1 _51476_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1787]),
    .B(_21973_),
    .S(_22072_),
    .Z(_01695_));
 MUX2_X1 _51477_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1788]),
    .B(_21837_),
    .S(_22072_),
    .Z(_01696_));
 MUX2_X1 _51478_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1789]),
    .B(_21919_),
    .S(_22072_),
    .Z(_01697_));
 MUX2_X1 _51479_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1790]),
    .B(_22028_),
    .S(_22072_),
    .Z(_01699_));
 MUX2_X1 _51480_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1791]),
    .B(_21952_),
    .S(_22072_),
    .Z(_01700_));
 MUX2_X1 _51481_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1792]),
    .B(_21991_),
    .S(_22072_),
    .Z(_01701_));
 BUF_X8 _51482_ (.A(_22062_),
    .Z(_22073_));
 MUX2_X1 _51483_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1793]),
    .B(_21860_),
    .S(_22073_),
    .Z(_01702_));
 MUX2_X1 _51484_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1794]),
    .B(_21955_),
    .S(_22073_),
    .Z(_01703_));
 MUX2_X1 _51485_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1795]),
    .B(_21862_),
    .S(_22073_),
    .Z(_01704_));
 MUX2_X1 _51486_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1796]),
    .B(_22033_),
    .S(_22073_),
    .Z(_01705_));
 MUX2_X1 _51487_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1797]),
    .B(_22034_),
    .S(_22073_),
    .Z(_01706_));
 MUX2_X1 _51488_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1798]),
    .B(_21879_),
    .S(_22073_),
    .Z(_01707_));
 MUX2_X1 _51489_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1799]),
    .B(_22035_),
    .S(_22073_),
    .Z(_01708_));
 BUF_X16 _51490_ (.A(_08629_),
    .Z(_22074_));
 MUX2_X1 _51491_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1800]),
    .B(_22074_),
    .S(_22073_),
    .Z(_01711_));
 NAND4_X1 _51492_ (.A1(_21672_),
    .A2(_21330_),
    .A3(_22067_),
    .A4(_22053_),
    .ZN(_22075_));
 INV_X1 _51493_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1801]),
    .ZN(_22076_));
 OAI21_X1 _51494_ (.A(_22075_),
    .B1(_22064_),
    .B2(_22076_),
    .ZN(_01712_));
 MUX2_X1 _51495_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1802]),
    .B(_21930_),
    .S(_22073_),
    .Z(_01713_));
 BUF_X16 _51496_ (.A(_21339_),
    .Z(_22077_));
 MUX2_X1 _51497_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1803]),
    .B(_22077_),
    .S(_22073_),
    .Z(_01714_));
 MUX2_X1 _51498_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1804]),
    .B(_21932_),
    .S(_22063_),
    .Z(_01715_));
 MUX2_X1 _51499_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1805]),
    .B(_21999_),
    .S(_22063_),
    .Z(_01716_));
 MUX2_X1 _51500_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1806]),
    .B(_22000_),
    .S(_22063_),
    .Z(_01717_));
 MUX2_X1 _51501_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1807]),
    .B(_22061_),
    .S(_22063_),
    .Z(_01718_));
 MUX2_X1 _51502_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1808]),
    .B(_21958_),
    .S(_22063_),
    .Z(_01719_));
 MUX2_X1 _51503_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1809]),
    .B(_21898_),
    .S(_22063_),
    .Z(_01720_));
 MUX2_X1 _51504_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1810]),
    .B(_21933_),
    .S(_22063_),
    .Z(_01722_));
 MUX2_X1 _51505_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1811]),
    .B(_21899_),
    .S(_22063_),
    .Z(_01723_));
 MUX2_X1 _51506_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1812]),
    .B(_21977_),
    .S(_22063_),
    .Z(_01724_));
 BUF_X16 _51507_ (.A(_11008_),
    .Z(_22078_));
 AND2_X4 _51508_ (.A1(_22078_),
    .A2(_21441_),
    .ZN(_22079_));
 BUF_X8 _51509_ (.A(_22079_),
    .Z(_22080_));
 BUF_X8 _51510_ (.A(_22080_),
    .Z(_22081_));
 MUX2_X1 _51511_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1715]),
    .B(_21863_),
    .S(_22081_),
    .Z(_01616_));
 MUX2_X1 _51512_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1716]),
    .B(_21867_),
    .S(_22081_),
    .Z(_01617_));
 MUX2_X1 _51513_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1717]),
    .B(_21967_),
    .S(_22081_),
    .Z(_01618_));
 BUF_X8 _51514_ (.A(_22079_),
    .Z(_22082_));
 MUX2_X1 _51515_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1718]),
    .B(_21868_),
    .S(_22082_),
    .Z(_01619_));
 NAND4_X2 _51516_ (.A1(_21890_),
    .A2(_21418_),
    .A3(_22067_),
    .A4(_22053_),
    .ZN(_22083_));
 INV_X1 _51517_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1719]),
    .ZN(_22084_));
 OAI21_X1 _51518_ (.A(_22083_),
    .B1(_22081_),
    .B2(_22084_),
    .ZN(_01620_));
 MUX2_X1 _51519_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1720]),
    .B(_21885_),
    .S(_22082_),
    .Z(_01622_));
 BUF_X16 _51520_ (.A(_21301_),
    .Z(_22085_));
 MUX2_X1 _51521_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1721]),
    .B(_22085_),
    .S(_22082_),
    .Z(_01623_));
 MUX2_X1 _51522_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1722]),
    .B(_21969_),
    .S(_22082_),
    .Z(_01624_));
 MUX2_X1 _51523_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1723]),
    .B(_22012_),
    .S(_22082_),
    .Z(_01625_));
 MUX2_X1 _51524_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1724]),
    .B(_21988_),
    .S(_22082_),
    .Z(_01626_));
 MUX2_X1 _51525_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1725]),
    .B(_21971_),
    .S(_22082_),
    .Z(_01627_));
 NAND4_X1 _51526_ (.A1(_21890_),
    .A2(_21717_),
    .A3(_22067_),
    .A4(_22053_),
    .ZN(_22086_));
 INV_X1 _51527_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1726]),
    .ZN(_22087_));
 OAI21_X1 _51528_ (.A(_22086_),
    .B1(_22081_),
    .B2(_22087_),
    .ZN(_01628_));
 BUF_X8 _51529_ (.A(_08551_),
    .Z(_22088_));
 MUX2_X1 _51530_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1727]),
    .B(_22088_),
    .S(_22082_),
    .Z(_01629_));
 MUX2_X1 _51531_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1728]),
    .B(_21852_),
    .S(_22082_),
    .Z(_01630_));
 MUX2_X1 _51532_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1729]),
    .B(_22050_),
    .S(_22082_),
    .Z(_01631_));
 BUF_X8 _51533_ (.A(_22079_),
    .Z(_22089_));
 MUX2_X1 _51534_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1730]),
    .B(_22066_),
    .S(_22089_),
    .Z(_01633_));
 BUF_X8 _51535_ (.A(_08564_),
    .Z(_22090_));
 MUX2_X1 _51536_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1731]),
    .B(_22090_),
    .S(_22089_),
    .Z(_01634_));
 MUX2_X1 _51537_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1732]),
    .B(_21948_),
    .S(_22089_),
    .Z(_01635_));
 MUX2_X1 _51538_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1733]),
    .B(_22052_),
    .S(_22089_),
    .Z(_01636_));
 MUX2_X1 _51539_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1734]),
    .B(_22019_),
    .S(_22089_),
    .Z(_01637_));
 MUX2_X1 _51540_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1735]),
    .B(_21778_),
    .S(_22089_),
    .Z(_01638_));
 MUX2_X1 _51541_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1736]),
    .B(_22022_),
    .S(_22089_),
    .Z(_01639_));
 MUX2_X1 _51542_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1737]),
    .B(_22023_),
    .S(_22089_),
    .Z(_01640_));
 MUX2_X1 _51543_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1738]),
    .B(_21973_),
    .S(_22089_),
    .Z(_01641_));
 MUX2_X1 _51544_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1739]),
    .B(_21837_),
    .S(_22089_),
    .Z(_01642_));
 NAND4_X2 _51545_ (.A1(_21890_),
    .A2(_21757_),
    .A3(_22067_),
    .A4(_22053_),
    .ZN(_22091_));
 INV_X1 _51546_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1740]),
    .ZN(_22092_));
 OAI21_X1 _51547_ (.A(_22091_),
    .B1(_22081_),
    .B2(_22092_),
    .ZN(_01644_));
 NAND4_X1 _51548_ (.A1(_21890_),
    .A2(_10583_),
    .A3(_22067_),
    .A4(_22053_),
    .ZN(_22093_));
 INV_X1 _51549_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1741]),
    .ZN(_22094_));
 OAI21_X1 _51550_ (.A(_22093_),
    .B1(_22081_),
    .B2(_22094_),
    .ZN(_01645_));
 BUF_X8 _51551_ (.A(_22079_),
    .Z(_22095_));
 MUX2_X1 _51552_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1742]),
    .B(_21952_),
    .S(_22095_),
    .Z(_01646_));
 MUX2_X1 _51553_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1743]),
    .B(_21991_),
    .S(_22095_),
    .Z(_01647_));
 MUX2_X1 _51554_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1744]),
    .B(_21860_),
    .S(_22095_),
    .Z(_01648_));
 BUF_X4 _51555_ (.A(_10990_),
    .Z(_22096_));
 NAND4_X1 _51556_ (.A1(_21890_),
    .A2(_21558_),
    .A3(_22067_),
    .A4(_22096_),
    .ZN(_22097_));
 INV_X1 _51557_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1745]),
    .ZN(_22098_));
 OAI21_X1 _51558_ (.A(_22097_),
    .B1(_22081_),
    .B2(_22098_),
    .ZN(_01649_));
 BUF_X8 _51559_ (.A(_08614_),
    .Z(_22099_));
 MUX2_X1 _51560_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1746]),
    .B(_22099_),
    .S(_22095_),
    .Z(_01650_));
 MUX2_X1 _51561_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1747]),
    .B(_22033_),
    .S(_22095_),
    .Z(_01651_));
 MUX2_X1 _51562_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1748]),
    .B(_22034_),
    .S(_22095_),
    .Z(_01652_));
 MUX2_X1 _51563_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1749]),
    .B(_21879_),
    .S(_22095_),
    .Z(_01653_));
 MUX2_X1 _51564_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1750]),
    .B(_22035_),
    .S(_22095_),
    .Z(_01655_));
 MUX2_X1 _51565_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1751]),
    .B(_22074_),
    .S(_22095_),
    .Z(_01656_));
 MUX2_X1 _51566_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1752]),
    .B(_21843_),
    .S(_22095_),
    .Z(_01657_));
 NAND4_X1 _51567_ (.A1(_21890_),
    .A2(_21591_),
    .A3(_22067_),
    .A4(_22096_),
    .ZN(_22100_));
 INV_X2 _51568_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1753]),
    .ZN(_22101_));
 OAI21_X1 _51569_ (.A(_22100_),
    .B1(_22081_),
    .B2(_22101_),
    .ZN(_01658_));
 MUX2_X1 _51570_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1754]),
    .B(_22077_),
    .S(_22080_),
    .Z(_01659_));
 MUX2_X1 _51571_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1755]),
    .B(_21932_),
    .S(_22080_),
    .Z(_01660_));
 MUX2_X1 _51572_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1756]),
    .B(_21999_),
    .S(_22080_),
    .Z(_01661_));
 MUX2_X1 _51573_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1757]),
    .B(_22000_),
    .S(_22080_),
    .Z(_01662_));
 NAND4_X1 _51574_ (.A1(_21890_),
    .A2(_21934_),
    .A3(_21983_),
    .A4(_21738_),
    .ZN(_22102_));
 INV_X1 _51575_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1758]),
    .ZN(_22103_));
 OAI21_X1 _51576_ (.A(_22102_),
    .B1(_22081_),
    .B2(_22103_),
    .ZN(_01663_));
 MUX2_X1 _51577_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1759]),
    .B(_21958_),
    .S(_22080_),
    .Z(_01664_));
 MUX2_X1 _51578_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1760]),
    .B(_21898_),
    .S(_22080_),
    .Z(_01666_));
 MUX2_X1 _51579_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1761]),
    .B(_21933_),
    .S(_22080_),
    .Z(_01667_));
 MUX2_X1 _51580_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1762]),
    .B(_21899_),
    .S(_22080_),
    .Z(_01668_));
 MUX2_X1 _51581_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1763]),
    .B(_21977_),
    .S(_22080_),
    .Z(_01669_));
 BUF_X16 _51582_ (.A(_21598_),
    .Z(_22104_));
 BUF_X8 _51583_ (.A(_11012_),
    .Z(_22105_));
 AND2_X4 _51584_ (.A1(_22105_),
    .A2(_21441_),
    .ZN(_22106_));
 BUF_X16 _51585_ (.A(_22106_),
    .Z(_22107_));
 BUF_X8 _51586_ (.A(_22107_),
    .Z(_22108_));
 MUX2_X1 _51587_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1666]),
    .B(_22104_),
    .S(_22108_),
    .Z(_01561_));
 BUF_X16 _51588_ (.A(_21605_),
    .Z(_22109_));
 MUX2_X1 _51589_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1667]),
    .B(_22109_),
    .S(_22108_),
    .Z(_01562_));
 MUX2_X1 _51590_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1668]),
    .B(_21967_),
    .S(_22108_),
    .Z(_01563_));
 BUF_X16 _51591_ (.A(_21608_),
    .Z(_22110_));
 BUF_X16 _51592_ (.A(_22106_),
    .Z(_22111_));
 MUX2_X1 _51593_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1669]),
    .B(_22110_),
    .S(_22111_),
    .Z(_01564_));
 BUF_X16 _51594_ (.A(_10859_),
    .Z(_22112_));
 NAND4_X2 _51595_ (.A1(_22112_),
    .A2(_21418_),
    .A3(_22067_),
    .A4(_22096_),
    .ZN(_22113_));
 INV_X1 _51596_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1670]),
    .ZN(_22114_));
 OAI21_X1 _51597_ (.A(_22113_),
    .B1(_22108_),
    .B2(_22114_),
    .ZN(_01566_));
 MUX2_X1 _51598_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1671]),
    .B(_21885_),
    .S(_22111_),
    .Z(_01567_));
 MUX2_X1 _51599_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1672]),
    .B(_22085_),
    .S(_22111_),
    .Z(_01568_));
 MUX2_X1 _51600_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1673]),
    .B(_21969_),
    .S(_22111_),
    .Z(_01569_));
 MUX2_X1 _51601_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1674]),
    .B(_22012_),
    .S(_22111_),
    .Z(_01570_));
 MUX2_X1 _51602_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1675]),
    .B(_21988_),
    .S(_22111_),
    .Z(_01571_));
 BUF_X4 _51603_ (.A(_21856_),
    .Z(_22115_));
 NAND4_X1 _51604_ (.A1(_22112_),
    .A2(_21309_),
    .A3(_22115_),
    .A4(_22096_),
    .ZN(_22116_));
 INV_X4 _51605_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1676]),
    .ZN(_22117_));
 OAI21_X1 _51606_ (.A(_22116_),
    .B1(_22108_),
    .B2(_22117_),
    .ZN(_01572_));
 NAND4_X1 _51607_ (.A1(_22112_),
    .A2(_21717_),
    .A3(_22115_),
    .A4(_22096_),
    .ZN(_22118_));
 INV_X1 _51608_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1677]),
    .ZN(_22119_));
 OAI21_X1 _51609_ (.A(_22118_),
    .B1(_22108_),
    .B2(_22119_),
    .ZN(_01573_));
 MUX2_X1 _51610_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1678]),
    .B(_22088_),
    .S(_22111_),
    .Z(_01574_));
 BUF_X16 _51611_ (.A(_08555_),
    .Z(_22120_));
 MUX2_X1 _51612_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1679]),
    .B(_22120_),
    .S(_22111_),
    .Z(_01575_));
 MUX2_X1 _51613_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1680]),
    .B(_22050_),
    .S(_22111_),
    .Z(_01577_));
 MUX2_X1 _51614_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1681]),
    .B(_22066_),
    .S(_22111_),
    .Z(_01578_));
 BUF_X8 _51615_ (.A(_22106_),
    .Z(_22121_));
 MUX2_X1 _51616_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1682]),
    .B(_22090_),
    .S(_22121_),
    .Z(_01579_));
 MUX2_X1 _51617_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1683]),
    .B(_21948_),
    .S(_22121_),
    .Z(_01580_));
 MUX2_X1 _51618_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1684]),
    .B(_22052_),
    .S(_22121_),
    .Z(_01581_));
 MUX2_X1 _51619_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1685]),
    .B(_22019_),
    .S(_22121_),
    .Z(_01582_));
 MUX2_X1 _51620_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1686]),
    .B(_21778_),
    .S(_22121_),
    .Z(_01583_));
 MUX2_X1 _51621_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1687]),
    .B(_22022_),
    .S(_22121_),
    .Z(_01584_));
 MUX2_X1 _51622_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1688]),
    .B(_22023_),
    .S(_22121_),
    .Z(_01585_));
 MUX2_X1 _51623_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1689]),
    .B(_21973_),
    .S(_22121_),
    .Z(_01586_));
 BUF_X8 _51624_ (.A(_08591_),
    .Z(_22122_));
 MUX2_X1 _51625_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1690]),
    .B(_22122_),
    .S(_22121_),
    .Z(_01588_));
 MUX2_X1 _51626_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1691]),
    .B(_21919_),
    .S(_22121_),
    .Z(_01589_));
 NAND4_X1 _51627_ (.A1(_22112_),
    .A2(_10583_),
    .A3(_22115_),
    .A4(_22096_),
    .ZN(_22123_));
 INV_X1 _51628_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1692]),
    .ZN(_22124_));
 OAI21_X1 _51629_ (.A(_22123_),
    .B1(_22108_),
    .B2(_22124_),
    .ZN(_01590_));
 BUF_X8 _51630_ (.A(_22106_),
    .Z(_22125_));
 MUX2_X1 _51631_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1693]),
    .B(_21952_),
    .S(_22125_),
    .Z(_01591_));
 MUX2_X1 _51632_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1694]),
    .B(_21991_),
    .S(_22125_),
    .Z(_01592_));
 MUX2_X1 _51633_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1695]),
    .B(_21860_),
    .S(_22125_),
    .Z(_01593_));
 NAND4_X1 _51634_ (.A1(_22112_),
    .A2(_21558_),
    .A3(_22115_),
    .A4(_22096_),
    .ZN(_22126_));
 INV_X1 _51635_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1696]),
    .ZN(_22127_));
 OAI21_X1 _51636_ (.A(_22126_),
    .B1(_22108_),
    .B2(_22127_),
    .ZN(_01594_));
 MUX2_X1 _51637_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1697]),
    .B(_22099_),
    .S(_22125_),
    .Z(_01595_));
 MUX2_X1 _51638_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1698]),
    .B(_22033_),
    .S(_22125_),
    .Z(_01596_));
 MUX2_X1 _51639_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1699]),
    .B(_22034_),
    .S(_22125_),
    .Z(_01597_));
 MUX2_X1 _51640_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1700]),
    .B(_21879_),
    .S(_22125_),
    .Z(_01600_));
 MUX2_X1 _51641_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1701]),
    .B(_22035_),
    .S(_22125_),
    .Z(_01601_));
 NAND4_X2 _51642_ (.A1(_22112_),
    .A2(_10593_),
    .A3(_22115_),
    .A4(_22096_),
    .ZN(_22128_));
 INV_X1 _51643_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1702]),
    .ZN(_22129_));
 OAI21_X1 _51644_ (.A(_22128_),
    .B1(_22108_),
    .B2(_22129_),
    .ZN(_01602_));
 MUX2_X1 _51645_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1703]),
    .B(_21843_),
    .S(_22125_),
    .Z(_01603_));
 MUX2_X1 _51646_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1704]),
    .B(_21930_),
    .S(_22125_),
    .Z(_01604_));
 MUX2_X1 _51647_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1705]),
    .B(_22077_),
    .S(_22107_),
    .Z(_01605_));
 MUX2_X1 _51648_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1706]),
    .B(_21932_),
    .S(_22107_),
    .Z(_01606_));
 MUX2_X1 _51649_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1707]),
    .B(_21999_),
    .S(_22107_),
    .Z(_01607_));
 MUX2_X1 _51650_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1708]),
    .B(_22000_),
    .S(_22107_),
    .Z(_01608_));
 NAND4_X1 _51651_ (.A1(_22112_),
    .A2(_21934_),
    .A3(_21983_),
    .A4(_21738_),
    .ZN(_22130_));
 INV_X1 _51652_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1709]),
    .ZN(_22131_));
 OAI21_X1 _51653_ (.A(_22130_),
    .B1(_22108_),
    .B2(_22131_),
    .ZN(_01609_));
 MUX2_X1 _51654_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1710]),
    .B(_21958_),
    .S(_22107_),
    .Z(_01611_));
 MUX2_X1 _51655_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1711]),
    .B(_21898_),
    .S(_22107_),
    .Z(_01612_));
 MUX2_X1 _51656_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1712]),
    .B(_21933_),
    .S(_22107_),
    .Z(_01613_));
 MUX2_X1 _51657_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1713]),
    .B(_21899_),
    .S(_22107_),
    .Z(_01614_));
 MUX2_X1 _51658_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1714]),
    .B(_21977_),
    .S(_22107_),
    .Z(_01615_));
 AND2_X4 _51659_ (.A1(_11019_),
    .A2(_21290_),
    .ZN(_22132_));
 BUF_X16 _51660_ (.A(_22132_),
    .Z(_22133_));
 BUF_X8 _51661_ (.A(_22133_),
    .Z(_22134_));
 MUX2_X1 _51662_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1617]),
    .B(_22104_),
    .S(_22134_),
    .Z(_01507_));
 MUX2_X1 _51663_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1618]),
    .B(_22109_),
    .S(_22134_),
    .Z(_01508_));
 BUF_X16 _51664_ (.A(_22132_),
    .Z(_22135_));
 MUX2_X1 _51665_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1619]),
    .B(_21967_),
    .S(_22135_),
    .Z(_01509_));
 MUX2_X1 _51666_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1620]),
    .B(_22110_),
    .S(_22135_),
    .Z(_01511_));
 MUX2_X1 _51667_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1621]),
    .B(_21968_),
    .S(_22135_),
    .Z(_01512_));
 BUF_X8 _51668_ (.A(_21299_),
    .Z(_22136_));
 MUX2_X1 _51669_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1622]),
    .B(_22136_),
    .S(_22135_),
    .Z(_01513_));
 MUX2_X1 _51670_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1623]),
    .B(_22085_),
    .S(_22135_),
    .Z(_01514_));
 MUX2_X1 _51671_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1624]),
    .B(_21969_),
    .S(_22135_),
    .Z(_01515_));
 MUX2_X1 _51672_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1625]),
    .B(_22012_),
    .S(_22135_),
    .Z(_01516_));
 MUX2_X1 _51673_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1626]),
    .B(_21988_),
    .S(_22135_),
    .Z(_01517_));
 MUX2_X1 _51674_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1627]),
    .B(_21971_),
    .S(_22135_),
    .Z(_01518_));
 NAND4_X1 _51675_ (.A1(_21961_),
    .A2(_21717_),
    .A3(_22115_),
    .A4(_22096_),
    .ZN(_22137_));
 INV_X1 _51676_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1628]),
    .ZN(_22138_));
 OAI21_X1 _51677_ (.A(_22137_),
    .B1(_22134_),
    .B2(_22138_),
    .ZN(_01519_));
 MUX2_X1 _51678_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1629]),
    .B(_22088_),
    .S(_22135_),
    .Z(_01520_));
 BUF_X8 _51679_ (.A(_22132_),
    .Z(_22139_));
 MUX2_X1 _51680_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1630]),
    .B(_22120_),
    .S(_22139_),
    .Z(_01522_));
 MUX2_X1 _51681_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1631]),
    .B(_22050_),
    .S(_22139_),
    .Z(_01523_));
 NAND4_X1 _51682_ (.A1(_21961_),
    .A2(_08561_),
    .A3(_22115_),
    .A4(_22096_),
    .ZN(_22140_));
 INV_X1 _51683_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1632]),
    .ZN(_22141_));
 OAI21_X1 _51684_ (.A(_22140_),
    .B1(_22134_),
    .B2(_22141_),
    .ZN(_01524_));
 BUF_X4 _51685_ (.A(_10990_),
    .Z(_22142_));
 NAND4_X1 _51686_ (.A1(_21961_),
    .A2(_10572_),
    .A3(_22115_),
    .A4(_22142_),
    .ZN(_22143_));
 INV_X2 _51687_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1633]),
    .ZN(_22144_));
 OAI21_X1 _51688_ (.A(_22143_),
    .B1(_22134_),
    .B2(_22144_),
    .ZN(_01525_));
 MUX2_X1 _51689_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1634]),
    .B(_21948_),
    .S(_22139_),
    .Z(_01526_));
 MUX2_X1 _51690_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1635]),
    .B(_22052_),
    .S(_22139_),
    .Z(_01527_));
 MUX2_X1 _51691_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1636]),
    .B(_22019_),
    .S(_22139_),
    .Z(_01528_));
 NAND4_X1 _51692_ (.A1(_21961_),
    .A2(_10614_),
    .A3(_22115_),
    .A4(_22142_),
    .ZN(_22145_));
 INV_X1 _51693_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1637]),
    .ZN(_22146_));
 OAI21_X1 _51694_ (.A(_22145_),
    .B1(_22134_),
    .B2(_22146_),
    .ZN(_01529_));
 MUX2_X1 _51695_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1638]),
    .B(_22022_),
    .S(_22139_),
    .Z(_01530_));
 MUX2_X1 _51696_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1639]),
    .B(_22023_),
    .S(_22139_),
    .Z(_01531_));
 MUX2_X1 _51697_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1640]),
    .B(_21973_),
    .S(_22139_),
    .Z(_01533_));
 MUX2_X1 _51698_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1641]),
    .B(_22122_),
    .S(_22139_),
    .Z(_01534_));
 MUX2_X1 _51699_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1642]),
    .B(_21919_),
    .S(_22139_),
    .Z(_01535_));
 NAND4_X1 _51700_ (.A1(_21961_),
    .A2(_10583_),
    .A3(_22115_),
    .A4(_22142_),
    .ZN(_22147_));
 INV_X1 _51701_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1643]),
    .ZN(_22148_));
 OAI21_X1 _51702_ (.A(_22147_),
    .B1(_22134_),
    .B2(_22148_),
    .ZN(_01536_));
 BUF_X8 _51703_ (.A(_21856_),
    .Z(_22149_));
 NAND4_X1 _51704_ (.A1(_21961_),
    .A2(_21520_),
    .A3(_22149_),
    .A4(_22142_),
    .ZN(_22150_));
 INV_X1 _51705_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1644]),
    .ZN(_22151_));
 OAI21_X1 _51706_ (.A(_22150_),
    .B1(_22134_),
    .B2(_22151_),
    .ZN(_01537_));
 BUF_X8 _51707_ (.A(_22132_),
    .Z(_22152_));
 MUX2_X1 _51708_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1645]),
    .B(_21991_),
    .S(_22152_),
    .Z(_01538_));
 MUX2_X1 _51709_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1646]),
    .B(_21860_),
    .S(_22152_),
    .Z(_01539_));
 MUX2_X1 _51710_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1647]),
    .B(_21955_),
    .S(_22152_),
    .Z(_01540_));
 MUX2_X1 _51711_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1648]),
    .B(_22099_),
    .S(_22152_),
    .Z(_01541_));
 MUX2_X1 _51712_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1649]),
    .B(_22033_),
    .S(_22152_),
    .Z(_01542_));
 MUX2_X1 _51713_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1650]),
    .B(_22034_),
    .S(_22152_),
    .Z(_01544_));
 BUF_X16 _51714_ (.A(_08623_),
    .Z(_22153_));
 MUX2_X1 _51715_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1651]),
    .B(_22153_),
    .S(_22152_),
    .Z(_01545_));
 MUX2_X1 _51716_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1652]),
    .B(_22035_),
    .S(_22152_),
    .Z(_01546_));
 MUX2_X1 _51717_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1653]),
    .B(_22074_),
    .S(_22152_),
    .Z(_01547_));
 MUX2_X1 _51718_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1654]),
    .B(_21843_),
    .S(_22152_),
    .Z(_01548_));
 MUX2_X1 _51719_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1655]),
    .B(_21930_),
    .S(_22133_),
    .Z(_01549_));
 MUX2_X1 _51720_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1656]),
    .B(_22077_),
    .S(_22133_),
    .Z(_01550_));
 MUX2_X1 _51721_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1657]),
    .B(_21932_),
    .S(_22133_),
    .Z(_01551_));
 MUX2_X1 _51722_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1658]),
    .B(_21999_),
    .S(_22133_),
    .Z(_01552_));
 MUX2_X1 _51723_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1659]),
    .B(_22000_),
    .S(_22133_),
    .Z(_01553_));
 BUF_X16 _51724_ (.A(_11015_),
    .Z(_22154_));
 NAND4_X1 _51725_ (.A1(_21961_),
    .A2(_22154_),
    .A3(_21983_),
    .A4(_21738_),
    .ZN(_22155_));
 INV_X1 _51726_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1660]),
    .ZN(_22156_));
 OAI21_X1 _51727_ (.A(_22155_),
    .B1(_22134_),
    .B2(_22156_),
    .ZN(_01555_));
 MUX2_X1 _51728_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1661]),
    .B(_21958_),
    .S(_22133_),
    .Z(_01556_));
 BUF_X8 _51729_ (.A(_21365_),
    .Z(_22157_));
 MUX2_X1 _51730_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1662]),
    .B(_22157_),
    .S(_22133_),
    .Z(_01557_));
 MUX2_X1 _51731_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1663]),
    .B(_21933_),
    .S(_22133_),
    .Z(_01558_));
 NAND4_X1 _51732_ (.A1(_21961_),
    .A2(_22154_),
    .A3(_21983_),
    .A4(_21373_),
    .ZN(_22158_));
 INV_X1 _51733_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1664]),
    .ZN(_22159_));
 OAI21_X1 _51734_ (.A(_22158_),
    .B1(_22134_),
    .B2(_22159_),
    .ZN(_01559_));
 MUX2_X1 _51735_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1665]),
    .B(_21977_),
    .S(_22133_),
    .Z(_01560_));
 AND2_X4 _51736_ (.A1(_11025_),
    .A2(_21441_),
    .ZN(_22160_));
 BUF_X16 _51737_ (.A(_22160_),
    .Z(_22161_));
 BUF_X4 _51738_ (.A(_22161_),
    .Z(_22162_));
 MUX2_X1 _51739_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1568]),
    .B(_22104_),
    .S(_22162_),
    .Z(_01452_));
 MUX2_X1 _51740_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1569]),
    .B(_22109_),
    .S(_22162_),
    .Z(_01453_));
 MUX2_X1 _51741_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1570]),
    .B(_21967_),
    .S(_22162_),
    .Z(_01455_));
 BUF_X16 _51742_ (.A(_22160_),
    .Z(_22163_));
 MUX2_X1 _51743_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1571]),
    .B(_22110_),
    .S(_22163_),
    .Z(_01456_));
 MUX2_X1 _51744_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1572]),
    .B(_21968_),
    .S(_22163_),
    .Z(_01457_));
 MUX2_X1 _51745_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1573]),
    .B(_22136_),
    .S(_22163_),
    .Z(_01458_));
 MUX2_X1 _51746_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1574]),
    .B(_22085_),
    .S(_22163_),
    .Z(_01459_));
 MUX2_X1 _51747_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1575]),
    .B(_21969_),
    .S(_22163_),
    .Z(_01460_));
 MUX2_X1 _51748_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1576]),
    .B(_22012_),
    .S(_22163_),
    .Z(_01461_));
 MUX2_X1 _51749_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1577]),
    .B(_21988_),
    .S(_22163_),
    .Z(_01462_));
 MUX2_X1 _51750_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1578]),
    .B(_21971_),
    .S(_22163_),
    .Z(_01463_));
 NAND4_X1 _51751_ (.A1(_21786_),
    .A2(_21717_),
    .A3(_22149_),
    .A4(_22142_),
    .ZN(_22164_));
 INV_X1 _51752_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1579]),
    .ZN(_22165_));
 OAI21_X1 _51753_ (.A(_22164_),
    .B1(_22162_),
    .B2(_22165_),
    .ZN(_01464_));
 MUX2_X1 _51754_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1580]),
    .B(_22088_),
    .S(_22163_),
    .Z(_01466_));
 MUX2_X1 _51755_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1581]),
    .B(_22120_),
    .S(_22163_),
    .Z(_01467_));
 BUF_X8 _51756_ (.A(_22160_),
    .Z(_22166_));
 MUX2_X1 _51757_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1582]),
    .B(_22050_),
    .S(_22166_),
    .Z(_01468_));
 MUX2_X1 _51758_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1583]),
    .B(_22066_),
    .S(_22166_),
    .Z(_01469_));
 MUX2_X1 _51759_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1584]),
    .B(_22090_),
    .S(_22166_),
    .Z(_01470_));
 MUX2_X1 _51760_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1585]),
    .B(_21948_),
    .S(_22166_),
    .Z(_01471_));
 MUX2_X1 _51761_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1586]),
    .B(_22052_),
    .S(_22166_),
    .Z(_01472_));
 MUX2_X1 _51762_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1587]),
    .B(_22019_),
    .S(_22166_),
    .Z(_01473_));
 BUF_X16 _51763_ (.A(_08578_),
    .Z(_22167_));
 MUX2_X1 _51764_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1588]),
    .B(_22167_),
    .S(_22166_),
    .Z(_01474_));
 MUX2_X1 _51765_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1589]),
    .B(_22022_),
    .S(_22166_),
    .Z(_01475_));
 MUX2_X1 _51766_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1590]),
    .B(_22023_),
    .S(_22166_),
    .Z(_01477_));
 MUX2_X1 _51767_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1591]),
    .B(_21973_),
    .S(_22166_),
    .Z(_01478_));
 BUF_X8 _51768_ (.A(_22160_),
    .Z(_22168_));
 MUX2_X1 _51769_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1592]),
    .B(_22122_),
    .S(_22168_),
    .Z(_01479_));
 NAND4_X1 _51770_ (.A1(_21786_),
    .A2(_21757_),
    .A3(_22149_),
    .A4(_22142_),
    .ZN(_22169_));
 INV_X1 _51771_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1593]),
    .ZN(_22170_));
 OAI21_X1 _51772_ (.A(_22169_),
    .B1(_22162_),
    .B2(_22170_),
    .ZN(_01480_));
 NAND4_X1 _51773_ (.A1(_21786_),
    .A2(_10583_),
    .A3(_22149_),
    .A4(_22142_),
    .ZN(_22171_));
 INV_X1 _51774_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1594]),
    .ZN(_22172_));
 OAI21_X1 _51775_ (.A(_22171_),
    .B1(_22162_),
    .B2(_22172_),
    .ZN(_01481_));
 NAND4_X1 _51776_ (.A1(_21786_),
    .A2(_21520_),
    .A3(_22149_),
    .A4(_22142_),
    .ZN(_22173_));
 INV_X1 _51777_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1595]),
    .ZN(_22174_));
 OAI21_X1 _51778_ (.A(_22173_),
    .B1(_22162_),
    .B2(_22174_),
    .ZN(_01482_));
 MUX2_X1 _51779_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1596]),
    .B(_21991_),
    .S(_22168_),
    .Z(_01483_));
 BUF_X16 _51780_ (.A(_08608_),
    .Z(_22175_));
 MUX2_X1 _51781_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1597]),
    .B(_22175_),
    .S(_22168_),
    .Z(_01484_));
 NAND4_X1 _51782_ (.A1(_21786_),
    .A2(_08611_),
    .A3(_22149_),
    .A4(_22142_),
    .ZN(_22176_));
 INV_X1 _51783_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1598]),
    .ZN(_22177_));
 OAI21_X1 _51784_ (.A(_22176_),
    .B1(_22162_),
    .B2(_22177_),
    .ZN(_01485_));
 MUX2_X1 _51785_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1599]),
    .B(_22099_),
    .S(_22168_),
    .Z(_01486_));
 MUX2_X1 _51786_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1600]),
    .B(_22033_),
    .S(_22168_),
    .Z(_01489_));
 MUX2_X1 _51787_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1601]),
    .B(_22034_),
    .S(_22168_),
    .Z(_01490_));
 MUX2_X1 _51788_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1602]),
    .B(_22153_),
    .S(_22168_),
    .Z(_01491_));
 MUX2_X1 _51789_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1603]),
    .B(_22035_),
    .S(_22168_),
    .Z(_01492_));
 NAND4_X2 _51790_ (.A1(_21786_),
    .A2(_08629_),
    .A3(_22149_),
    .A4(_22142_),
    .ZN(_22178_));
 INV_X1 _51791_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1604]),
    .ZN(_22179_));
 OAI21_X1 _51792_ (.A(_22178_),
    .B1(_22162_),
    .B2(_22179_),
    .ZN(_01493_));
 BUF_X4 _51793_ (.A(_08632_),
    .Z(_22180_));
 MUX2_X1 _51794_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1605]),
    .B(_22180_),
    .S(_22168_),
    .Z(_01494_));
 MUX2_X1 _51795_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1606]),
    .B(_21930_),
    .S(_22168_),
    .Z(_01495_));
 MUX2_X1 _51796_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1607]),
    .B(_22077_),
    .S(_22161_),
    .Z(_01496_));
 BUF_X16 _51797_ (.A(_21343_),
    .Z(_22181_));
 MUX2_X1 _51798_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1608]),
    .B(_22181_),
    .S(_22161_),
    .Z(_01497_));
 MUX2_X1 _51799_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1609]),
    .B(_21999_),
    .S(_22161_),
    .Z(_01498_));
 MUX2_X1 _51800_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1610]),
    .B(_22000_),
    .S(_22161_),
    .Z(_01500_));
 NAND4_X1 _51801_ (.A1(_21786_),
    .A2(_22154_),
    .A3(_21983_),
    .A4(_21738_),
    .ZN(_22182_));
 INV_X1 _51802_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1611]),
    .ZN(_22183_));
 OAI21_X1 _51803_ (.A(_22182_),
    .B1(_22162_),
    .B2(_22183_),
    .ZN(_01501_));
 MUX2_X1 _51804_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1612]),
    .B(_21958_),
    .S(_22161_),
    .Z(_01502_));
 MUX2_X1 _51805_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1613]),
    .B(_22157_),
    .S(_22161_),
    .Z(_01503_));
 MUX2_X1 _51806_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1614]),
    .B(_21933_),
    .S(_22161_),
    .Z(_01504_));
 MUX2_X1 _51807_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1615]),
    .B(_21899_),
    .S(_22161_),
    .Z(_01505_));
 MUX2_X1 _51808_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1616]),
    .B(_21977_),
    .S(_22161_),
    .Z(_01506_));
 AND2_X4 _51809_ (.A1(_11031_),
    .A2(_21441_),
    .ZN(_22184_));
 BUF_X8 _51810_ (.A(_22184_),
    .Z(_22185_));
 BUF_X8 _51811_ (.A(_22185_),
    .Z(_22186_));
 MUX2_X1 _51812_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1519]),
    .B(_22104_),
    .S(_22186_),
    .Z(_01398_));
 MUX2_X1 _51813_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1520]),
    .B(_22109_),
    .S(_22186_),
    .Z(_01400_));
 MUX2_X1 _51814_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1521]),
    .B(_21967_),
    .S(_22186_),
    .Z(_01401_));
 BUF_X8 _51815_ (.A(_22184_),
    .Z(_22187_));
 MUX2_X1 _51816_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1522]),
    .B(_22110_),
    .S(_22187_),
    .Z(_01402_));
 BUF_X8 _51817_ (.A(_10805_),
    .Z(_22188_));
 BUF_X8 _51818_ (.A(_11038_),
    .Z(_22189_));
 NAND4_X1 _51819_ (.A1(_22188_),
    .A2(_21418_),
    .A3(_22149_),
    .A4(_22189_),
    .ZN(_22190_));
 INV_X1 _51820_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1523]),
    .ZN(_22191_));
 OAI21_X1 _51821_ (.A(_22190_),
    .B1(_22186_),
    .B2(_22191_),
    .ZN(_01403_));
 MUX2_X1 _51822_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1524]),
    .B(_22136_),
    .S(_22187_),
    .Z(_01404_));
 MUX2_X1 _51823_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1525]),
    .B(_22085_),
    .S(_22187_),
    .Z(_01405_));
 MUX2_X1 _51824_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1526]),
    .B(_21969_),
    .S(_22187_),
    .Z(_01406_));
 NAND4_X1 _51825_ (.A1(_22188_),
    .A2(_21392_),
    .A3(_22149_),
    .A4(_22189_),
    .ZN(_22192_));
 INV_X1 _51826_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1527]),
    .ZN(_22193_));
 OAI21_X1 _51827_ (.A(_22192_),
    .B1(_22186_),
    .B2(_22193_),
    .ZN(_01407_));
 MUX2_X1 _51828_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1528]),
    .B(_21988_),
    .S(_22187_),
    .Z(_01408_));
 MUX2_X1 _51829_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1529]),
    .B(_21971_),
    .S(_22187_),
    .Z(_01409_));
 MUX2_X1 _51830_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1530]),
    .B(_22049_),
    .S(_22187_),
    .Z(_01411_));
 MUX2_X1 _51831_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1531]),
    .B(_22088_),
    .S(_22187_),
    .Z(_01412_));
 MUX2_X1 _51832_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1532]),
    .B(_22120_),
    .S(_22187_),
    .Z(_01413_));
 MUX2_X1 _51833_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1533]),
    .B(_22050_),
    .S(_22187_),
    .Z(_01414_));
 BUF_X8 _51834_ (.A(_22184_),
    .Z(_22194_));
 MUX2_X1 _51835_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1534]),
    .B(_22066_),
    .S(_22194_),
    .Z(_01415_));
 MUX2_X1 _51836_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1535]),
    .B(_22090_),
    .S(_22194_),
    .Z(_01416_));
 MUX2_X1 _51837_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1536]),
    .B(_21948_),
    .S(_22194_),
    .Z(_01417_));
 MUX2_X1 _51838_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1537]),
    .B(_22052_),
    .S(_22194_),
    .Z(_01418_));
 MUX2_X1 _51839_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1538]),
    .B(_22019_),
    .S(_22194_),
    .Z(_01419_));
 NAND4_X1 _51840_ (.A1(_22188_),
    .A2(_10614_),
    .A3(_22149_),
    .A4(_22189_),
    .ZN(_22195_));
 INV_X1 _51841_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1539]),
    .ZN(_22196_));
 OAI21_X1 _51842_ (.A(_22195_),
    .B1(_22186_),
    .B2(_22196_),
    .ZN(_01420_));
 MUX2_X1 _51843_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1540]),
    .B(_22022_),
    .S(_22194_),
    .Z(_01422_));
 BUF_X4 _51844_ (.A(_21856_),
    .Z(_22197_));
 NAND4_X2 _51845_ (.A1(_22188_),
    .A2(_10579_),
    .A3(_22197_),
    .A4(_22189_),
    .ZN(_22198_));
 INV_X4 _51846_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1541]),
    .ZN(_22199_));
 OAI21_X1 _51847_ (.A(_22198_),
    .B1(_22186_),
    .B2(_22199_),
    .ZN(_01423_));
 BUF_X4 _51848_ (.A(_11038_),
    .Z(_22200_));
 NAND4_X1 _51849_ (.A1(_22188_),
    .A2(_08588_),
    .A3(_22197_),
    .A4(_22200_),
    .ZN(_22201_));
 INV_X1 _51850_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1542]),
    .ZN(_22202_));
 OAI21_X1 _51851_ (.A(_22201_),
    .B1(_22186_),
    .B2(_22202_),
    .ZN(_01424_));
 MUX2_X1 _51852_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1543]),
    .B(_22122_),
    .S(_22194_),
    .Z(_01425_));
 MUX2_X1 _51853_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1544]),
    .B(_21919_),
    .S(_22194_),
    .Z(_01426_));
 NAND4_X1 _51854_ (.A1(_22188_),
    .A2(_08597_),
    .A3(_22197_),
    .A4(_22200_),
    .ZN(_22203_));
 INV_X1 _51855_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1545]),
    .ZN(_22204_));
 OAI21_X1 _51856_ (.A(_22203_),
    .B1(_22186_),
    .B2(_22204_),
    .ZN(_01427_));
 MUX2_X1 _51857_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1546]),
    .B(_21952_),
    .S(_22194_),
    .Z(_01428_));
 MUX2_X1 _51858_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1547]),
    .B(_21991_),
    .S(_22194_),
    .Z(_01429_));
 BUF_X8 _51859_ (.A(_22184_),
    .Z(_22205_));
 MUX2_X1 _51860_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1548]),
    .B(_22175_),
    .S(_22205_),
    .Z(_01430_));
 MUX2_X1 _51861_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1549]),
    .B(_21955_),
    .S(_22205_),
    .Z(_01431_));
 MUX2_X1 _51862_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1550]),
    .B(_22099_),
    .S(_22205_),
    .Z(_01433_));
 MUX2_X1 _51863_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1551]),
    .B(_22033_),
    .S(_22205_),
    .Z(_01434_));
 MUX2_X1 _51864_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1552]),
    .B(_22034_),
    .S(_22205_),
    .Z(_01435_));
 MUX2_X1 _51865_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1553]),
    .B(_22153_),
    .S(_22205_),
    .Z(_01436_));
 MUX2_X1 _51866_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1554]),
    .B(_22035_),
    .S(_22205_),
    .Z(_01437_));
 MUX2_X1 _51867_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1555]),
    .B(_22074_),
    .S(_22205_),
    .Z(_01438_));
 MUX2_X1 _51868_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1556]),
    .B(_22180_),
    .S(_22205_),
    .Z(_01439_));
 MUX2_X1 _51869_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1557]),
    .B(_21930_),
    .S(_22205_),
    .Z(_01440_));
 MUX2_X1 _51870_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1558]),
    .B(_22077_),
    .S(_22185_),
    .Z(_01441_));
 NAND4_X1 _51871_ (.A1(_22188_),
    .A2(_22154_),
    .A3(_11039_),
    .A4(_21763_),
    .ZN(_22206_));
 INV_X1 _51872_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1559]),
    .ZN(_22207_));
 OAI21_X1 _51873_ (.A(_22206_),
    .B1(_22186_),
    .B2(_22207_),
    .ZN(_01442_));
 MUX2_X1 _51874_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1560]),
    .B(_21999_),
    .S(_22185_),
    .Z(_01444_));
 MUX2_X1 _51875_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1561]),
    .B(_22000_),
    .S(_22185_),
    .Z(_01445_));
 MUX2_X1 _51876_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1562]),
    .B(_22061_),
    .S(_22185_),
    .Z(_01446_));
 BUF_X8 _51877_ (.A(_21359_),
    .Z(_22208_));
 MUX2_X1 _51878_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1563]),
    .B(_22208_),
    .S(_22185_),
    .Z(_01447_));
 MUX2_X1 _51879_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1564]),
    .B(_22157_),
    .S(_22185_),
    .Z(_01448_));
 BUF_X8 _51880_ (.A(_21369_),
    .Z(_22209_));
 MUX2_X1 _51881_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1565]),
    .B(_22209_),
    .S(_22185_),
    .Z(_01449_));
 MUX2_X1 _51882_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1566]),
    .B(_21899_),
    .S(_22185_),
    .Z(_01450_));
 MUX2_X1 _51883_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1567]),
    .B(_21977_),
    .S(_22185_),
    .Z(_01451_));
 BUF_X8 _51884_ (.A(_11041_),
    .Z(_22210_));
 AND2_X4 _51885_ (.A1(_22210_),
    .A2(_21679_),
    .ZN(_22211_));
 BUF_X8 _51886_ (.A(_22211_),
    .Z(_22212_));
 BUF_X8 _51887_ (.A(_22212_),
    .Z(_22213_));
 MUX2_X1 _51888_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1470]),
    .B(_22104_),
    .S(_22213_),
    .Z(_01344_));
 MUX2_X1 _51889_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1471]),
    .B(_22109_),
    .S(_22213_),
    .Z(_01345_));
 BUF_X8 _51890_ (.A(_21294_),
    .Z(_22214_));
 MUX2_X1 _51891_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1472]),
    .B(_22214_),
    .S(_22213_),
    .Z(_01346_));
 MUX2_X1 _51892_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1473]),
    .B(_22110_),
    .S(_22213_),
    .Z(_01347_));
 NAND4_X1 _51893_ (.A1(_22041_),
    .A2(_21418_),
    .A3(_22197_),
    .A4(_22200_),
    .ZN(_22215_));
 INV_X1 _51894_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1474]),
    .ZN(_22216_));
 OAI21_X1 _51895_ (.A(_22215_),
    .B1(_22213_),
    .B2(_22216_),
    .ZN(_01348_));
 BUF_X8 _51896_ (.A(_22211_),
    .Z(_22217_));
 MUX2_X1 _51897_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1475]),
    .B(_22136_),
    .S(_22217_),
    .Z(_01349_));
 MUX2_X1 _51898_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1476]),
    .B(_22085_),
    .S(_22217_),
    .Z(_01350_));
 MUX2_X1 _51899_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1477]),
    .B(_21969_),
    .S(_22217_),
    .Z(_01351_));
 NAND4_X1 _51900_ (.A1(_22041_),
    .A2(_21392_),
    .A3(_22197_),
    .A4(_22200_),
    .ZN(_22218_));
 INV_X1 _51901_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1478]),
    .ZN(_22219_));
 OAI21_X1 _51902_ (.A(_22218_),
    .B1(_22213_),
    .B2(_22219_),
    .ZN(_01352_));
 MUX2_X1 _51903_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1479]),
    .B(_21988_),
    .S(_22217_),
    .Z(_01353_));
 MUX2_X1 _51904_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1480]),
    .B(_21971_),
    .S(_22217_),
    .Z(_01355_));
 MUX2_X1 _51905_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1481]),
    .B(_22049_),
    .S(_22217_),
    .Z(_01356_));
 MUX2_X1 _51906_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1482]),
    .B(_22088_),
    .S(_22217_),
    .Z(_01357_));
 MUX2_X1 _51907_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1483]),
    .B(_22120_),
    .S(_22217_),
    .Z(_01358_));
 MUX2_X1 _51908_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1484]),
    .B(_22050_),
    .S(_22217_),
    .Z(_01359_));
 MUX2_X1 _51909_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1485]),
    .B(_22066_),
    .S(_22217_),
    .Z(_01360_));
 BUF_X8 _51910_ (.A(_22211_),
    .Z(_22220_));
 MUX2_X1 _51911_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1486]),
    .B(_22090_),
    .S(_22220_),
    .Z(_01361_));
 BUF_X8 _51912_ (.A(_08567_),
    .Z(_22221_));
 MUX2_X1 _51913_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1487]),
    .B(_22221_),
    .S(_22220_),
    .Z(_01362_));
 MUX2_X1 _51914_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1488]),
    .B(_22052_),
    .S(_22220_),
    .Z(_01363_));
 MUX2_X1 _51915_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1489]),
    .B(_22019_),
    .S(_22220_),
    .Z(_01364_));
 NAND4_X1 _51916_ (.A1(_22041_),
    .A2(_10614_),
    .A3(_22197_),
    .A4(_22200_),
    .ZN(_22222_));
 INV_X1 _51917_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1490]),
    .ZN(_22223_));
 OAI21_X1 _51918_ (.A(_22222_),
    .B1(_22213_),
    .B2(_22223_),
    .ZN(_01366_));
 MUX2_X1 _51919_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1491]),
    .B(_22022_),
    .S(_22220_),
    .Z(_01367_));
 MUX2_X1 _51920_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1492]),
    .B(_22023_),
    .S(_22220_),
    .Z(_01368_));
 MUX2_X1 _51921_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1493]),
    .B(_21973_),
    .S(_22220_),
    .Z(_01369_));
 MUX2_X1 _51922_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1494]),
    .B(_22122_),
    .S(_22220_),
    .Z(_01370_));
 MUX2_X1 _51923_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1495]),
    .B(_21919_),
    .S(_22220_),
    .Z(_01371_));
 MUX2_X1 _51924_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1496]),
    .B(_22028_),
    .S(_22220_),
    .Z(_01372_));
 BUF_X8 _51925_ (.A(_22211_),
    .Z(_22224_));
 MUX2_X1 _51926_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1497]),
    .B(_21952_),
    .S(_22224_),
    .Z(_01373_));
 MUX2_X1 _51927_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1498]),
    .B(_21991_),
    .S(_22224_),
    .Z(_01374_));
 MUX2_X1 _51928_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1499]),
    .B(_22175_),
    .S(_22224_),
    .Z(_01375_));
 MUX2_X1 _51929_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1500]),
    .B(_21955_),
    .S(_22224_),
    .Z(_01378_));
 MUX2_X1 _51930_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1501]),
    .B(_22099_),
    .S(_22224_),
    .Z(_01379_));
 MUX2_X1 _51931_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1502]),
    .B(_22033_),
    .S(_22224_),
    .Z(_01380_));
 MUX2_X1 _51932_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1503]),
    .B(_22034_),
    .S(_22224_),
    .Z(_01381_));
 MUX2_X1 _51933_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1504]),
    .B(_22153_),
    .S(_22224_),
    .Z(_01382_));
 MUX2_X1 _51934_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1505]),
    .B(_22035_),
    .S(_22224_),
    .Z(_01383_));
 MUX2_X1 _51935_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1506]),
    .B(_22074_),
    .S(_22224_),
    .Z(_01384_));
 MUX2_X1 _51936_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1507]),
    .B(_22180_),
    .S(_22212_),
    .Z(_01385_));
 NAND4_X1 _51937_ (.A1(_22041_),
    .A2(_21591_),
    .A3(_22197_),
    .A4(_22200_),
    .ZN(_22225_));
 INV_X4 _51938_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1508]),
    .ZN(_22226_));
 OAI21_X1 _51939_ (.A(_22225_),
    .B1(_22213_),
    .B2(_22226_),
    .ZN(_01386_));
 MUX2_X1 _51940_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1509]),
    .B(_22077_),
    .S(_22212_),
    .Z(_01387_));
 NAND4_X1 _51941_ (.A1(_22041_),
    .A2(_22154_),
    .A3(_11039_),
    .A4(_21763_),
    .ZN(_22227_));
 INV_X1 _51942_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1510]),
    .ZN(_22228_));
 OAI21_X1 _51943_ (.A(_22227_),
    .B1(_22213_),
    .B2(_22228_),
    .ZN(_01389_));
 MUX2_X1 _51944_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1511]),
    .B(_21999_),
    .S(_22212_),
    .Z(_01390_));
 MUX2_X1 _51945_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1512]),
    .B(_22000_),
    .S(_22212_),
    .Z(_01391_));
 MUX2_X1 _51946_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1513]),
    .B(_22061_),
    .S(_22212_),
    .Z(_01392_));
 MUX2_X1 _51947_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1514]),
    .B(_22208_),
    .S(_22212_),
    .Z(_01393_));
 NAND4_X1 _51948_ (.A1(_22041_),
    .A2(_22154_),
    .A3(_22189_),
    .A4(_21365_),
    .ZN(_22229_));
 INV_X4 _51949_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1515]),
    .ZN(_22230_));
 OAI21_X1 _51950_ (.A(_22229_),
    .B1(_22213_),
    .B2(_22230_),
    .ZN(_01394_));
 MUX2_X1 _51951_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1516]),
    .B(_22209_),
    .S(_22212_),
    .Z(_01395_));
 MUX2_X1 _51952_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1517]),
    .B(_21899_),
    .S(_22212_),
    .Z(_01396_));
 BUF_X4 _51953_ (.A(_21377_),
    .Z(_22231_));
 MUX2_X1 _51954_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1518]),
    .B(_22231_),
    .S(_22212_),
    .Z(_01397_));
 BUF_X16 _51955_ (.A(_11045_),
    .Z(_22232_));
 AND2_X4 _51956_ (.A1(_22232_),
    .A2(_21432_),
    .ZN(_22233_));
 BUF_X16 _51957_ (.A(_22233_),
    .Z(_22234_));
 BUF_X16 _51958_ (.A(_22234_),
    .Z(_22235_));
 MUX2_X1 _51959_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1421]),
    .B(_22104_),
    .S(_22235_),
    .Z(_01290_));
 MUX2_X1 _51960_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1422]),
    .B(_22109_),
    .S(_22235_),
    .Z(_01291_));
 MUX2_X1 _51961_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1423]),
    .B(_22214_),
    .S(_22235_),
    .Z(_01292_));
 MUX2_X1 _51962_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1424]),
    .B(_22110_),
    .S(_22235_),
    .Z(_01293_));
 MUX2_X1 _51963_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1425]),
    .B(_21968_),
    .S(_22235_),
    .Z(_01294_));
 MUX2_X1 _51964_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1426]),
    .B(_22136_),
    .S(_22235_),
    .Z(_01295_));
 MUX2_X1 _51965_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1427]),
    .B(_22085_),
    .S(_22235_),
    .Z(_01296_));
 MUX2_X1 _51966_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1428]),
    .B(_21969_),
    .S(_22235_),
    .Z(_01297_));
 BUF_X8 _51967_ (.A(_22233_),
    .Z(_22236_));
 MUX2_X1 _51968_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1429]),
    .B(_22012_),
    .S(_22236_),
    .Z(_01298_));
 BUF_X16 _51969_ (.A(_21307_),
    .Z(_22237_));
 MUX2_X1 _51970_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1430]),
    .B(_22237_),
    .S(_22236_),
    .Z(_01300_));
 MUX2_X1 _51971_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1431]),
    .B(_21971_),
    .S(_22236_),
    .Z(_01301_));
 MUX2_X1 _51972_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1432]),
    .B(_22049_),
    .S(_22236_),
    .Z(_01302_));
 MUX2_X1 _51973_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1433]),
    .B(_22088_),
    .S(_22236_),
    .Z(_01303_));
 MUX2_X1 _51974_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1434]),
    .B(_22120_),
    .S(_22236_),
    .Z(_01304_));
 MUX2_X1 _51975_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1435]),
    .B(_22050_),
    .S(_22236_),
    .Z(_01305_));
 MUX2_X1 _51976_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1436]),
    .B(_22066_),
    .S(_22236_),
    .Z(_01306_));
 MUX2_X1 _51977_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1437]),
    .B(_22090_),
    .S(_22236_),
    .Z(_01307_));
 MUX2_X1 _51978_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1438]),
    .B(_22221_),
    .S(_22236_),
    .Z(_01308_));
 BUF_X8 _51979_ (.A(_22233_),
    .Z(_22238_));
 MUX2_X1 _51980_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1439]),
    .B(_22052_),
    .S(_22238_),
    .Z(_01309_));
 MUX2_X1 _51981_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1440]),
    .B(_22019_),
    .S(_22238_),
    .Z(_01311_));
 MUX2_X1 _51982_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1441]),
    .B(_22167_),
    .S(_22238_),
    .Z(_01312_));
 MUX2_X1 _51983_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1442]),
    .B(_22022_),
    .S(_22238_),
    .Z(_01313_));
 MUX2_X1 _51984_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1443]),
    .B(_22023_),
    .S(_22238_),
    .Z(_01314_));
 BUF_X4 _51985_ (.A(_08588_),
    .Z(_22239_));
 MUX2_X1 _51986_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1444]),
    .B(_22239_),
    .S(_22238_),
    .Z(_01315_));
 BUF_X32 _51987_ (.A(_10824_),
    .Z(_22240_));
 BUF_X32 _51988_ (.A(_22240_),
    .Z(_22241_));
 BUF_X32 _51989_ (.A(_22241_),
    .Z(_22242_));
 BUF_X8 _51990_ (.A(_22242_),
    .Z(_22243_));
 NAND4_X1 _51991_ (.A1(_22243_),
    .A2(_22025_),
    .A3(_22197_),
    .A4(_22200_),
    .ZN(_22244_));
 INV_X1 _51992_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1445]),
    .ZN(_22245_));
 OAI21_X1 _51993_ (.A(_22244_),
    .B1(_22235_),
    .B2(_22245_),
    .ZN(_01316_));
 MUX2_X1 _51994_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1446]),
    .B(_21919_),
    .S(_22238_),
    .Z(_01317_));
 NAND4_X1 _51995_ (.A1(_22243_),
    .A2(_08597_),
    .A3(_22197_),
    .A4(_22200_),
    .ZN(_22246_));
 INV_X1 _51996_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1447]),
    .ZN(_22247_));
 OAI21_X1 _51997_ (.A(_22246_),
    .B1(_22235_),
    .B2(_22247_),
    .ZN(_01318_));
 MUX2_X1 _51998_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1448]),
    .B(_21952_),
    .S(_22238_),
    .Z(_01319_));
 BUF_X8 _51999_ (.A(_08604_),
    .Z(_22248_));
 MUX2_X1 _52000_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1449]),
    .B(_22248_),
    .S(_22238_),
    .Z(_01320_));
 MUX2_X1 _52001_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1450]),
    .B(_22175_),
    .S(_22238_),
    .Z(_01322_));
 BUF_X16 _52002_ (.A(_22233_),
    .Z(_22249_));
 MUX2_X1 _52003_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1451]),
    .B(_21955_),
    .S(_22249_),
    .Z(_01323_));
 MUX2_X1 _52004_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1452]),
    .B(_22099_),
    .S(_22249_),
    .Z(_01324_));
 MUX2_X1 _52005_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1453]),
    .B(_22033_),
    .S(_22249_),
    .Z(_01325_));
 MUX2_X1 _52006_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1454]),
    .B(_22034_),
    .S(_22249_),
    .Z(_01326_));
 MUX2_X1 _52007_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1455]),
    .B(_22153_),
    .S(_22249_),
    .Z(_01327_));
 MUX2_X1 _52008_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1456]),
    .B(_22035_),
    .S(_22249_),
    .Z(_01328_));
 MUX2_X1 _52009_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1457]),
    .B(_22074_),
    .S(_22249_),
    .Z(_01329_));
 MUX2_X1 _52010_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1458]),
    .B(_22180_),
    .S(_22249_),
    .Z(_01330_));
 BUF_X4 _52011_ (.A(_08635_),
    .Z(_22250_));
 MUX2_X1 _52012_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1459]),
    .B(_22250_),
    .S(_22249_),
    .Z(_01331_));
 MUX2_X1 _52013_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1460]),
    .B(_22077_),
    .S(_22249_),
    .Z(_01333_));
 MUX2_X1 _52014_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1461]),
    .B(_22181_),
    .S(_22234_),
    .Z(_01334_));
 BUF_X16 _52015_ (.A(_21347_),
    .Z(_22251_));
 MUX2_X1 _52016_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1462]),
    .B(_22251_),
    .S(_22234_),
    .Z(_01335_));
 MUX2_X1 _52017_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1463]),
    .B(_22000_),
    .S(_22234_),
    .Z(_01336_));
 MUX2_X1 _52018_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1464]),
    .B(_22061_),
    .S(_22234_),
    .Z(_01337_));
 MUX2_X1 _52019_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1465]),
    .B(_22208_),
    .S(_22234_),
    .Z(_01338_));
 MUX2_X1 _52020_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1466]),
    .B(_22157_),
    .S(_22234_),
    .Z(_01339_));
 MUX2_X1 _52021_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1467]),
    .B(_22209_),
    .S(_22234_),
    .Z(_01340_));
 BUF_X4 _52022_ (.A(_21373_),
    .Z(_22252_));
 MUX2_X1 _52023_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1468]),
    .B(_22252_),
    .S(_22234_),
    .Z(_01341_));
 MUX2_X1 _52024_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1469]),
    .B(_22231_),
    .S(_22234_),
    .Z(_01342_));
 AND2_X4 _52025_ (.A1(_11050_),
    .A2(_21412_),
    .ZN(_22253_));
 BUF_X16 _52026_ (.A(_22253_),
    .Z(_22254_));
 BUF_X8 _52027_ (.A(_22254_),
    .Z(_22255_));
 MUX2_X1 _52028_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1372]),
    .B(_22104_),
    .S(_22255_),
    .Z(_01235_));
 MUX2_X1 _52029_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1373]),
    .B(_22109_),
    .S(_22255_),
    .Z(_01236_));
 MUX2_X1 _52030_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1374]),
    .B(_22214_),
    .S(_22255_),
    .Z(_01237_));
 MUX2_X1 _52031_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1375]),
    .B(_22110_),
    .S(_22255_),
    .Z(_01238_));
 MUX2_X1 _52032_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1376]),
    .B(_21968_),
    .S(_22255_),
    .Z(_01239_));
 BUF_X8 _52033_ (.A(_22253_),
    .Z(_22256_));
 MUX2_X1 _52034_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1377]),
    .B(_22136_),
    .S(_22256_),
    .Z(_01240_));
 MUX2_X1 _52035_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1378]),
    .B(_22085_),
    .S(_22256_),
    .Z(_01241_));
 BUF_X8 _52036_ (.A(_21303_),
    .Z(_22257_));
 MUX2_X1 _52037_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1379]),
    .B(_22257_),
    .S(_22256_),
    .Z(_01242_));
 NAND4_X1 _52038_ (.A1(_21672_),
    .A2(_21392_),
    .A3(_22197_),
    .A4(_22200_),
    .ZN(_22258_));
 INV_X1 _52039_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1380]),
    .ZN(_22259_));
 OAI21_X1 _52040_ (.A(_22258_),
    .B1(_22255_),
    .B2(_22259_),
    .ZN(_01244_));
 MUX2_X1 _52041_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1381]),
    .B(_22237_),
    .S(_22256_),
    .Z(_01245_));
 BUF_X8 _52042_ (.A(_10845_),
    .Z(_22260_));
 BUF_X4 _52043_ (.A(_21856_),
    .Z(_22261_));
 NAND4_X1 _52044_ (.A1(_22260_),
    .A2(_21309_),
    .A3(_22261_),
    .A4(_22200_),
    .ZN(_22262_));
 INV_X1 _52045_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1382]),
    .ZN(_22263_));
 OAI21_X1 _52046_ (.A(_22262_),
    .B1(_22255_),
    .B2(_22263_),
    .ZN(_01246_));
 BUF_X4 _52047_ (.A(_11038_),
    .Z(_22264_));
 NAND4_X2 _52048_ (.A1(_22260_),
    .A2(_21717_),
    .A3(_22261_),
    .A4(_22264_),
    .ZN(_22265_));
 INV_X1 _52049_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1383]),
    .ZN(_22266_));
 OAI21_X1 _52050_ (.A(_22265_),
    .B1(_22255_),
    .B2(_22266_),
    .ZN(_01247_));
 MUX2_X1 _52051_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1384]),
    .B(_22088_),
    .S(_22256_),
    .Z(_01248_));
 MUX2_X1 _52052_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1385]),
    .B(_22120_),
    .S(_22256_),
    .Z(_01249_));
 MUX2_X1 _52053_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1386]),
    .B(_22050_),
    .S(_22256_),
    .Z(_01250_));
 MUX2_X1 _52054_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1387]),
    .B(_22066_),
    .S(_22256_),
    .Z(_01251_));
 MUX2_X1 _52055_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1388]),
    .B(_22090_),
    .S(_22256_),
    .Z(_01252_));
 MUX2_X1 _52056_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1389]),
    .B(_22221_),
    .S(_22256_),
    .Z(_01253_));
 BUF_X8 _52057_ (.A(_22253_),
    .Z(_22267_));
 MUX2_X1 _52058_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1390]),
    .B(_22052_),
    .S(_22267_),
    .Z(_01255_));
 BUF_X8 _52059_ (.A(_08575_),
    .Z(_22268_));
 MUX2_X1 _52060_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1391]),
    .B(_22268_),
    .S(_22267_),
    .Z(_01256_));
 MUX2_X1 _52061_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1392]),
    .B(_22167_),
    .S(_22267_),
    .Z(_01257_));
 BUF_X8 _52062_ (.A(_08581_),
    .Z(_22269_));
 MUX2_X1 _52063_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1393]),
    .B(_22269_),
    .S(_22267_),
    .Z(_01258_));
 MUX2_X1 _52064_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1394]),
    .B(_22023_),
    .S(_22267_),
    .Z(_01259_));
 MUX2_X1 _52065_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1395]),
    .B(_22239_),
    .S(_22267_),
    .Z(_01260_));
 MUX2_X1 _52066_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1396]),
    .B(_22122_),
    .S(_22267_),
    .Z(_01261_));
 BUF_X8 _52067_ (.A(_08594_),
    .Z(_22270_));
 MUX2_X1 _52068_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1397]),
    .B(_22270_),
    .S(_22267_),
    .Z(_01262_));
 MUX2_X1 _52069_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1398]),
    .B(_22028_),
    .S(_22267_),
    .Z(_01263_));
 BUF_X4 _52070_ (.A(_08600_),
    .Z(_22271_));
 MUX2_X1 _52071_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1399]),
    .B(_22271_),
    .S(_22267_),
    .Z(_01264_));
 BUF_X8 _52072_ (.A(_22253_),
    .Z(_22272_));
 MUX2_X1 _52073_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1400]),
    .B(_22248_),
    .S(_22272_),
    .Z(_01267_));
 MUX2_X1 _52074_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1401]),
    .B(_22175_),
    .S(_22272_),
    .Z(_01268_));
 MUX2_X1 _52075_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1402]),
    .B(_21955_),
    .S(_22272_),
    .Z(_01269_));
 MUX2_X1 _52076_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1403]),
    .B(_22099_),
    .S(_22272_),
    .Z(_01270_));
 BUF_X8 _52077_ (.A(_08617_),
    .Z(_22273_));
 MUX2_X1 _52078_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1404]),
    .B(_22273_),
    .S(_22272_),
    .Z(_01271_));
 BUF_X8 _52079_ (.A(_08620_),
    .Z(_22274_));
 MUX2_X1 _52080_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1405]),
    .B(_22274_),
    .S(_22272_),
    .Z(_01272_));
 MUX2_X1 _52081_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1406]),
    .B(_22153_),
    .S(_22272_),
    .Z(_01273_));
 BUF_X4 _52082_ (.A(_08626_),
    .Z(_22275_));
 MUX2_X1 _52083_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1407]),
    .B(_22275_),
    .S(_22272_),
    .Z(_01274_));
 MUX2_X1 _52084_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1408]),
    .B(_22074_),
    .S(_22272_),
    .Z(_01275_));
 MUX2_X1 _52085_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1409]),
    .B(_22180_),
    .S(_22272_),
    .Z(_01276_));
 MUX2_X1 _52086_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1410]),
    .B(_22250_),
    .S(_22254_),
    .Z(_01278_));
 MUX2_X1 _52087_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1411]),
    .B(_22077_),
    .S(_22254_),
    .Z(_01279_));
 NAND4_X2 _52088_ (.A1(_22260_),
    .A2(_22154_),
    .A3(_22189_),
    .A4(_21343_),
    .ZN(_22276_));
 INV_X1 _52089_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1412]),
    .ZN(_22277_));
 OAI21_X1 _52090_ (.A(_22276_),
    .B1(_22255_),
    .B2(_22277_),
    .ZN(_01280_));
 MUX2_X1 _52091_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1413]),
    .B(_22251_),
    .S(_22254_),
    .Z(_01281_));
 NAND4_X1 _52092_ (.A1(_22260_),
    .A2(_22154_),
    .A3(_22189_),
    .A4(_21351_),
    .ZN(_22278_));
 INV_X1 _52093_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1414]),
    .ZN(_22279_));
 OAI21_X1 _52094_ (.A(_22278_),
    .B1(_22255_),
    .B2(_22279_),
    .ZN(_01282_));
 MUX2_X1 _52095_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1415]),
    .B(_22061_),
    .S(_22254_),
    .Z(_01283_));
 MUX2_X1 _52096_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1416]),
    .B(_22208_),
    .S(_22254_),
    .Z(_01284_));
 MUX2_X1 _52097_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1417]),
    .B(_22157_),
    .S(_22254_),
    .Z(_01285_));
 MUX2_X1 _52098_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1418]),
    .B(_22209_),
    .S(_22254_),
    .Z(_01286_));
 MUX2_X1 _52099_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1419]),
    .B(_22252_),
    .S(_22254_),
    .Z(_01287_));
 MUX2_X1 _52100_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1420]),
    .B(_22231_),
    .S(_22254_),
    .Z(_01289_));
 BUF_X4 _52101_ (.A(_10781_),
    .Z(_22280_));
 NAND4_X1 _52102_ (.A1(_22280_),
    .A2(_21598_),
    .A3(_22261_),
    .A4(_22264_),
    .ZN(_22281_));
 BUF_X16 _52103_ (.A(_11054_),
    .Z(_22282_));
 AND2_X4 _52104_ (.A1(_22282_),
    .A2(_21290_),
    .ZN(_22283_));
 BUF_X8 _52105_ (.A(_22283_),
    .Z(_22284_));
 BUF_X4 _52106_ (.A(_22284_),
    .Z(_22285_));
 INV_X1 _52107_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1323]),
    .ZN(_22286_));
 OAI21_X1 _52108_ (.A(_22281_),
    .B1(_22285_),
    .B2(_22286_),
    .ZN(_01181_));
 MUX2_X1 _52109_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1324]),
    .B(_22109_),
    .S(_22284_),
    .Z(_01182_));
 MUX2_X1 _52110_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1325]),
    .B(_22214_),
    .S(_22284_),
    .Z(_01183_));
 MUX2_X1 _52111_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1326]),
    .B(_22110_),
    .S(_22284_),
    .Z(_01184_));
 MUX2_X1 _52112_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1327]),
    .B(_21968_),
    .S(_22284_),
    .Z(_01185_));
 MUX2_X1 _52113_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1328]),
    .B(_22136_),
    .S(_22284_),
    .Z(_01186_));
 MUX2_X1 _52114_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1329]),
    .B(_22085_),
    .S(_22284_),
    .Z(_01187_));
 MUX2_X1 _52115_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1330]),
    .B(_22257_),
    .S(_22284_),
    .Z(_01189_));
 MUX2_X1 _52116_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1331]),
    .B(_22012_),
    .S(_22284_),
    .Z(_01190_));
 MUX2_X1 _52117_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1332]),
    .B(_22237_),
    .S(_22284_),
    .Z(_01191_));
 BUF_X8 _52118_ (.A(_21309_),
    .Z(_22287_));
 BUF_X8 _52119_ (.A(_22283_),
    .Z(_22288_));
 MUX2_X1 _52120_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1333]),
    .B(_22287_),
    .S(_22288_),
    .Z(_01192_));
 MUX2_X1 _52121_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1334]),
    .B(_22049_),
    .S(_22288_),
    .Z(_01193_));
 NAND4_X1 _52122_ (.A1(_22280_),
    .A2(_10563_),
    .A3(_22261_),
    .A4(_22264_),
    .ZN(_22289_));
 INV_X1 _52123_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1335]),
    .ZN(_22290_));
 OAI21_X1 _52124_ (.A(_22289_),
    .B1(_22285_),
    .B2(_22290_),
    .ZN(_01194_));
 NAND4_X1 _52125_ (.A1(_22280_),
    .A2(_08555_),
    .A3(_22261_),
    .A4(_22264_),
    .ZN(_22291_));
 INV_X1 _52126_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1336]),
    .ZN(_22292_));
 OAI21_X1 _52127_ (.A(_22291_),
    .B1(_22285_),
    .B2(_22292_),
    .ZN(_01195_));
 BUF_X8 _52128_ (.A(_08558_),
    .Z(_22293_));
 MUX2_X1 _52129_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1337]),
    .B(_22293_),
    .S(_22288_),
    .Z(_01196_));
 MUX2_X1 _52130_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1338]),
    .B(_22066_),
    .S(_22288_),
    .Z(_01197_));
 MUX2_X1 _52131_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1339]),
    .B(_22090_),
    .S(_22288_),
    .Z(_01198_));
 MUX2_X1 _52132_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1340]),
    .B(_22221_),
    .S(_22288_),
    .Z(_01200_));
 BUF_X4 _52133_ (.A(_08571_),
    .Z(_22294_));
 MUX2_X1 _52134_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1341]),
    .B(_22294_),
    .S(_22288_),
    .Z(_01201_));
 MUX2_X1 _52135_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1342]),
    .B(_22268_),
    .S(_22288_),
    .Z(_01202_));
 MUX2_X1 _52136_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1343]),
    .B(_22167_),
    .S(_22288_),
    .Z(_01203_));
 NAND4_X1 _52137_ (.A1(_22280_),
    .A2(_10578_),
    .A3(_22261_),
    .A4(_22264_),
    .ZN(_22295_));
 INV_X1 _52138_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1344]),
    .ZN(_22296_));
 OAI21_X1 _52139_ (.A(_22295_),
    .B1(_22285_),
    .B2(_22296_),
    .ZN(_01204_));
 BUF_X8 _52140_ (.A(_08584_),
    .Z(_22297_));
 MUX2_X1 _52141_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1345]),
    .B(_22297_),
    .S(_22288_),
    .Z(_01205_));
 BUF_X16 _52142_ (.A(_22283_),
    .Z(_22298_));
 MUX2_X1 _52143_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1346]),
    .B(_22239_),
    .S(_22298_),
    .Z(_01206_));
 NAND4_X1 _52144_ (.A1(_22280_),
    .A2(_22025_),
    .A3(_22261_),
    .A4(_22264_),
    .ZN(_22299_));
 INV_X1 _52145_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1347]),
    .ZN(_22300_));
 OAI21_X1 _52146_ (.A(_22299_),
    .B1(_22285_),
    .B2(_22300_),
    .ZN(_01207_));
 NAND4_X1 _52147_ (.A1(_22280_),
    .A2(_21757_),
    .A3(_22261_),
    .A4(_22264_),
    .ZN(_22301_));
 INV_X1 _52148_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1348]),
    .ZN(_22302_));
 OAI21_X1 _52149_ (.A(_22301_),
    .B1(_22285_),
    .B2(_22302_),
    .ZN(_01208_));
 MUX2_X1 _52150_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1349]),
    .B(_22028_),
    .S(_22298_),
    .Z(_01209_));
 MUX2_X1 _52151_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1350]),
    .B(_22271_),
    .S(_22298_),
    .Z(_01211_));
 NAND4_X1 _52152_ (.A1(_22280_),
    .A2(_21725_),
    .A3(_22261_),
    .A4(_22264_),
    .ZN(_22303_));
 INV_X1 _52153_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1351]),
    .ZN(_22304_));
 OAI21_X1 _52154_ (.A(_22303_),
    .B1(_22285_),
    .B2(_22304_),
    .ZN(_01212_));
 MUX2_X1 _52155_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1352]),
    .B(_22175_),
    .S(_22298_),
    .Z(_01213_));
 MUX2_X1 _52156_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1353]),
    .B(_21955_),
    .S(_22298_),
    .Z(_01214_));
 MUX2_X1 _52157_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1354]),
    .B(_22099_),
    .S(_22298_),
    .Z(_01215_));
 NAND4_X1 _52158_ (.A1(_22280_),
    .A2(_10603_),
    .A3(_22261_),
    .A4(_22264_),
    .ZN(_22305_));
 INV_X1 _52159_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1355]),
    .ZN(_22306_));
 OAI21_X1 _52160_ (.A(_22305_),
    .B1(_22285_),
    .B2(_22306_),
    .ZN(_01216_));
 MUX2_X1 _52161_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1356]),
    .B(_22274_),
    .S(_22298_),
    .Z(_01217_));
 MUX2_X1 _52162_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1357]),
    .B(_22153_),
    .S(_22298_),
    .Z(_01218_));
 MUX2_X1 _52163_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1358]),
    .B(_22275_),
    .S(_22298_),
    .Z(_01219_));
 MUX2_X1 _52164_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1359]),
    .B(_22074_),
    .S(_22298_),
    .Z(_01220_));
 BUF_X16 _52165_ (.A(_22283_),
    .Z(_22307_));
 MUX2_X1 _52166_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1360]),
    .B(_22180_),
    .S(_22307_),
    .Z(_01222_));
 MUX2_X1 _52167_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1361]),
    .B(_22250_),
    .S(_22307_),
    .Z(_01223_));
 MUX2_X1 _52168_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1362]),
    .B(_22077_),
    .S(_22307_),
    .Z(_01224_));
 MUX2_X1 _52169_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1363]),
    .B(_22181_),
    .S(_22307_),
    .Z(_01225_));
 MUX2_X1 _52170_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1364]),
    .B(_22251_),
    .S(_22307_),
    .Z(_01226_));
 BUF_X8 _52171_ (.A(_21351_),
    .Z(_22308_));
 MUX2_X1 _52172_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1365]),
    .B(_22308_),
    .S(_22307_),
    .Z(_01227_));
 MUX2_X1 _52173_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1366]),
    .B(_22061_),
    .S(_22307_),
    .Z(_01228_));
 NAND4_X1 _52174_ (.A1(_22280_),
    .A2(_22154_),
    .A3(_22189_),
    .A4(_21360_),
    .ZN(_22309_));
 INV_X1 _52175_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1367]),
    .ZN(_22310_));
 OAI21_X1 _52176_ (.A(_22309_),
    .B1(_22285_),
    .B2(_22310_),
    .ZN(_01229_));
 NAND4_X1 _52177_ (.A1(_22280_),
    .A2(_22154_),
    .A3(_22189_),
    .A4(_21365_),
    .ZN(_22311_));
 INV_X2 _52178_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1368]),
    .ZN(_22312_));
 OAI21_X1 _52179_ (.A(_22311_),
    .B1(_22285_),
    .B2(_22312_),
    .ZN(_01230_));
 MUX2_X1 _52180_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1369]),
    .B(_22209_),
    .S(_22307_),
    .Z(_01231_));
 MUX2_X1 _52181_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1370]),
    .B(_22252_),
    .S(_22307_),
    .Z(_01233_));
 MUX2_X1 _52182_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1371]),
    .B(_22231_),
    .S(_22307_),
    .Z(_01234_));
 AND2_X4 _52183_ (.A1(_11059_),
    .A2(_21432_),
    .ZN(_22313_));
 BUF_X8 _52184_ (.A(_22313_),
    .Z(_22314_));
 BUF_X4 _52185_ (.A(_22314_),
    .Z(_22315_));
 MUX2_X1 _52186_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1274]),
    .B(_22104_),
    .S(_22315_),
    .Z(_01126_));
 MUX2_X1 _52187_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1275]),
    .B(_22109_),
    .S(_22315_),
    .Z(_01127_));
 MUX2_X1 _52188_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1276]),
    .B(_22214_),
    .S(_22315_),
    .Z(_01128_));
 MUX2_X1 _52189_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1277]),
    .B(_22110_),
    .S(_22315_),
    .Z(_01129_));
 BUF_X16 _52190_ (.A(_21297_),
    .Z(_22316_));
 MUX2_X1 _52191_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1278]),
    .B(_22316_),
    .S(_22315_),
    .Z(_01130_));
 MUX2_X1 _52192_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1279]),
    .B(_22136_),
    .S(_22315_),
    .Z(_01131_));
 MUX2_X1 _52193_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1280]),
    .B(_22085_),
    .S(_22315_),
    .Z(_01133_));
 BUF_X8 _52194_ (.A(_22313_),
    .Z(_22317_));
 MUX2_X1 _52195_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1281]),
    .B(_22257_),
    .S(_22317_),
    .Z(_01134_));
 MUX2_X1 _52196_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1282]),
    .B(_22012_),
    .S(_22317_),
    .Z(_01135_));
 MUX2_X1 _52197_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1283]),
    .B(_22237_),
    .S(_22317_),
    .Z(_01136_));
 MUX2_X1 _52198_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1284]),
    .B(_22287_),
    .S(_22317_),
    .Z(_01137_));
 MUX2_X1 _52199_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1285]),
    .B(_22049_),
    .S(_22317_),
    .Z(_01138_));
 MUX2_X1 _52200_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1286]),
    .B(_22088_),
    .S(_22317_),
    .Z(_01139_));
 MUX2_X1 _52201_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1287]),
    .B(_22120_),
    .S(_22317_),
    .Z(_01140_));
 MUX2_X1 _52202_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1288]),
    .B(_22293_),
    .S(_22317_),
    .Z(_01141_));
 MUX2_X1 _52203_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1289]),
    .B(_22066_),
    .S(_22317_),
    .Z(_01142_));
 MUX2_X1 _52204_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1290]),
    .B(_22090_),
    .S(_22317_),
    .Z(_01144_));
 BUF_X8 _52205_ (.A(_22313_),
    .Z(_22318_));
 MUX2_X1 _52206_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1291]),
    .B(_22221_),
    .S(_22318_),
    .Z(_01145_));
 MUX2_X1 _52207_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1292]),
    .B(_22294_),
    .S(_22318_),
    .Z(_01146_));
 MUX2_X1 _52208_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1293]),
    .B(_22268_),
    .S(_22318_),
    .Z(_01147_));
 MUX2_X1 _52209_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1294]),
    .B(_22167_),
    .S(_22318_),
    .Z(_01148_));
 BUF_X4 _52210_ (.A(_21856_),
    .Z(_22319_));
 NAND4_X1 _52211_ (.A1(_22112_),
    .A2(_10578_),
    .A3(_22319_),
    .A4(_22264_),
    .ZN(_22320_));
 INV_X1 _52212_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1295]),
    .ZN(_22321_));
 OAI21_X1 _52213_ (.A(_22320_),
    .B1(_22315_),
    .B2(_22321_),
    .ZN(_01149_));
 MUX2_X1 _52214_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1296]),
    .B(_22297_),
    .S(_22318_),
    .Z(_01150_));
 MUX2_X1 _52215_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1297]),
    .B(_22239_),
    .S(_22318_),
    .Z(_01151_));
 BUF_X4 _52216_ (.A(_11038_),
    .Z(_22322_));
 NAND4_X1 _52217_ (.A1(_22112_),
    .A2(_22025_),
    .A3(_22319_),
    .A4(_22322_),
    .ZN(_22323_));
 INV_X1 _52218_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1298]),
    .ZN(_22324_));
 OAI21_X1 _52219_ (.A(_22323_),
    .B1(_22315_),
    .B2(_22324_),
    .ZN(_01152_));
 NAND4_X1 _52220_ (.A1(_22112_),
    .A2(_21757_),
    .A3(_22319_),
    .A4(_22322_),
    .ZN(_22325_));
 INV_X1 _52221_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1299]),
    .ZN(_22326_));
 OAI21_X1 _52222_ (.A(_22325_),
    .B1(_22315_),
    .B2(_22326_),
    .ZN(_01153_));
 MUX2_X1 _52223_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1300]),
    .B(_22028_),
    .S(_22318_),
    .Z(_01156_));
 MUX2_X1 _52224_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1301]),
    .B(_22271_),
    .S(_22318_),
    .Z(_01157_));
 MUX2_X1 _52225_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1302]),
    .B(_22248_),
    .S(_22318_),
    .Z(_01158_));
 MUX2_X1 _52226_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1303]),
    .B(_22175_),
    .S(_22318_),
    .Z(_01159_));
 BUF_X8 _52227_ (.A(_08611_),
    .Z(_22327_));
 BUF_X16 _52228_ (.A(_22313_),
    .Z(_22328_));
 MUX2_X1 _52229_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1304]),
    .B(_22327_),
    .S(_22328_),
    .Z(_01160_));
 MUX2_X1 _52230_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1305]),
    .B(_22099_),
    .S(_22328_),
    .Z(_01161_));
 MUX2_X1 _52231_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1306]),
    .B(_22273_),
    .S(_22328_),
    .Z(_01162_));
 MUX2_X1 _52232_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1307]),
    .B(_22274_),
    .S(_22328_),
    .Z(_01163_));
 MUX2_X1 _52233_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1308]),
    .B(_22153_),
    .S(_22328_),
    .Z(_01164_));
 MUX2_X1 _52234_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1309]),
    .B(_22275_),
    .S(_22328_),
    .Z(_01165_));
 MUX2_X1 _52235_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1310]),
    .B(_22074_),
    .S(_22328_),
    .Z(_01167_));
 MUX2_X1 _52236_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1311]),
    .B(_22180_),
    .S(_22328_),
    .Z(_01168_));
 MUX2_X1 _52237_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1312]),
    .B(_22250_),
    .S(_22328_),
    .Z(_01169_));
 BUF_X16 _52238_ (.A(_21339_),
    .Z(_22329_));
 MUX2_X1 _52239_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1313]),
    .B(_22329_),
    .S(_22328_),
    .Z(_01170_));
 MUX2_X1 _52240_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1314]),
    .B(_22181_),
    .S(_22314_),
    .Z(_01171_));
 MUX2_X1 _52241_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1315]),
    .B(_22251_),
    .S(_22314_),
    .Z(_01172_));
 MUX2_X1 _52242_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1316]),
    .B(_22308_),
    .S(_22314_),
    .Z(_01173_));
 MUX2_X1 _52243_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1317]),
    .B(_22061_),
    .S(_22314_),
    .Z(_01174_));
 MUX2_X1 _52244_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1318]),
    .B(_22208_),
    .S(_22314_),
    .Z(_01175_));
 MUX2_X1 _52245_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1319]),
    .B(_22157_),
    .S(_22314_),
    .Z(_01176_));
 MUX2_X1 _52246_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1320]),
    .B(_22209_),
    .S(_22314_),
    .Z(_01178_));
 MUX2_X1 _52247_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1321]),
    .B(_22252_),
    .S(_22314_),
    .Z(_01179_));
 MUX2_X1 _52248_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1322]),
    .B(_22231_),
    .S(_22314_),
    .Z(_01180_));
 AND2_X4 _52249_ (.A1(_11065_),
    .A2(_21441_),
    .ZN(_22330_));
 BUF_X16 _52250_ (.A(_22330_),
    .Z(_22331_));
 BUF_X4 _52251_ (.A(_22331_),
    .Z(_22332_));
 MUX2_X1 _52252_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1225]),
    .B(_22104_),
    .S(_22332_),
    .Z(_01072_));
 MUX2_X1 _52253_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1226]),
    .B(_22109_),
    .S(_22332_),
    .Z(_01073_));
 NAND4_X1 _52254_ (.A1(_21961_),
    .A2(_21383_),
    .A3(_22319_),
    .A4(_22322_),
    .ZN(_22333_));
 INV_X1 _52255_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1227]),
    .ZN(_22334_));
 OAI21_X1 _52256_ (.A(_22333_),
    .B1(_22332_),
    .B2(_22334_),
    .ZN(_01074_));
 MUX2_X1 _52257_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1228]),
    .B(_22110_),
    .S(_22332_),
    .Z(_01075_));
 BUF_X8 _52258_ (.A(_22330_),
    .Z(_22335_));
 MUX2_X1 _52259_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1229]),
    .B(_22316_),
    .S(_22335_),
    .Z(_01076_));
 MUX2_X1 _52260_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1230]),
    .B(_22136_),
    .S(_22335_),
    .Z(_01078_));
 BUF_X8 _52261_ (.A(_21301_),
    .Z(_22336_));
 MUX2_X1 _52262_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1231]),
    .B(_22336_),
    .S(_22335_),
    .Z(_01079_));
 MUX2_X1 _52263_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1232]),
    .B(_22257_),
    .S(_22335_),
    .Z(_01080_));
 BUF_X16 _52264_ (.A(_21305_),
    .Z(_22337_));
 MUX2_X1 _52265_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1233]),
    .B(_22337_),
    .S(_22335_),
    .Z(_01081_));
 MUX2_X1 _52266_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1234]),
    .B(_22237_),
    .S(_22335_),
    .Z(_01082_));
 MUX2_X1 _52267_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1235]),
    .B(_22287_),
    .S(_22335_),
    .Z(_01083_));
 MUX2_X1 _52268_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1236]),
    .B(_22049_),
    .S(_22335_),
    .Z(_01084_));
 MUX2_X1 _52269_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1237]),
    .B(_22088_),
    .S(_22335_),
    .Z(_01085_));
 MUX2_X1 _52270_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1238]),
    .B(_22120_),
    .S(_22335_),
    .Z(_01086_));
 BUF_X8 _52271_ (.A(_22330_),
    .Z(_22338_));
 MUX2_X1 _52272_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1239]),
    .B(_22293_),
    .S(_22338_),
    .Z(_01087_));
 BUF_X8 _52273_ (.A(_08561_),
    .Z(_22339_));
 MUX2_X1 _52274_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1240]),
    .B(_22339_),
    .S(_22338_),
    .Z(_01089_));
 BUF_X8 _52275_ (.A(_10869_),
    .Z(_22340_));
 NAND4_X1 _52276_ (.A1(_22340_),
    .A2(_10572_),
    .A3(_22319_),
    .A4(_22322_),
    .ZN(_22341_));
 INV_X1 _52277_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1241]),
    .ZN(_22342_));
 OAI21_X1 _52278_ (.A(_22341_),
    .B1(_22332_),
    .B2(_22342_),
    .ZN(_01090_));
 MUX2_X1 _52279_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1242]),
    .B(_22221_),
    .S(_22338_),
    .Z(_01091_));
 MUX2_X1 _52280_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1243]),
    .B(_22294_),
    .S(_22338_),
    .Z(_01092_));
 MUX2_X1 _52281_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1244]),
    .B(_22268_),
    .S(_22338_),
    .Z(_01093_));
 MUX2_X1 _52282_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1245]),
    .B(_22167_),
    .S(_22338_),
    .Z(_01094_));
 NAND4_X1 _52283_ (.A1(_22340_),
    .A2(_10578_),
    .A3(_22319_),
    .A4(_22322_),
    .ZN(_22343_));
 INV_X1 _52284_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1246]),
    .ZN(_22344_));
 OAI21_X1 _52285_ (.A(_22343_),
    .B1(_22332_),
    .B2(_22344_),
    .ZN(_01095_));
 MUX2_X1 _52286_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1247]),
    .B(_22297_),
    .S(_22338_),
    .Z(_01096_));
 MUX2_X1 _52287_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1248]),
    .B(_22239_),
    .S(_22338_),
    .Z(_01097_));
 MUX2_X1 _52288_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1249]),
    .B(_22122_),
    .S(_22338_),
    .Z(_01098_));
 MUX2_X1 _52289_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1250]),
    .B(_22270_),
    .S(_22338_),
    .Z(_01100_));
 BUF_X16 _52290_ (.A(_22330_),
    .Z(_22345_));
 MUX2_X1 _52291_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1251]),
    .B(_22028_),
    .S(_22345_),
    .Z(_01101_));
 NAND4_X4 _52292_ (.A1(_22340_),
    .A2(_21520_),
    .A3(_22319_),
    .A4(_22322_),
    .ZN(_22346_));
 INV_X1 _52293_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1252]),
    .ZN(_22347_));
 OAI21_X1 _52294_ (.A(_22346_),
    .B1(_22332_),
    .B2(_22347_),
    .ZN(_01102_));
 NAND4_X1 _52295_ (.A1(_22340_),
    .A2(_21725_),
    .A3(_22319_),
    .A4(_22322_),
    .ZN(_22348_));
 INV_X1 _52296_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1253]),
    .ZN(_22349_));
 OAI21_X1 _52297_ (.A(_22348_),
    .B1(_22332_),
    .B2(_22349_),
    .ZN(_01103_));
 NAND4_X1 _52298_ (.A1(_22340_),
    .A2(_10616_),
    .A3(_22319_),
    .A4(_22322_),
    .ZN(_22350_));
 INV_X1 _52299_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1254]),
    .ZN(_22351_));
 OAI21_X1 _52300_ (.A(_22350_),
    .B1(_22332_),
    .B2(_22351_),
    .ZN(_01104_));
 MUX2_X1 _52301_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1255]),
    .B(_22327_),
    .S(_22345_),
    .Z(_01105_));
 BUF_X4 _52302_ (.A(_08614_),
    .Z(_22352_));
 MUX2_X1 _52303_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1256]),
    .B(_22352_),
    .S(_22345_),
    .Z(_01106_));
 MUX2_X1 _52304_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1257]),
    .B(_22273_),
    .S(_22345_),
    .Z(_01107_));
 MUX2_X1 _52305_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1258]),
    .B(_22274_),
    .S(_22345_),
    .Z(_01108_));
 NAND4_X1 _52306_ (.A1(_22340_),
    .A2(_21562_),
    .A3(_22319_),
    .A4(_22322_),
    .ZN(_22353_));
 INV_X1 _52307_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1259]),
    .ZN(_22354_));
 OAI21_X1 _52308_ (.A(_22353_),
    .B1(_22332_),
    .B2(_22354_),
    .ZN(_01109_));
 MUX2_X1 _52309_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1260]),
    .B(_22275_),
    .S(_22345_),
    .Z(_01111_));
 MUX2_X1 _52310_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1261]),
    .B(_22074_),
    .S(_22345_),
    .Z(_01112_));
 MUX2_X1 _52311_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1262]),
    .B(_22180_),
    .S(_22345_),
    .Z(_01113_));
 MUX2_X1 _52312_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1263]),
    .B(_22250_),
    .S(_22345_),
    .Z(_01114_));
 MUX2_X1 _52313_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1264]),
    .B(_22329_),
    .S(_22345_),
    .Z(_01115_));
 MUX2_X1 _52314_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1265]),
    .B(_22181_),
    .S(_22331_),
    .Z(_01116_));
 MUX2_X1 _52315_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1266]),
    .B(_22251_),
    .S(_22331_),
    .Z(_01117_));
 MUX2_X1 _52316_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1267]),
    .B(_22308_),
    .S(_22331_),
    .Z(_01118_));
 MUX2_X1 _52317_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1268]),
    .B(_22061_),
    .S(_22331_),
    .Z(_01119_));
 MUX2_X1 _52318_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1269]),
    .B(_22208_),
    .S(_22331_),
    .Z(_01120_));
 MUX2_X1 _52319_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1270]),
    .B(_22157_),
    .S(_22331_),
    .Z(_01122_));
 MUX2_X1 _52320_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1271]),
    .B(_22209_),
    .S(_22331_),
    .Z(_01123_));
 MUX2_X1 _52321_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1272]),
    .B(_22252_),
    .S(_22331_),
    .Z(_01124_));
 MUX2_X1 _52322_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1273]),
    .B(_22231_),
    .S(_22331_),
    .Z(_01125_));
 AND2_X4 _52323_ (.A1(_11069_),
    .A2(_21441_),
    .ZN(_22355_));
 BUF_X16 _52324_ (.A(_22355_),
    .Z(_22356_));
 BUF_X4 _52325_ (.A(_22356_),
    .Z(_22357_));
 MUX2_X1 _52326_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1176]),
    .B(_22104_),
    .S(_22357_),
    .Z(_01017_));
 BUF_X8 _52327_ (.A(_21605_),
    .Z(_22358_));
 MUX2_X1 _52328_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1177]),
    .B(_22358_),
    .S(_22357_),
    .Z(_01018_));
 BUF_X8 _52329_ (.A(_10880_),
    .Z(_22359_));
 BUF_X16 _52330_ (.A(_10784_),
    .Z(_22360_));
 BUF_X4 _52331_ (.A(_22360_),
    .Z(_22361_));
 NAND4_X1 _52332_ (.A1(_22359_),
    .A2(_21383_),
    .A3(_22361_),
    .A4(_22322_),
    .ZN(_22362_));
 INV_X1 _52333_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1178]),
    .ZN(_22363_));
 OAI21_X1 _52334_ (.A(_22362_),
    .B1(_22357_),
    .B2(_22363_),
    .ZN(_01019_));
 BUF_X8 _52335_ (.A(_21608_),
    .Z(_22364_));
 MUX2_X1 _52336_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1179]),
    .B(_22364_),
    .S(_22357_),
    .Z(_01020_));
 BUF_X16 _52337_ (.A(_22355_),
    .Z(_22365_));
 MUX2_X1 _52338_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1180]),
    .B(_22316_),
    .S(_22365_),
    .Z(_01022_));
 MUX2_X1 _52339_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1181]),
    .B(_22136_),
    .S(_22365_),
    .Z(_01023_));
 MUX2_X1 _52340_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1182]),
    .B(_22336_),
    .S(_22365_),
    .Z(_01024_));
 MUX2_X1 _52341_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1183]),
    .B(_22257_),
    .S(_22365_),
    .Z(_01025_));
 NAND4_X1 _52342_ (.A1(_22359_),
    .A2(_21392_),
    .A3(_22361_),
    .A4(_11038_),
    .ZN(_22366_));
 INV_X1 _52343_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1184]),
    .ZN(_22367_));
 OAI21_X1 _52344_ (.A(_22366_),
    .B1(_22357_),
    .B2(_22367_),
    .ZN(_01026_));
 MUX2_X1 _52345_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1185]),
    .B(_22237_),
    .S(_22365_),
    .Z(_01027_));
 MUX2_X1 _52346_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1186]),
    .B(_22287_),
    .S(_22365_),
    .Z(_01028_));
 NAND4_X1 _52347_ (.A1(_22359_),
    .A2(_21717_),
    .A3(_22361_),
    .A4(_11038_),
    .ZN(_22368_));
 INV_X1 _52348_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1187]),
    .ZN(_22369_));
 OAI21_X1 _52349_ (.A(_22368_),
    .B1(_22357_),
    .B2(_22369_),
    .ZN(_01029_));
 BUF_X16 _52350_ (.A(_08551_),
    .Z(_22370_));
 MUX2_X1 _52351_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1188]),
    .B(_22370_),
    .S(_22365_),
    .Z(_01030_));
 MUX2_X1 _52352_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1189]),
    .B(_22120_),
    .S(_22365_),
    .Z(_01031_));
 MUX2_X1 _52353_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1190]),
    .B(_22293_),
    .S(_22365_),
    .Z(_01033_));
 MUX2_X1 _52354_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1191]),
    .B(_22339_),
    .S(_22365_),
    .Z(_01034_));
 BUF_X8 _52355_ (.A(_08564_),
    .Z(_22371_));
 NAND4_X1 _52356_ (.A1(_22359_),
    .A2(_22371_),
    .A3(_22361_),
    .A4(_11038_),
    .ZN(_22372_));
 INV_X1 _52357_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1192]),
    .ZN(_22373_));
 OAI21_X1 _52358_ (.A(_22372_),
    .B1(_22357_),
    .B2(_22373_),
    .ZN(_01035_));
 BUF_X16 _52359_ (.A(_22355_),
    .Z(_22374_));
 MUX2_X1 _52360_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1193]),
    .B(_22221_),
    .S(_22374_),
    .Z(_01036_));
 MUX2_X1 _52361_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1194]),
    .B(_22294_),
    .S(_22374_),
    .Z(_01037_));
 MUX2_X1 _52362_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1195]),
    .B(_22268_),
    .S(_22374_),
    .Z(_01038_));
 MUX2_X1 _52363_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1196]),
    .B(_22167_),
    .S(_22374_),
    .Z(_01039_));
 MUX2_X1 _52364_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1197]),
    .B(_22269_),
    .S(_22374_),
    .Z(_01040_));
 MUX2_X1 _52365_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1198]),
    .B(_22297_),
    .S(_22374_),
    .Z(_01041_));
 MUX2_X1 _52366_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1199]),
    .B(_22239_),
    .S(_22374_),
    .Z(_01042_));
 MUX2_X1 _52367_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1200]),
    .B(_22122_),
    .S(_22374_),
    .Z(_01045_));
 MUX2_X1 _52368_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1201]),
    .B(_22270_),
    .S(_22374_),
    .Z(_01046_));
 MUX2_X1 _52369_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1202]),
    .B(_22028_),
    .S(_22374_),
    .Z(_01047_));
 BUF_X16 _52370_ (.A(_22355_),
    .Z(_22375_));
 MUX2_X1 _52371_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1203]),
    .B(_22271_),
    .S(_22375_),
    .Z(_01048_));
 MUX2_X1 _52372_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1204]),
    .B(_22248_),
    .S(_22375_),
    .Z(_01049_));
 NAND4_X1 _52373_ (.A1(_22359_),
    .A2(_10616_),
    .A3(_22361_),
    .A4(_11038_),
    .ZN(_22376_));
 INV_X1 _52374_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1205]),
    .ZN(_22377_));
 OAI21_X1 _52375_ (.A(_22376_),
    .B1(_22357_),
    .B2(_22377_),
    .ZN(_01050_));
 MUX2_X1 _52376_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1206]),
    .B(_22327_),
    .S(_22375_),
    .Z(_01051_));
 MUX2_X1 _52377_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1207]),
    .B(_22352_),
    .S(_22375_),
    .Z(_01052_));
 MUX2_X1 _52378_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1208]),
    .B(_22273_),
    .S(_22375_),
    .Z(_01053_));
 MUX2_X1 _52379_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1209]),
    .B(_22274_),
    .S(_22375_),
    .Z(_01054_));
 NAND4_X1 _52380_ (.A1(_22359_),
    .A2(_21562_),
    .A3(_22361_),
    .A4(_11038_),
    .ZN(_22378_));
 INV_X1 _52381_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1210]),
    .ZN(_22379_));
 OAI21_X1 _52382_ (.A(_22378_),
    .B1(_22357_),
    .B2(_22379_),
    .ZN(_01056_));
 MUX2_X1 _52383_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1211]),
    .B(_22275_),
    .S(_22375_),
    .Z(_01057_));
 BUF_X16 _52384_ (.A(_08629_),
    .Z(_22380_));
 MUX2_X1 _52385_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1212]),
    .B(_22380_),
    .S(_22375_),
    .Z(_01058_));
 MUX2_X1 _52386_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1213]),
    .B(_22180_),
    .S(_22375_),
    .Z(_01059_));
 MUX2_X1 _52387_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1214]),
    .B(_22250_),
    .S(_22375_),
    .Z(_01060_));
 MUX2_X1 _52388_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1215]),
    .B(_22329_),
    .S(_22356_),
    .Z(_01061_));
 BUF_X16 _52389_ (.A(_11015_),
    .Z(_22381_));
 NAND4_X2 _52390_ (.A1(_22359_),
    .A2(_22381_),
    .A3(_22189_),
    .A4(_21343_),
    .ZN(_22382_));
 INV_X1 _52391_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1216]),
    .ZN(_22383_));
 OAI21_X1 _52392_ (.A(_22382_),
    .B1(_22357_),
    .B2(_22383_),
    .ZN(_01062_));
 MUX2_X1 _52393_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1217]),
    .B(_22251_),
    .S(_22356_),
    .Z(_01063_));
 MUX2_X1 _52394_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1218]),
    .B(_22308_),
    .S(_22356_),
    .Z(_01064_));
 MUX2_X1 _52395_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1219]),
    .B(_22061_),
    .S(_22356_),
    .Z(_01065_));
 MUX2_X1 _52396_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1220]),
    .B(_22208_),
    .S(_22356_),
    .Z(_01067_));
 MUX2_X1 _52397_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1221]),
    .B(_22157_),
    .S(_22356_),
    .Z(_01068_));
 MUX2_X1 _52398_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1222]),
    .B(_22209_),
    .S(_22356_),
    .Z(_01069_));
 MUX2_X1 _52399_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1223]),
    .B(_22252_),
    .S(_22356_),
    .Z(_01070_));
 MUX2_X1 _52400_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1224]),
    .B(_22231_),
    .S(_22356_),
    .Z(_01071_));
 BUF_X8 _52401_ (.A(_21598_),
    .Z(_22384_));
 AND2_X4 _52402_ (.A1(_11075_),
    .A2(_21441_),
    .ZN(_22385_));
 BUF_X16 _52403_ (.A(_22385_),
    .Z(_22386_));
 BUF_X4 _52404_ (.A(_22386_),
    .Z(_22387_));
 MUX2_X1 _52405_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1127]),
    .B(_22384_),
    .S(_22387_),
    .Z(_00963_));
 MUX2_X1 _52406_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1128]),
    .B(_22358_),
    .S(_22387_),
    .Z(_00964_));
 BUF_X4 _52407_ (.A(_11082_),
    .Z(_22388_));
 NAND4_X1 _52408_ (.A1(_22188_),
    .A2(_21383_),
    .A3(_22361_),
    .A4(_22388_),
    .ZN(_22389_));
 INV_X1 _52409_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1129]),
    .ZN(_22390_));
 OAI21_X1 _52410_ (.A(_22389_),
    .B1(_22387_),
    .B2(_22390_),
    .ZN(_00965_));
 MUX2_X1 _52411_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1130]),
    .B(_22364_),
    .S(_22387_),
    .Z(_00967_));
 BUF_X8 _52412_ (.A(_22385_),
    .Z(_22391_));
 MUX2_X1 _52413_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1131]),
    .B(_22316_),
    .S(_22391_),
    .Z(_00968_));
 BUF_X8 _52414_ (.A(_21299_),
    .Z(_22392_));
 MUX2_X1 _52415_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1132]),
    .B(_22392_),
    .S(_22391_),
    .Z(_00969_));
 MUX2_X1 _52416_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1133]),
    .B(_22336_),
    .S(_22391_),
    .Z(_00970_));
 MUX2_X1 _52417_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1134]),
    .B(_22257_),
    .S(_22391_),
    .Z(_00971_));
 NAND4_X1 _52418_ (.A1(_22188_),
    .A2(_21305_),
    .A3(_22361_),
    .A4(_22388_),
    .ZN(_22393_));
 INV_X1 _52419_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1135]),
    .ZN(_22394_));
 OAI21_X1 _52420_ (.A(_22393_),
    .B1(_22387_),
    .B2(_22394_),
    .ZN(_00972_));
 MUX2_X1 _52421_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1136]),
    .B(_22237_),
    .S(_22391_),
    .Z(_00973_));
 NAND4_X1 _52422_ (.A1(_22188_),
    .A2(_21309_),
    .A3(_22361_),
    .A4(_22388_),
    .ZN(_22395_));
 INV_X8 _52423_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1137]),
    .ZN(_22396_));
 OAI21_X1 _52424_ (.A(_22395_),
    .B1(_22387_),
    .B2(_22396_),
    .ZN(_00974_));
 MUX2_X1 _52425_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1138]),
    .B(_22049_),
    .S(_22391_),
    .Z(_00975_));
 MUX2_X1 _52426_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1139]),
    .B(_22370_),
    .S(_22391_),
    .Z(_00976_));
 BUF_X4 _52427_ (.A(_08555_),
    .Z(_22397_));
 MUX2_X1 _52428_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1140]),
    .B(_22397_),
    .S(_22391_),
    .Z(_00978_));
 MUX2_X1 _52429_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1141]),
    .B(_22293_),
    .S(_22391_),
    .Z(_00979_));
 MUX2_X1 _52430_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1142]),
    .B(_22339_),
    .S(_22391_),
    .Z(_00980_));
 BUF_X16 _52431_ (.A(_22385_),
    .Z(_22398_));
 MUX2_X1 _52432_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1143]),
    .B(_22090_),
    .S(_22398_),
    .Z(_00981_));
 MUX2_X1 _52433_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1144]),
    .B(_22221_),
    .S(_22398_),
    .Z(_00982_));
 MUX2_X1 _52434_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1145]),
    .B(_22294_),
    .S(_22398_),
    .Z(_00983_));
 MUX2_X1 _52435_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1146]),
    .B(_22268_),
    .S(_22398_),
    .Z(_00984_));
 MUX2_X1 _52436_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1147]),
    .B(_22167_),
    .S(_22398_),
    .Z(_00985_));
 MUX2_X1 _52437_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1148]),
    .B(_22269_),
    .S(_22398_),
    .Z(_00986_));
 MUX2_X1 _52438_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1149]),
    .B(_22297_),
    .S(_22398_),
    .Z(_00987_));
 MUX2_X1 _52439_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1150]),
    .B(_22239_),
    .S(_22398_),
    .Z(_00989_));
 BUF_X8 _52440_ (.A(_10805_),
    .Z(_22399_));
 NAND4_X1 _52441_ (.A1(_22399_),
    .A2(_22025_),
    .A3(_22361_),
    .A4(_22388_),
    .ZN(_22400_));
 INV_X1 _52442_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1151]),
    .ZN(_22401_));
 OAI21_X1 _52443_ (.A(_22400_),
    .B1(_22387_),
    .B2(_22401_),
    .ZN(_00990_));
 MUX2_X1 _52444_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1152]),
    .B(_22270_),
    .S(_22398_),
    .Z(_00991_));
 MUX2_X1 _52445_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1153]),
    .B(_22028_),
    .S(_22398_),
    .Z(_00992_));
 BUF_X16 _52446_ (.A(_22385_),
    .Z(_22402_));
 MUX2_X1 _52447_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1154]),
    .B(_22271_),
    .S(_22402_),
    .Z(_00993_));
 MUX2_X1 _52448_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1155]),
    .B(_22248_),
    .S(_22402_),
    .Z(_00994_));
 MUX2_X1 _52449_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1156]),
    .B(_22175_),
    .S(_22402_),
    .Z(_00995_));
 MUX2_X1 _52450_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1157]),
    .B(_22327_),
    .S(_22402_),
    .Z(_00996_));
 MUX2_X1 _52451_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1158]),
    .B(_22352_),
    .S(_22402_),
    .Z(_00997_));
 MUX2_X1 _52452_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1159]),
    .B(_22273_),
    .S(_22402_),
    .Z(_00998_));
 MUX2_X1 _52453_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1160]),
    .B(_22274_),
    .S(_22402_),
    .Z(_01000_));
 MUX2_X1 _52454_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1161]),
    .B(_22153_),
    .S(_22402_),
    .Z(_01001_));
 MUX2_X1 _52455_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1162]),
    .B(_22275_),
    .S(_22402_),
    .Z(_01002_));
 MUX2_X1 _52456_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1163]),
    .B(_22380_),
    .S(_22402_),
    .Z(_01003_));
 MUX2_X1 _52457_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1164]),
    .B(_22180_),
    .S(_22386_),
    .Z(_01004_));
 BUF_X4 _52458_ (.A(_22360_),
    .Z(_22403_));
 NAND4_X1 _52459_ (.A1(_22399_),
    .A2(_21591_),
    .A3(_22403_),
    .A4(_22388_),
    .ZN(_22404_));
 INV_X4 _52460_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1165]),
    .ZN(_22405_));
 OAI21_X1 _52461_ (.A(_22404_),
    .B1(_22387_),
    .B2(_22405_),
    .ZN(_01005_));
 NAND4_X2 _52462_ (.A1(_22399_),
    .A2(_22381_),
    .A3(_11083_),
    .A4(_21339_),
    .ZN(_22406_));
 INV_X1 _52463_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1166]),
    .ZN(_22407_));
 OAI21_X1 _52464_ (.A(_22406_),
    .B1(_22387_),
    .B2(_22407_),
    .ZN(_01006_));
 MUX2_X1 _52465_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1167]),
    .B(_22181_),
    .S(_22386_),
    .Z(_01007_));
 MUX2_X1 _52466_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1168]),
    .B(_22251_),
    .S(_22386_),
    .Z(_01008_));
 MUX2_X1 _52467_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1169]),
    .B(_22308_),
    .S(_22386_),
    .Z(_01009_));
 NAND4_X2 _52468_ (.A1(_22399_),
    .A2(_22381_),
    .A3(_11083_),
    .A4(_21738_),
    .ZN(_22408_));
 INV_X1 _52469_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1170]),
    .ZN(_22409_));
 OAI21_X1 _52470_ (.A(_22408_),
    .B1(_22387_),
    .B2(_22409_),
    .ZN(_01011_));
 MUX2_X1 _52471_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1171]),
    .B(_22208_),
    .S(_22386_),
    .Z(_01012_));
 MUX2_X1 _52472_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1172]),
    .B(_22157_),
    .S(_22386_),
    .Z(_01013_));
 MUX2_X1 _52473_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1173]),
    .B(_22209_),
    .S(_22386_),
    .Z(_01014_));
 MUX2_X1 _52474_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1174]),
    .B(_22252_),
    .S(_22386_),
    .Z(_01015_));
 MUX2_X1 _52475_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1175]),
    .B(_22231_),
    .S(_22386_),
    .Z(_01016_));
 BUF_X16 _52476_ (.A(_11085_),
    .Z(_22410_));
 AND2_X4 _52477_ (.A1(_22410_),
    .A2(_21679_),
    .ZN(_22411_));
 BUF_X8 _52478_ (.A(_22411_),
    .Z(_22412_));
 BUF_X4 _52479_ (.A(_22412_),
    .Z(_22413_));
 MUX2_X1 _52480_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1078]),
    .B(_22384_),
    .S(_22413_),
    .Z(_00908_));
 MUX2_X1 _52481_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1079]),
    .B(_22358_),
    .S(_22413_),
    .Z(_00909_));
 BUF_X4 _52482_ (.A(_11082_),
    .Z(_22414_));
 NAND4_X1 _52483_ (.A1(_22041_),
    .A2(_21383_),
    .A3(_22403_),
    .A4(_22414_),
    .ZN(_22415_));
 INV_X1 _52484_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1080]),
    .ZN(_22416_));
 OAI21_X1 _52485_ (.A(_22415_),
    .B1(_22413_),
    .B2(_22416_),
    .ZN(_00911_));
 MUX2_X1 _52486_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1081]),
    .B(_22364_),
    .S(_22413_),
    .Z(_00912_));
 BUF_X8 _52487_ (.A(_22411_),
    .Z(_22417_));
 MUX2_X1 _52488_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1082]),
    .B(_22316_),
    .S(_22417_),
    .Z(_00913_));
 MUX2_X1 _52489_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1083]),
    .B(_22392_),
    .S(_22417_),
    .Z(_00914_));
 MUX2_X1 _52490_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1084]),
    .B(_22336_),
    .S(_22417_),
    .Z(_00915_));
 MUX2_X1 _52491_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1085]),
    .B(_22257_),
    .S(_22417_),
    .Z(_00916_));
 NAND4_X1 _52492_ (.A1(_22041_),
    .A2(_21305_),
    .A3(_22403_),
    .A4(_22414_),
    .ZN(_22418_));
 INV_X1 _52493_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1086]),
    .ZN(_22419_));
 OAI21_X1 _52494_ (.A(_22418_),
    .B1(_22413_),
    .B2(_22419_),
    .ZN(_00917_));
 MUX2_X1 _52495_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1087]),
    .B(_22237_),
    .S(_22417_),
    .Z(_00918_));
 MUX2_X1 _52496_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1088]),
    .B(_22287_),
    .S(_22417_),
    .Z(_00919_));
 NAND4_X2 _52497_ (.A1(_22041_),
    .A2(_21717_),
    .A3(_22403_),
    .A4(_22414_),
    .ZN(_22420_));
 INV_X1 _52498_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1089]),
    .ZN(_22421_));
 OAI21_X1 _52499_ (.A(_22420_),
    .B1(_22413_),
    .B2(_22421_),
    .ZN(_00920_));
 MUX2_X1 _52500_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1090]),
    .B(_22370_),
    .S(_22417_),
    .Z(_00922_));
 MUX2_X1 _52501_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1091]),
    .B(_22397_),
    .S(_22417_),
    .Z(_00923_));
 MUX2_X1 _52502_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1092]),
    .B(_22293_),
    .S(_22417_),
    .Z(_00924_));
 MUX2_X1 _52503_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1093]),
    .B(_22339_),
    .S(_22417_),
    .Z(_00925_));
 BUF_X8 _52504_ (.A(_10819_),
    .Z(_22422_));
 NAND4_X1 _52505_ (.A1(_22422_),
    .A2(_22371_),
    .A3(_22403_),
    .A4(_22414_),
    .ZN(_22423_));
 INV_X1 _52506_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1094]),
    .ZN(_22424_));
 OAI21_X1 _52507_ (.A(_22423_),
    .B1(_22413_),
    .B2(_22424_),
    .ZN(_00926_));
 BUF_X16 _52508_ (.A(_22411_),
    .Z(_22425_));
 MUX2_X1 _52509_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1095]),
    .B(_22221_),
    .S(_22425_),
    .Z(_00927_));
 MUX2_X1 _52510_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1096]),
    .B(_22294_),
    .S(_22425_),
    .Z(_00928_));
 MUX2_X1 _52511_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1097]),
    .B(_22268_),
    .S(_22425_),
    .Z(_00929_));
 MUX2_X1 _52512_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1098]),
    .B(_22167_),
    .S(_22425_),
    .Z(_00930_));
 MUX2_X1 _52513_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1099]),
    .B(_22269_),
    .S(_22425_),
    .Z(_00931_));
 MUX2_X1 _52514_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1100]),
    .B(_22297_),
    .S(_22425_),
    .Z(_00934_));
 MUX2_X1 _52515_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1101]),
    .B(_22239_),
    .S(_22425_),
    .Z(_00935_));
 MUX2_X1 _52516_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1102]),
    .B(_22122_),
    .S(_22425_),
    .Z(_00936_));
 MUX2_X1 _52517_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1103]),
    .B(_22270_),
    .S(_22425_),
    .Z(_00937_));
 BUF_X8 _52518_ (.A(_08597_),
    .Z(_22426_));
 MUX2_X1 _52519_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1104]),
    .B(_22426_),
    .S(_22425_),
    .Z(_00938_));
 BUF_X8 _52520_ (.A(_22411_),
    .Z(_22427_));
 MUX2_X1 _52521_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1105]),
    .B(_22271_),
    .S(_22427_),
    .Z(_00939_));
 MUX2_X1 _52522_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1106]),
    .B(_22248_),
    .S(_22427_),
    .Z(_00940_));
 MUX2_X1 _52523_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1107]),
    .B(_22175_),
    .S(_22427_),
    .Z(_00941_));
 MUX2_X1 _52524_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1108]),
    .B(_22327_),
    .S(_22427_),
    .Z(_00942_));
 MUX2_X1 _52525_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1109]),
    .B(_22352_),
    .S(_22427_),
    .Z(_00943_));
 MUX2_X1 _52526_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1110]),
    .B(_22273_),
    .S(_22427_),
    .Z(_00945_));
 MUX2_X1 _52527_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1111]),
    .B(_22274_),
    .S(_22427_),
    .Z(_00946_));
 MUX2_X1 _52528_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1112]),
    .B(_22153_),
    .S(_22427_),
    .Z(_00947_));
 MUX2_X1 _52529_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1113]),
    .B(_22275_),
    .S(_22427_),
    .Z(_00948_));
 MUX2_X1 _52530_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1114]),
    .B(_22380_),
    .S(_22427_),
    .Z(_00949_));
 BUF_X8 _52531_ (.A(_08632_),
    .Z(_22428_));
 MUX2_X1 _52532_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1115]),
    .B(_22428_),
    .S(_22412_),
    .Z(_00950_));
 MUX2_X1 _52533_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1116]),
    .B(_22250_),
    .S(_22412_),
    .Z(_00951_));
 NAND4_X1 _52534_ (.A1(_22422_),
    .A2(_22381_),
    .A3(_22388_),
    .A4(_21339_),
    .ZN(_22429_));
 INV_X1 _52535_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1117]),
    .ZN(_22430_));
 OAI21_X1 _52536_ (.A(_22429_),
    .B1(_22413_),
    .B2(_22430_),
    .ZN(_00952_));
 NAND4_X1 _52537_ (.A1(_22422_),
    .A2(_22381_),
    .A3(_22388_),
    .A4(_21343_),
    .ZN(_22431_));
 INV_X1 _52538_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1118]),
    .ZN(_22432_));
 OAI21_X1 _52539_ (.A(_22431_),
    .B1(_22413_),
    .B2(_22432_),
    .ZN(_00953_));
 MUX2_X1 _52540_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1119]),
    .B(_22251_),
    .S(_22412_),
    .Z(_00954_));
 MUX2_X1 _52541_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1120]),
    .B(_22308_),
    .S(_22412_),
    .Z(_00956_));
 NAND4_X1 _52542_ (.A1(_22422_),
    .A2(_22381_),
    .A3(_22388_),
    .A4(_21738_),
    .ZN(_22433_));
 INV_X1 _52543_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1121]),
    .ZN(_22434_));
 OAI21_X1 _52544_ (.A(_22433_),
    .B1(_22413_),
    .B2(_22434_),
    .ZN(_00957_));
 MUX2_X1 _52545_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1122]),
    .B(_22208_),
    .S(_22412_),
    .Z(_00958_));
 MUX2_X1 _52546_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1123]),
    .B(_22157_),
    .S(_22412_),
    .Z(_00959_));
 MUX2_X1 _52547_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1124]),
    .B(_22209_),
    .S(_22412_),
    .Z(_00960_));
 MUX2_X1 _52548_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1125]),
    .B(_22252_),
    .S(_22412_),
    .Z(_00961_));
 MUX2_X1 _52549_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1126]),
    .B(_22231_),
    .S(_22412_),
    .Z(_00962_));
 BUF_X8 _52550_ (.A(_11090_),
    .Z(_22435_));
 AND2_X4 _52551_ (.A1(_22435_),
    .A2(_21679_),
    .ZN(_22436_));
 BUF_X8 _52552_ (.A(_22436_),
    .Z(_22437_));
 BUF_X8 _52553_ (.A(_22437_),
    .Z(_22438_));
 MUX2_X1 _52554_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1029]),
    .B(_22384_),
    .S(_22438_),
    .Z(_00854_));
 NAND4_X1 _52555_ (.A1(_22243_),
    .A2(_21605_),
    .A3(_22403_),
    .A4(_22414_),
    .ZN(_22439_));
 INV_X1 _52556_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1030]),
    .ZN(_22440_));
 OAI21_X1 _52557_ (.A(_22439_),
    .B1(_22438_),
    .B2(_22440_),
    .ZN(_00856_));
 NAND4_X1 _52558_ (.A1(_22243_),
    .A2(_21383_),
    .A3(_22403_),
    .A4(_22414_),
    .ZN(_22441_));
 INV_X1 _52559_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1031]),
    .ZN(_22442_));
 OAI21_X1 _52560_ (.A(_22441_),
    .B1(_22438_),
    .B2(_22442_),
    .ZN(_00857_));
 MUX2_X1 _52561_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1032]),
    .B(_22364_),
    .S(_22438_),
    .Z(_00858_));
 MUX2_X1 _52562_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1033]),
    .B(_22316_),
    .S(_22438_),
    .Z(_00859_));
 MUX2_X1 _52563_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1034]),
    .B(_22392_),
    .S(_22438_),
    .Z(_00860_));
 BUF_X8 _52564_ (.A(_22436_),
    .Z(_22443_));
 MUX2_X1 _52565_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1035]),
    .B(_22336_),
    .S(_22443_),
    .Z(_00861_));
 MUX2_X1 _52566_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1036]),
    .B(_22257_),
    .S(_22443_),
    .Z(_00862_));
 NAND4_X1 _52567_ (.A1(_22243_),
    .A2(_21305_),
    .A3(_22403_),
    .A4(_22414_),
    .ZN(_22444_));
 INV_X1 _52568_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1037]),
    .ZN(_22445_));
 OAI21_X1 _52569_ (.A(_22444_),
    .B1(_22438_),
    .B2(_22445_),
    .ZN(_00863_));
 MUX2_X1 _52570_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1038]),
    .B(_22237_),
    .S(_22443_),
    .Z(_00864_));
 MUX2_X1 _52571_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1039]),
    .B(_22287_),
    .S(_22443_),
    .Z(_00865_));
 MUX2_X1 _52572_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1040]),
    .B(_22049_),
    .S(_22443_),
    .Z(_00867_));
 MUX2_X1 _52573_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1041]),
    .B(_22370_),
    .S(_22443_),
    .Z(_00868_));
 MUX2_X1 _52574_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1042]),
    .B(_22397_),
    .S(_22443_),
    .Z(_00869_));
 MUX2_X1 _52575_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1043]),
    .B(_22293_),
    .S(_22443_),
    .Z(_00870_));
 MUX2_X1 _52576_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1044]),
    .B(_22339_),
    .S(_22443_),
    .Z(_00871_));
 NAND4_X1 _52577_ (.A1(_22243_),
    .A2(_22371_),
    .A3(_22403_),
    .A4(_22414_),
    .ZN(_22446_));
 INV_X1 _52578_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1045]),
    .ZN(_22447_));
 OAI21_X1 _52579_ (.A(_22446_),
    .B1(_22438_),
    .B2(_22447_),
    .ZN(_00872_));
 MUX2_X1 _52580_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1046]),
    .B(_22221_),
    .S(_22443_),
    .Z(_00873_));
 BUF_X8 _52581_ (.A(_22436_),
    .Z(_22448_));
 MUX2_X1 _52582_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1047]),
    .B(_22294_),
    .S(_22448_),
    .Z(_00874_));
 MUX2_X1 _52583_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1048]),
    .B(_22268_),
    .S(_22448_),
    .Z(_00875_));
 MUX2_X1 _52584_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1049]),
    .B(_22167_),
    .S(_22448_),
    .Z(_00876_));
 MUX2_X1 _52585_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1050]),
    .B(_22269_),
    .S(_22448_),
    .Z(_00878_));
 MUX2_X1 _52586_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1051]),
    .B(_22297_),
    .S(_22448_),
    .Z(_00879_));
 MUX2_X1 _52587_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1052]),
    .B(_22239_),
    .S(_22448_),
    .Z(_00880_));
 MUX2_X1 _52588_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1053]),
    .B(_22122_),
    .S(_22448_),
    .Z(_00881_));
 MUX2_X1 _52589_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1054]),
    .B(_22270_),
    .S(_22448_),
    .Z(_00882_));
 MUX2_X1 _52590_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1055]),
    .B(_22426_),
    .S(_22448_),
    .Z(_00883_));
 MUX2_X1 _52591_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1056]),
    .B(_22271_),
    .S(_22448_),
    .Z(_00884_));
 BUF_X16 _52592_ (.A(_22436_),
    .Z(_22449_));
 MUX2_X1 _52593_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1057]),
    .B(_22248_),
    .S(_22449_),
    .Z(_00885_));
 MUX2_X1 _52594_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1058]),
    .B(_22175_),
    .S(_22449_),
    .Z(_00886_));
 MUX2_X1 _52595_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1059]),
    .B(_22327_),
    .S(_22449_),
    .Z(_00887_));
 MUX2_X1 _52596_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1060]),
    .B(_22352_),
    .S(_22449_),
    .Z(_00889_));
 MUX2_X1 _52597_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1061]),
    .B(_22273_),
    .S(_22449_),
    .Z(_00890_));
 NAND4_X1 _52598_ (.A1(_22243_),
    .A2(_10604_),
    .A3(_22403_),
    .A4(_22414_),
    .ZN(_22450_));
 INV_X1 _52599_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1062]),
    .ZN(_22451_));
 OAI21_X1 _52600_ (.A(_22450_),
    .B1(_22438_),
    .B2(_22451_),
    .ZN(_00891_));
 BUF_X16 _52601_ (.A(_08623_),
    .Z(_22452_));
 MUX2_X1 _52602_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1063]),
    .B(_22452_),
    .S(_22449_),
    .Z(_00892_));
 MUX2_X1 _52603_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1064]),
    .B(_22275_),
    .S(_22449_),
    .Z(_00893_));
 MUX2_X1 _52604_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1065]),
    .B(_22380_),
    .S(_22449_),
    .Z(_00894_));
 MUX2_X1 _52605_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1066]),
    .B(_22428_),
    .S(_22449_),
    .Z(_00895_));
 MUX2_X1 _52606_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1067]),
    .B(_22250_),
    .S(_22449_),
    .Z(_00896_));
 MUX2_X1 _52607_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1068]),
    .B(_22329_),
    .S(_22437_),
    .Z(_00897_));
 MUX2_X1 _52608_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1069]),
    .B(_22181_),
    .S(_22437_),
    .Z(_00898_));
 MUX2_X1 _52609_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1070]),
    .B(_22251_),
    .S(_22437_),
    .Z(_00900_));
 MUX2_X1 _52610_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1071]),
    .B(_22308_),
    .S(_22437_),
    .Z(_00901_));
 NAND4_X4 _52611_ (.A1(_22243_),
    .A2(_22381_),
    .A3(_22388_),
    .A4(_21738_),
    .ZN(_22453_));
 INV_X1 _52612_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1072]),
    .ZN(_22454_));
 OAI21_X1 _52613_ (.A(_22453_),
    .B1(_22438_),
    .B2(_22454_),
    .ZN(_00902_));
 MUX2_X1 _52614_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1073]),
    .B(_22208_),
    .S(_22437_),
    .Z(_00903_));
 BUF_X4 _52615_ (.A(_21365_),
    .Z(_22455_));
 MUX2_X1 _52616_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1074]),
    .B(_22455_),
    .S(_22437_),
    .Z(_00904_));
 BUF_X4 _52617_ (.A(_21369_),
    .Z(_22456_));
 MUX2_X1 _52618_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1075]),
    .B(_22456_),
    .S(_22437_),
    .Z(_00905_));
 MUX2_X1 _52619_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1076]),
    .B(_22252_),
    .S(_22437_),
    .Z(_00906_));
 MUX2_X1 _52620_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1077]),
    .B(_22231_),
    .S(_22437_),
    .Z(_00907_));
 BUF_X4 _52621_ (.A(_22360_),
    .Z(_22457_));
 NAND4_X1 _52622_ (.A1(_22260_),
    .A2(_21598_),
    .A3(_22457_),
    .A4(_22414_),
    .ZN(_22458_));
 BUF_X16 _52623_ (.A(_11094_),
    .Z(_22459_));
 AND2_X4 _52624_ (.A1(_22459_),
    .A2(_21290_),
    .ZN(_22460_));
 BUF_X8 _52625_ (.A(_22460_),
    .Z(_22461_));
 BUF_X4 _52626_ (.A(_22461_),
    .Z(_22462_));
 INV_X4 _52627_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [980]),
    .ZN(_22463_));
 OAI21_X1 _52628_ (.A(_22458_),
    .B1(_22462_),
    .B2(_22463_),
    .ZN(_03935_));
 MUX2_X1 _52629_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [981]),
    .B(_22358_),
    .S(_22461_),
    .Z(_03936_));
 MUX2_X1 _52630_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [982]),
    .B(_22214_),
    .S(_22461_),
    .Z(_03937_));
 MUX2_X1 _52631_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [983]),
    .B(_22364_),
    .S(_22461_),
    .Z(_03938_));
 MUX2_X1 _52632_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [984]),
    .B(_22316_),
    .S(_22461_),
    .Z(_03939_));
 MUX2_X1 _52633_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [985]),
    .B(_22392_),
    .S(_22461_),
    .Z(_03940_));
 MUX2_X1 _52634_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [986]),
    .B(_22336_),
    .S(_22461_),
    .Z(_03941_));
 MUX2_X1 _52635_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [987]),
    .B(_22257_),
    .S(_22461_),
    .Z(_03942_));
 MUX2_X1 _52636_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [988]),
    .B(_22337_),
    .S(_22461_),
    .Z(_03943_));
 BUF_X16 _52637_ (.A(_22460_),
    .Z(_22464_));
 MUX2_X1 _52638_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [989]),
    .B(_22237_),
    .S(_22464_),
    .Z(_03944_));
 MUX2_X1 _52639_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [990]),
    .B(_22287_),
    .S(_22464_),
    .Z(_03946_));
 BUF_X4 _52640_ (.A(_11082_),
    .Z(_22465_));
 NAND4_X2 _52641_ (.A1(_22260_),
    .A2(_21311_),
    .A3(_22457_),
    .A4(_22465_),
    .ZN(_22466_));
 INV_X1 _52642_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [991]),
    .ZN(_22467_));
 OAI21_X1 _52643_ (.A(_22466_),
    .B1(_22462_),
    .B2(_22467_),
    .ZN(_03947_));
 MUX2_X1 _52644_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [992]),
    .B(_22370_),
    .S(_22464_),
    .Z(_03948_));
 MUX2_X1 _52645_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [993]),
    .B(_22397_),
    .S(_22464_),
    .Z(_03949_));
 MUX2_X1 _52646_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [994]),
    .B(_22293_),
    .S(_22464_),
    .Z(_03950_));
 MUX2_X1 _52647_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [995]),
    .B(_22339_),
    .S(_22464_),
    .Z(_03951_));
 NAND4_X1 _52648_ (.A1(_22260_),
    .A2(_22371_),
    .A3(_22457_),
    .A4(_22465_),
    .ZN(_22468_));
 INV_X1 _52649_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [996]),
    .ZN(_22469_));
 OAI21_X1 _52650_ (.A(_22468_),
    .B1(_22462_),
    .B2(_22469_),
    .ZN(_03952_));
 BUF_X4 _52651_ (.A(_08567_),
    .Z(_22470_));
 MUX2_X1 _52652_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [997]),
    .B(_22470_),
    .S(_22464_),
    .Z(_03953_));
 MUX2_X1 _52653_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [998]),
    .B(_22294_),
    .S(_22464_),
    .Z(_03954_));
 MUX2_X1 _52654_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [999]),
    .B(_22268_),
    .S(_22464_),
    .Z(_03955_));
 BUF_X4 _52655_ (.A(_08578_),
    .Z(_22471_));
 MUX2_X1 _52656_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1000]),
    .B(_22471_),
    .S(_22464_),
    .Z(_00823_));
 BUF_X16 _52657_ (.A(_22460_),
    .Z(_22472_));
 MUX2_X1 _52658_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1001]),
    .B(_22269_),
    .S(_22472_),
    .Z(_00824_));
 MUX2_X1 _52659_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1002]),
    .B(_22297_),
    .S(_22472_),
    .Z(_00825_));
 MUX2_X1 _52660_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1003]),
    .B(_22239_),
    .S(_22472_),
    .Z(_00826_));
 NAND4_X1 _52661_ (.A1(_22260_),
    .A2(_22025_),
    .A3(_22457_),
    .A4(_22465_),
    .ZN(_22473_));
 INV_X1 _52662_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1004]),
    .ZN(_22474_));
 OAI21_X1 _52663_ (.A(_22473_),
    .B1(_22462_),
    .B2(_22474_),
    .ZN(_00827_));
 MUX2_X1 _52664_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1005]),
    .B(_22270_),
    .S(_22472_),
    .Z(_00828_));
 MUX2_X1 _52665_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1006]),
    .B(_22426_),
    .S(_22472_),
    .Z(_00829_));
 NAND4_X1 _52666_ (.A1(_22260_),
    .A2(_08600_),
    .A3(_22457_),
    .A4(_22465_),
    .ZN(_22475_));
 INV_X1 _52667_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1007]),
    .ZN(_22476_));
 OAI21_X1 _52668_ (.A(_22475_),
    .B1(_22462_),
    .B2(_22476_),
    .ZN(_00830_));
 NAND4_X1 _52669_ (.A1(_22260_),
    .A2(_21725_),
    .A3(_22457_),
    .A4(_22465_),
    .ZN(_22477_));
 INV_X1 _52670_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1008]),
    .ZN(_22478_));
 OAI21_X1 _52671_ (.A(_22477_),
    .B1(_22462_),
    .B2(_22478_),
    .ZN(_00831_));
 BUF_X4 _52672_ (.A(_08608_),
    .Z(_22479_));
 MUX2_X1 _52673_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1009]),
    .B(_22479_),
    .S(_22472_),
    .Z(_00832_));
 BUF_X8 _52674_ (.A(_10845_),
    .Z(_22480_));
 NAND4_X1 _52675_ (.A1(_22480_),
    .A2(_08611_),
    .A3(_22457_),
    .A4(_22465_),
    .ZN(_22481_));
 INV_X2 _52676_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1010]),
    .ZN(_22482_));
 OAI21_X1 _52677_ (.A(_22481_),
    .B1(_22462_),
    .B2(_22482_),
    .ZN(_00834_));
 MUX2_X1 _52678_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1011]),
    .B(_22352_),
    .S(_22472_),
    .Z(_00835_));
 NAND4_X1 _52679_ (.A1(_22480_),
    .A2(_10603_),
    .A3(_22457_),
    .A4(_22465_),
    .ZN(_22483_));
 INV_X4 _52680_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1012]),
    .ZN(_22484_));
 OAI21_X1 _52681_ (.A(_22483_),
    .B1(_22462_),
    .B2(_22484_),
    .ZN(_00836_));
 MUX2_X1 _52682_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1013]),
    .B(_22274_),
    .S(_22472_),
    .Z(_00837_));
 MUX2_X1 _52683_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1014]),
    .B(_22452_),
    .S(_22472_),
    .Z(_00838_));
 MUX2_X1 _52684_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1015]),
    .B(_22275_),
    .S(_22472_),
    .Z(_00839_));
 NAND4_X1 _52685_ (.A1(_22480_),
    .A2(_08629_),
    .A3(_22457_),
    .A4(_22465_),
    .ZN(_22485_));
 INV_X1 _52686_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1016]),
    .ZN(_22486_));
 OAI21_X1 _52687_ (.A(_22485_),
    .B1(_22462_),
    .B2(_22486_),
    .ZN(_00840_));
 NAND4_X1 _52688_ (.A1(_22480_),
    .A2(_21330_),
    .A3(_22457_),
    .A4(_22465_),
    .ZN(_22487_));
 INV_X2 _52689_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1017]),
    .ZN(_22488_));
 OAI21_X1 _52690_ (.A(_22487_),
    .B1(_22462_),
    .B2(_22488_),
    .ZN(_00841_));
 BUF_X16 _52691_ (.A(_22460_),
    .Z(_22489_));
 MUX2_X1 _52692_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1018]),
    .B(_22250_),
    .S(_22489_),
    .Z(_00842_));
 MUX2_X1 _52693_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1019]),
    .B(_22329_),
    .S(_22489_),
    .Z(_00843_));
 NAND4_X2 _52694_ (.A1(_22480_),
    .A2(_22381_),
    .A3(_22388_),
    .A4(_21343_),
    .ZN(_22490_));
 INV_X1 _52695_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1020]),
    .ZN(_22491_));
 OAI21_X1 _52696_ (.A(_22490_),
    .B1(_22461_),
    .B2(_22491_),
    .ZN(_00845_));
 MUX2_X1 _52697_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1021]),
    .B(_22251_),
    .S(_22489_),
    .Z(_00846_));
 MUX2_X1 _52698_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1022]),
    .B(_22308_),
    .S(_22489_),
    .Z(_00847_));
 BUF_X8 _52699_ (.A(_21355_),
    .Z(_22492_));
 MUX2_X1 _52700_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1023]),
    .B(_22492_),
    .S(_22489_),
    .Z(_00848_));
 BUF_X8 _52701_ (.A(_21359_),
    .Z(_22493_));
 MUX2_X1 _52702_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1024]),
    .B(_22493_),
    .S(_22489_),
    .Z(_00849_));
 MUX2_X1 _52703_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1025]),
    .B(_22455_),
    .S(_22489_),
    .Z(_00850_));
 MUX2_X1 _52704_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1026]),
    .B(_22456_),
    .S(_22489_),
    .Z(_00851_));
 MUX2_X1 _52705_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1027]),
    .B(_22252_),
    .S(_22489_),
    .Z(_00852_));
 BUF_X4 _52706_ (.A(_21377_),
    .Z(_22494_));
 MUX2_X1 _52707_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1028]),
    .B(_22494_),
    .S(_22489_),
    .Z(_00853_));
 AND2_X4 _52708_ (.A1(_11100_),
    .A2(_21574_),
    .ZN(_22495_));
 BUF_X16 _52709_ (.A(_22495_),
    .Z(_22496_));
 BUF_X8 _52710_ (.A(_22496_),
    .Z(_22497_));
 MUX2_X1 _52711_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [931]),
    .B(_22384_),
    .S(_22497_),
    .Z(_03881_));
 MUX2_X1 _52712_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [932]),
    .B(_22358_),
    .S(_22497_),
    .Z(_03882_));
 MUX2_X1 _52713_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [933]),
    .B(_22214_),
    .S(_22497_),
    .Z(_03883_));
 MUX2_X1 _52714_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [934]),
    .B(_22364_),
    .S(_22497_),
    .Z(_03884_));
 BUF_X8 _52715_ (.A(_10781_),
    .Z(_22498_));
 BUF_X4 _52716_ (.A(_22360_),
    .Z(_22499_));
 NAND4_X1 _52717_ (.A1(_22498_),
    .A2(_21418_),
    .A3(_22499_),
    .A4(_22465_),
    .ZN(_22500_));
 INV_X1 _52718_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [935]),
    .ZN(_22501_));
 OAI21_X1 _52719_ (.A(_22500_),
    .B1(_22497_),
    .B2(_22501_),
    .ZN(_03885_));
 MUX2_X1 _52720_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [936]),
    .B(_22392_),
    .S(_22497_),
    .Z(_03886_));
 MUX2_X1 _52721_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [937]),
    .B(_22336_),
    .S(_22497_),
    .Z(_03887_));
 BUF_X16 _52722_ (.A(_22495_),
    .Z(_22502_));
 MUX2_X1 _52723_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [938]),
    .B(_22257_),
    .S(_22502_),
    .Z(_03888_));
 MUX2_X1 _52724_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [939]),
    .B(_22337_),
    .S(_22502_),
    .Z(_03889_));
 BUF_X16 _52725_ (.A(_21307_),
    .Z(_22503_));
 MUX2_X1 _52726_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [940]),
    .B(_22503_),
    .S(_22502_),
    .Z(_03891_));
 MUX2_X1 _52727_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [941]),
    .B(_22287_),
    .S(_22502_),
    .Z(_03892_));
 BUF_X4 _52728_ (.A(_21311_),
    .Z(_22504_));
 MUX2_X1 _52729_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [942]),
    .B(_22504_),
    .S(_22502_),
    .Z(_03893_));
 MUX2_X1 _52730_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [943]),
    .B(_22370_),
    .S(_22502_),
    .Z(_03894_));
 MUX2_X1 _52731_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [944]),
    .B(_22397_),
    .S(_22502_),
    .Z(_03895_));
 MUX2_X1 _52732_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [945]),
    .B(_22293_),
    .S(_22502_),
    .Z(_03896_));
 MUX2_X1 _52733_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [946]),
    .B(_22339_),
    .S(_22502_),
    .Z(_03897_));
 BUF_X4 _52734_ (.A(_11082_),
    .Z(_22505_));
 NAND4_X2 _52735_ (.A1(_22498_),
    .A2(_22371_),
    .A3(_22499_),
    .A4(_22505_),
    .ZN(_22506_));
 INV_X1 _52736_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [947]),
    .ZN(_22507_));
 OAI21_X1 _52737_ (.A(_22506_),
    .B1(_22497_),
    .B2(_22507_),
    .ZN(_03898_));
 MUX2_X1 _52738_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [948]),
    .B(_22470_),
    .S(_22502_),
    .Z(_03899_));
 BUF_X16 _52739_ (.A(_22495_),
    .Z(_22508_));
 MUX2_X1 _52740_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [949]),
    .B(_22294_),
    .S(_22508_),
    .Z(_03900_));
 MUX2_X1 _52741_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [950]),
    .B(_22268_),
    .S(_22508_),
    .Z(_03902_));
 NAND4_X4 _52742_ (.A1(_22498_),
    .A2(_10614_),
    .A3(_22499_),
    .A4(_22505_),
    .ZN(_22509_));
 INV_X1 _52743_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [951]),
    .ZN(_22510_));
 OAI21_X1 _52744_ (.A(_22509_),
    .B1(_22497_),
    .B2(_22510_),
    .ZN(_03903_));
 MUX2_X1 _52745_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [952]),
    .B(_22269_),
    .S(_22508_),
    .Z(_03904_));
 MUX2_X1 _52746_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [953]),
    .B(_22297_),
    .S(_22508_),
    .Z(_03905_));
 BUF_X8 _52747_ (.A(_08588_),
    .Z(_22511_));
 MUX2_X1 _52748_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [954]),
    .B(_22511_),
    .S(_22508_),
    .Z(_03906_));
 BUF_X8 _52749_ (.A(_08591_),
    .Z(_22512_));
 MUX2_X1 _52750_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [955]),
    .B(_22512_),
    .S(_22508_),
    .Z(_03907_));
 MUX2_X1 _52751_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [956]),
    .B(_22270_),
    .S(_22508_),
    .Z(_03908_));
 MUX2_X1 _52752_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [957]),
    .B(_22426_),
    .S(_22508_),
    .Z(_03909_));
 MUX2_X1 _52753_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [958]),
    .B(_22271_),
    .S(_22508_),
    .Z(_03910_));
 MUX2_X1 _52754_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [959]),
    .B(_22248_),
    .S(_22508_),
    .Z(_03911_));
 BUF_X16 _52755_ (.A(_22495_),
    .Z(_22513_));
 MUX2_X1 _52756_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [960]),
    .B(_22479_),
    .S(_22513_),
    .Z(_03913_));
 MUX2_X1 _52757_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [961]),
    .B(_22327_),
    .S(_22513_),
    .Z(_03914_));
 MUX2_X1 _52758_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [962]),
    .B(_22352_),
    .S(_22513_),
    .Z(_03915_));
 MUX2_X1 _52759_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [963]),
    .B(_22273_),
    .S(_22513_),
    .Z(_03916_));
 MUX2_X1 _52760_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [964]),
    .B(_22274_),
    .S(_22513_),
    .Z(_03917_));
 NAND4_X1 _52761_ (.A1(_22498_),
    .A2(_21562_),
    .A3(_22499_),
    .A4(_22505_),
    .ZN(_22514_));
 INV_X1 _52762_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [965]),
    .ZN(_22515_));
 OAI21_X1 _52763_ (.A(_22514_),
    .B1(_22497_),
    .B2(_22515_),
    .ZN(_03918_));
 MUX2_X1 _52764_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [966]),
    .B(_22275_),
    .S(_22513_),
    .Z(_03919_));
 MUX2_X1 _52765_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [967]),
    .B(_22380_),
    .S(_22513_),
    .Z(_03920_));
 MUX2_X1 _52766_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [968]),
    .B(_22428_),
    .S(_22513_),
    .Z(_03921_));
 MUX2_X1 _52767_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [969]),
    .B(_22250_),
    .S(_22513_),
    .Z(_03922_));
 MUX2_X1 _52768_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [970]),
    .B(_22329_),
    .S(_22513_),
    .Z(_03924_));
 MUX2_X1 _52769_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [971]),
    .B(_22181_),
    .S(_22496_),
    .Z(_03925_));
 BUF_X16 _52770_ (.A(_21347_),
    .Z(_22516_));
 MUX2_X1 _52771_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [972]),
    .B(_22516_),
    .S(_22496_),
    .Z(_03926_));
 MUX2_X1 _52772_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [973]),
    .B(_22308_),
    .S(_22496_),
    .Z(_03927_));
 MUX2_X1 _52773_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [974]),
    .B(_22492_),
    .S(_22496_),
    .Z(_03928_));
 MUX2_X1 _52774_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [975]),
    .B(_22493_),
    .S(_22496_),
    .Z(_03929_));
 MUX2_X1 _52775_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [976]),
    .B(_22455_),
    .S(_22496_),
    .Z(_03930_));
 MUX2_X1 _52776_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [977]),
    .B(_22456_),
    .S(_22496_),
    .Z(_03931_));
 BUF_X8 _52777_ (.A(_21373_),
    .Z(_22517_));
 MUX2_X1 _52778_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [978]),
    .B(_22517_),
    .S(_22496_),
    .Z(_03932_));
 MUX2_X1 _52779_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [979]),
    .B(_22494_),
    .S(_22496_),
    .Z(_03933_));
 AND2_X4 _52780_ (.A1(_11106_),
    .A2(_21412_),
    .ZN(_22518_));
 BUF_X16 _52781_ (.A(_22518_),
    .Z(_22519_));
 BUF_X8 _52782_ (.A(_22519_),
    .Z(_22520_));
 MUX2_X1 _52783_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [882]),
    .B(_22384_),
    .S(_22520_),
    .Z(_03826_));
 MUX2_X1 _52784_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [883]),
    .B(_22358_),
    .S(_22520_),
    .Z(_03827_));
 MUX2_X1 _52785_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [884]),
    .B(_22214_),
    .S(_22520_),
    .Z(_03828_));
 MUX2_X1 _52786_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [885]),
    .B(_22364_),
    .S(_22520_),
    .Z(_03829_));
 BUF_X32 _52787_ (.A(_10854_),
    .Z(_22521_));
 BUF_X32 _52788_ (.A(_22521_),
    .Z(_22522_));
 BUF_X32 _52789_ (.A(_22522_),
    .Z(_22523_));
 BUF_X16 _52790_ (.A(_22523_),
    .Z(_22524_));
 BUF_X8 _52791_ (.A(_22524_),
    .Z(_22525_));
 NAND4_X1 _52792_ (.A1(_22525_),
    .A2(_21418_),
    .A3(_22499_),
    .A4(_22505_),
    .ZN(_22526_));
 INV_X1 _52793_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [886]),
    .ZN(_22527_));
 OAI21_X1 _52794_ (.A(_22526_),
    .B1(_22520_),
    .B2(_22527_),
    .ZN(_03830_));
 MUX2_X1 _52795_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [887]),
    .B(_22392_),
    .S(_22520_),
    .Z(_03831_));
 BUF_X16 _52796_ (.A(_22518_),
    .Z(_22528_));
 MUX2_X1 _52797_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [888]),
    .B(_22336_),
    .S(_22528_),
    .Z(_03832_));
 BUF_X8 _52798_ (.A(_21303_),
    .Z(_22529_));
 MUX2_X1 _52799_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [889]),
    .B(_22529_),
    .S(_22528_),
    .Z(_03833_));
 MUX2_X1 _52800_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [890]),
    .B(_22337_),
    .S(_22528_),
    .Z(_03835_));
 MUX2_X1 _52801_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [891]),
    .B(_22503_),
    .S(_22528_),
    .Z(_03836_));
 MUX2_X1 _52802_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [892]),
    .B(_22287_),
    .S(_22528_),
    .Z(_03837_));
 MUX2_X1 _52803_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [893]),
    .B(_22504_),
    .S(_22528_),
    .Z(_03838_));
 MUX2_X1 _52804_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [894]),
    .B(_22370_),
    .S(_22528_),
    .Z(_03839_));
 MUX2_X1 _52805_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [895]),
    .B(_22397_),
    .S(_22528_),
    .Z(_03840_));
 MUX2_X1 _52806_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [896]),
    .B(_22293_),
    .S(_22528_),
    .Z(_03841_));
 MUX2_X1 _52807_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [897]),
    .B(_22339_),
    .S(_22528_),
    .Z(_03842_));
 NAND4_X2 _52808_ (.A1(_22525_),
    .A2(_22371_),
    .A3(_22499_),
    .A4(_22505_),
    .ZN(_22530_));
 INV_X1 _52809_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [898]),
    .ZN(_22531_));
 OAI21_X1 _52810_ (.A(_22530_),
    .B1(_22520_),
    .B2(_22531_),
    .ZN(_03843_));
 BUF_X16 _52811_ (.A(_22518_),
    .Z(_22532_));
 MUX2_X1 _52812_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [899]),
    .B(_22470_),
    .S(_22532_),
    .Z(_03844_));
 MUX2_X1 _52813_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [900]),
    .B(_22294_),
    .S(_22532_),
    .Z(_03847_));
 BUF_X8 _52814_ (.A(_08575_),
    .Z(_22533_));
 MUX2_X1 _52815_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [901]),
    .B(_22533_),
    .S(_22532_),
    .Z(_03848_));
 MUX2_X1 _52816_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [902]),
    .B(_22471_),
    .S(_22532_),
    .Z(_03849_));
 MUX2_X1 _52817_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [903]),
    .B(_22269_),
    .S(_22532_),
    .Z(_03850_));
 MUX2_X1 _52818_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [904]),
    .B(_22297_),
    .S(_22532_),
    .Z(_03851_));
 MUX2_X1 _52819_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [905]),
    .B(_22511_),
    .S(_22532_),
    .Z(_03852_));
 MUX2_X1 _52820_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [906]),
    .B(_22512_),
    .S(_22532_),
    .Z(_03853_));
 NAND4_X4 _52821_ (.A1(_22525_),
    .A2(_21757_),
    .A3(_22499_),
    .A4(_22505_),
    .ZN(_22534_));
 INV_X1 _52822_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [907]),
    .ZN(_22535_));
 OAI21_X1 _52823_ (.A(_22534_),
    .B1(_22520_),
    .B2(_22535_),
    .ZN(_03854_));
 MUX2_X1 _52824_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [908]),
    .B(_22426_),
    .S(_22532_),
    .Z(_03855_));
 MUX2_X1 _52825_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [909]),
    .B(_22271_),
    .S(_22532_),
    .Z(_03856_));
 NAND4_X1 _52826_ (.A1(_22525_),
    .A2(_21725_),
    .A3(_22499_),
    .A4(_22505_),
    .ZN(_22536_));
 INV_X1 _52827_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [910]),
    .ZN(_22537_));
 OAI21_X1 _52828_ (.A(_22536_),
    .B1(_22520_),
    .B2(_22537_),
    .ZN(_03858_));
 BUF_X16 _52829_ (.A(_22518_),
    .Z(_22538_));
 MUX2_X1 _52830_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [911]),
    .B(_22479_),
    .S(_22538_),
    .Z(_03859_));
 MUX2_X1 _52831_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [912]),
    .B(_22327_),
    .S(_22538_),
    .Z(_03860_));
 MUX2_X1 _52832_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [913]),
    .B(_22352_),
    .S(_22538_),
    .Z(_03861_));
 MUX2_X1 _52833_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [914]),
    .B(_22273_),
    .S(_22538_),
    .Z(_03862_));
 MUX2_X1 _52834_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [915]),
    .B(_22274_),
    .S(_22538_),
    .Z(_03863_));
 NAND4_X1 _52835_ (.A1(_22525_),
    .A2(_21562_),
    .A3(_22499_),
    .A4(_22505_),
    .ZN(_22539_));
 INV_X1 _52836_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [916]),
    .ZN(_22540_));
 OAI21_X1 _52837_ (.A(_22539_),
    .B1(_22520_),
    .B2(_22540_),
    .ZN(_03864_));
 BUF_X8 _52838_ (.A(_08626_),
    .Z(_22541_));
 MUX2_X1 _52839_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [917]),
    .B(_22541_),
    .S(_22538_),
    .Z(_03865_));
 MUX2_X1 _52840_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [918]),
    .B(_22380_),
    .S(_22538_),
    .Z(_03866_));
 MUX2_X1 _52841_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [919]),
    .B(_22428_),
    .S(_22538_),
    .Z(_03867_));
 BUF_X4 _52842_ (.A(_08635_),
    .Z(_22542_));
 MUX2_X1 _52843_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [920]),
    .B(_22542_),
    .S(_22538_),
    .Z(_03869_));
 MUX2_X1 _52844_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [921]),
    .B(_22329_),
    .S(_22538_),
    .Z(_03870_));
 MUX2_X1 _52845_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [922]),
    .B(_22181_),
    .S(_22519_),
    .Z(_03871_));
 MUX2_X1 _52846_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [923]),
    .B(_22516_),
    .S(_22519_),
    .Z(_03872_));
 MUX2_X1 _52847_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [924]),
    .B(_22308_),
    .S(_22519_),
    .Z(_03873_));
 MUX2_X1 _52848_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [925]),
    .B(_22492_),
    .S(_22519_),
    .Z(_03874_));
 MUX2_X1 _52849_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [926]),
    .B(_22493_),
    .S(_22519_),
    .Z(_03875_));
 MUX2_X1 _52850_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [927]),
    .B(_22455_),
    .S(_22519_),
    .Z(_03876_));
 MUX2_X1 _52851_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [928]),
    .B(_22456_),
    .S(_22519_),
    .Z(_03877_));
 MUX2_X1 _52852_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [929]),
    .B(_22517_),
    .S(_22519_),
    .Z(_03878_));
 MUX2_X1 _52853_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [930]),
    .B(_22494_),
    .S(_22519_),
    .Z(_03880_));
 NAND4_X1 _52854_ (.A1(_22340_),
    .A2(_21598_),
    .A3(_22499_),
    .A4(_22505_),
    .ZN(_22543_));
 BUF_X16 _52855_ (.A(_11110_),
    .Z(_22544_));
 AND2_X4 _52856_ (.A1(_22544_),
    .A2(_21290_),
    .ZN(_22545_));
 BUF_X16 _52857_ (.A(_22545_),
    .Z(_22546_));
 BUF_X4 _52858_ (.A(_22546_),
    .Z(_22547_));
 INV_X4 _52859_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [833]),
    .ZN(_22548_));
 OAI21_X1 _52860_ (.A(_22543_),
    .B1(_22547_),
    .B2(_22548_),
    .ZN(_03772_));
 MUX2_X1 _52861_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [834]),
    .B(_22358_),
    .S(_22547_),
    .Z(_03773_));
 MUX2_X1 _52862_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [835]),
    .B(_22214_),
    .S(_22547_),
    .Z(_03774_));
 BUF_X8 _52863_ (.A(_22545_),
    .Z(_22549_));
 MUX2_X1 _52864_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [836]),
    .B(_22364_),
    .S(_22549_),
    .Z(_03775_));
 BUF_X4 _52865_ (.A(_22360_),
    .Z(_22550_));
 NAND4_X1 _52866_ (.A1(_22340_),
    .A2(_21418_),
    .A3(_22550_),
    .A4(_22505_),
    .ZN(_22551_));
 INV_X1 _52867_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [837]),
    .ZN(_22552_));
 OAI21_X1 _52868_ (.A(_22551_),
    .B1(_22547_),
    .B2(_22552_),
    .ZN(_03776_));
 MUX2_X1 _52869_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [838]),
    .B(_22392_),
    .S(_22549_),
    .Z(_03777_));
 MUX2_X1 _52870_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [839]),
    .B(_22336_),
    .S(_22549_),
    .Z(_03778_));
 MUX2_X1 _52871_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [840]),
    .B(_22529_),
    .S(_22549_),
    .Z(_03780_));
 BUF_X4 _52872_ (.A(_11082_),
    .Z(_22553_));
 NAND4_X1 _52873_ (.A1(_22340_),
    .A2(_21305_),
    .A3(_22550_),
    .A4(_22553_),
    .ZN(_22554_));
 INV_X1 _52874_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [841]),
    .ZN(_22555_));
 OAI21_X1 _52875_ (.A(_22554_),
    .B1(_22547_),
    .B2(_22555_),
    .ZN(_03781_));
 MUX2_X1 _52876_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [842]),
    .B(_22503_),
    .S(_22549_),
    .Z(_03782_));
 MUX2_X1 _52877_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [843]),
    .B(_22287_),
    .S(_22549_),
    .Z(_03783_));
 MUX2_X1 _52878_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [844]),
    .B(_22504_),
    .S(_22549_),
    .Z(_03784_));
 MUX2_X1 _52879_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [845]),
    .B(_22370_),
    .S(_22549_),
    .Z(_03785_));
 MUX2_X1 _52880_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [846]),
    .B(_22397_),
    .S(_22549_),
    .Z(_03786_));
 BUF_X8 _52881_ (.A(_08558_),
    .Z(_22556_));
 MUX2_X1 _52882_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [847]),
    .B(_22556_),
    .S(_22549_),
    .Z(_03787_));
 BUF_X16 _52883_ (.A(_22545_),
    .Z(_22557_));
 MUX2_X1 _52884_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [848]),
    .B(_22339_),
    .S(_22557_),
    .Z(_03788_));
 NAND4_X1 _52885_ (.A1(_22340_),
    .A2(_22371_),
    .A3(_22550_),
    .A4(_22553_),
    .ZN(_22558_));
 INV_X1 _52886_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [849]),
    .ZN(_22559_));
 OAI21_X1 _52887_ (.A(_22558_),
    .B1(_22547_),
    .B2(_22559_),
    .ZN(_03789_));
 MUX2_X1 _52888_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [850]),
    .B(_22470_),
    .S(_22557_),
    .Z(_03791_));
 BUF_X8 _52889_ (.A(_08571_),
    .Z(_22560_));
 MUX2_X1 _52890_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [851]),
    .B(_22560_),
    .S(_22557_),
    .Z(_03792_));
 MUX2_X1 _52891_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [852]),
    .B(_22533_),
    .S(_22557_),
    .Z(_03793_));
 MUX2_X1 _52892_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [853]),
    .B(_22471_),
    .S(_22557_),
    .Z(_03794_));
 MUX2_X1 _52893_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [854]),
    .B(_22269_),
    .S(_22557_),
    .Z(_03795_));
 BUF_X8 _52894_ (.A(_08584_),
    .Z(_22561_));
 MUX2_X1 _52895_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [855]),
    .B(_22561_),
    .S(_22557_),
    .Z(_03796_));
 MUX2_X1 _52896_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [856]),
    .B(_22511_),
    .S(_22557_),
    .Z(_03797_));
 MUX2_X1 _52897_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [857]),
    .B(_22512_),
    .S(_22557_),
    .Z(_03798_));
 MUX2_X1 _52898_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [858]),
    .B(_22270_),
    .S(_22557_),
    .Z(_03799_));
 BUF_X16 _52899_ (.A(_22545_),
    .Z(_22562_));
 MUX2_X1 _52900_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [859]),
    .B(_22426_),
    .S(_22562_),
    .Z(_03800_));
 MUX2_X1 _52901_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [860]),
    .B(_22271_),
    .S(_22562_),
    .Z(_03802_));
 BUF_X8 _52902_ (.A(_10869_),
    .Z(_22563_));
 NAND4_X1 _52903_ (.A1(_22563_),
    .A2(_21725_),
    .A3(_22550_),
    .A4(_22553_),
    .ZN(_22564_));
 INV_X1 _52904_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [861]),
    .ZN(_22565_));
 OAI21_X1 _52905_ (.A(_22564_),
    .B1(_22547_),
    .B2(_22565_),
    .ZN(_03803_));
 NAND4_X2 _52906_ (.A1(_22563_),
    .A2(_10616_),
    .A3(_22550_),
    .A4(_22553_),
    .ZN(_22566_));
 INV_X1 _52907_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [862]),
    .ZN(_22567_));
 OAI21_X1 _52908_ (.A(_22566_),
    .B1(_22547_),
    .B2(_22567_),
    .ZN(_03804_));
 MUX2_X1 _52909_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [863]),
    .B(_22327_),
    .S(_22562_),
    .Z(_03805_));
 MUX2_X1 _52910_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [864]),
    .B(_22352_),
    .S(_22562_),
    .Z(_03806_));
 NAND4_X1 _52911_ (.A1(_22563_),
    .A2(_08617_),
    .A3(_22550_),
    .A4(_22553_),
    .ZN(_22568_));
 INV_X4 _52912_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [865]),
    .ZN(_22569_));
 OAI21_X1 _52913_ (.A(_22568_),
    .B1(_22547_),
    .B2(_22569_),
    .ZN(_03807_));
 BUF_X8 _52914_ (.A(_08620_),
    .Z(_22570_));
 MUX2_X1 _52915_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [866]),
    .B(_22570_),
    .S(_22562_),
    .Z(_03808_));
 NAND4_X2 _52916_ (.A1(_22563_),
    .A2(_21562_),
    .A3(_22550_),
    .A4(_22553_),
    .ZN(_22571_));
 INV_X1 _52917_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [867]),
    .ZN(_22572_));
 OAI21_X1 _52918_ (.A(_22571_),
    .B1(_22547_),
    .B2(_22572_),
    .ZN(_03809_));
 MUX2_X1 _52919_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [868]),
    .B(_22541_),
    .S(_22562_),
    .Z(_03810_));
 MUX2_X1 _52920_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [869]),
    .B(_22380_),
    .S(_22562_),
    .Z(_03811_));
 MUX2_X1 _52921_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [870]),
    .B(_22428_),
    .S(_22562_),
    .Z(_03813_));
 MUX2_X1 _52922_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [871]),
    .B(_22542_),
    .S(_22562_),
    .Z(_03814_));
 MUX2_X1 _52923_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [872]),
    .B(_22329_),
    .S(_22562_),
    .Z(_03815_));
 MUX2_X1 _52924_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [873]),
    .B(_22181_),
    .S(_22546_),
    .Z(_03816_));
 MUX2_X1 _52925_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [874]),
    .B(_22516_),
    .S(_22546_),
    .Z(_03817_));
 BUF_X8 _52926_ (.A(_21351_),
    .Z(_22573_));
 MUX2_X1 _52927_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [875]),
    .B(_22573_),
    .S(_22546_),
    .Z(_03818_));
 MUX2_X1 _52928_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [876]),
    .B(_22492_),
    .S(_22546_),
    .Z(_03819_));
 MUX2_X1 _52929_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [877]),
    .B(_22493_),
    .S(_22546_),
    .Z(_03820_));
 MUX2_X1 _52930_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [878]),
    .B(_22455_),
    .S(_22546_),
    .Z(_03821_));
 MUX2_X1 _52931_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [879]),
    .B(_22456_),
    .S(_22546_),
    .Z(_03822_));
 MUX2_X1 _52932_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [880]),
    .B(_22517_),
    .S(_22546_),
    .Z(_03824_));
 MUX2_X1 _52933_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [881]),
    .B(_22494_),
    .S(_22546_),
    .Z(_03825_));
 AND2_X4 _52934_ (.A1(_11114_),
    .A2(_21679_),
    .ZN(_22574_));
 BUF_X16 _52935_ (.A(_22574_),
    .Z(_22575_));
 BUF_X8 _52936_ (.A(_22575_),
    .Z(_22576_));
 MUX2_X1 _52937_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [784]),
    .B(_22384_),
    .S(_22576_),
    .Z(_03717_));
 NAND4_X1 _52938_ (.A1(_22359_),
    .A2(_21605_),
    .A3(_22550_),
    .A4(_22553_),
    .ZN(_22577_));
 INV_X1 _52939_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [785]),
    .ZN(_22578_));
 OAI21_X1 _52940_ (.A(_22577_),
    .B1(_22576_),
    .B2(_22578_),
    .ZN(_03718_));
 MUX2_X1 _52941_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [786]),
    .B(_22214_),
    .S(_22576_),
    .Z(_03719_));
 MUX2_X1 _52942_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [787]),
    .B(_22364_),
    .S(_22576_),
    .Z(_03720_));
 NAND4_X1 _52943_ (.A1(_22359_),
    .A2(_21418_),
    .A3(_22550_),
    .A4(_22553_),
    .ZN(_22579_));
 INV_X1 _52944_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [788]),
    .ZN(_22580_));
 OAI21_X1 _52945_ (.A(_22579_),
    .B1(_22576_),
    .B2(_22580_),
    .ZN(_03721_));
 MUX2_X1 _52946_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [789]),
    .B(_22392_),
    .S(_22576_),
    .Z(_03722_));
 BUF_X8 _52947_ (.A(_22574_),
    .Z(_22581_));
 MUX2_X1 _52948_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [790]),
    .B(_22336_),
    .S(_22581_),
    .Z(_03724_));
 MUX2_X1 _52949_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [791]),
    .B(_22529_),
    .S(_22581_),
    .Z(_03725_));
 MUX2_X1 _52950_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [792]),
    .B(_22337_),
    .S(_22581_),
    .Z(_03726_));
 MUX2_X1 _52951_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [793]),
    .B(_22503_),
    .S(_22581_),
    .Z(_03727_));
 BUF_X8 _52952_ (.A(_21309_),
    .Z(_22582_));
 MUX2_X1 _52953_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [794]),
    .B(_22582_),
    .S(_22581_),
    .Z(_03728_));
 MUX2_X1 _52954_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [795]),
    .B(_22504_),
    .S(_22581_),
    .Z(_03729_));
 MUX2_X1 _52955_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [796]),
    .B(_22370_),
    .S(_22581_),
    .Z(_03730_));
 MUX2_X1 _52956_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [797]),
    .B(_22397_),
    .S(_22581_),
    .Z(_03731_));
 MUX2_X1 _52957_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [798]),
    .B(_22556_),
    .S(_22581_),
    .Z(_03732_));
 MUX2_X1 _52958_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [799]),
    .B(_22339_),
    .S(_22581_),
    .Z(_03733_));
 BUF_X8 _52959_ (.A(_08564_),
    .Z(_22583_));
 BUF_X16 _52960_ (.A(_22574_),
    .Z(_22584_));
 MUX2_X1 _52961_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [800]),
    .B(_22583_),
    .S(_22584_),
    .Z(_03736_));
 MUX2_X1 _52962_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [801]),
    .B(_22470_),
    .S(_22584_),
    .Z(_03737_));
 MUX2_X1 _52963_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [802]),
    .B(_22560_),
    .S(_22584_),
    .Z(_03738_));
 MUX2_X1 _52964_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [803]),
    .B(_22533_),
    .S(_22584_),
    .Z(_03739_));
 MUX2_X1 _52965_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [804]),
    .B(_22471_),
    .S(_22584_),
    .Z(_03740_));
 MUX2_X1 _52966_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [805]),
    .B(_22269_),
    .S(_22584_),
    .Z(_03741_));
 MUX2_X1 _52967_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [806]),
    .B(_22561_),
    .S(_22584_),
    .Z(_03742_));
 MUX2_X1 _52968_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [807]),
    .B(_22511_),
    .S(_22584_),
    .Z(_03743_));
 MUX2_X1 _52969_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [808]),
    .B(_22512_),
    .S(_22584_),
    .Z(_03744_));
 MUX2_X1 _52970_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [809]),
    .B(_22270_),
    .S(_22584_),
    .Z(_03745_));
 BUF_X8 _52971_ (.A(_22574_),
    .Z(_22585_));
 MUX2_X1 _52972_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [810]),
    .B(_22426_),
    .S(_22585_),
    .Z(_03747_));
 NAND4_X1 _52973_ (.A1(_22359_),
    .A2(_08600_),
    .A3(_22550_),
    .A4(_22553_),
    .ZN(_22586_));
 INV_X1 _52974_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [811]),
    .ZN(_22587_));
 OAI21_X1 _52975_ (.A(_22586_),
    .B1(_22576_),
    .B2(_22587_),
    .ZN(_03748_));
 MUX2_X1 _52976_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [812]),
    .B(_22248_),
    .S(_22585_),
    .Z(_03749_));
 BUF_X8 _52977_ (.A(_10880_),
    .Z(_22588_));
 BUF_X8 _52978_ (.A(_22360_),
    .Z(_22589_));
 NAND4_X2 _52979_ (.A1(_22588_),
    .A2(_08608_),
    .A3(_22589_),
    .A4(_22553_),
    .ZN(_22590_));
 INV_X1 _52980_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [813]),
    .ZN(_22591_));
 OAI21_X1 _52981_ (.A(_22590_),
    .B1(_22576_),
    .B2(_22591_),
    .ZN(_03750_));
 MUX2_X1 _52982_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [814]),
    .B(_22327_),
    .S(_22585_),
    .Z(_03751_));
 MUX2_X1 _52983_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [815]),
    .B(_22352_),
    .S(_22585_),
    .Z(_03752_));
 MUX2_X1 _52984_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [816]),
    .B(_22273_),
    .S(_22585_),
    .Z(_03753_));
 NAND4_X1 _52985_ (.A1(_22588_),
    .A2(_08620_),
    .A3(_22589_),
    .A4(_11082_),
    .ZN(_22592_));
 INV_X1 _52986_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [817]),
    .ZN(_22593_));
 OAI21_X1 _52987_ (.A(_22592_),
    .B1(_22576_),
    .B2(_22593_),
    .ZN(_03754_));
 NAND4_X2 _52988_ (.A1(_22588_),
    .A2(_21562_),
    .A3(_22589_),
    .A4(_11082_),
    .ZN(_22594_));
 INV_X1 _52989_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [818]),
    .ZN(_22595_));
 OAI21_X1 _52990_ (.A(_22594_),
    .B1(_22576_),
    .B2(_22595_),
    .ZN(_03755_));
 MUX2_X1 _52991_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [819]),
    .B(_22541_),
    .S(_22585_),
    .Z(_03756_));
 MUX2_X1 _52992_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [820]),
    .B(_22380_),
    .S(_22585_),
    .Z(_03758_));
 MUX2_X1 _52993_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [821]),
    .B(_22428_),
    .S(_22585_),
    .Z(_03759_));
 MUX2_X1 _52994_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [822]),
    .B(_22542_),
    .S(_22585_),
    .Z(_03760_));
 MUX2_X1 _52995_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [823]),
    .B(_22329_),
    .S(_22585_),
    .Z(_03761_));
 BUF_X16 _52996_ (.A(_21343_),
    .Z(_22596_));
 MUX2_X1 _52997_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [824]),
    .B(_22596_),
    .S(_22575_),
    .Z(_03762_));
 MUX2_X1 _52998_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [825]),
    .B(_22516_),
    .S(_22575_),
    .Z(_03763_));
 MUX2_X1 _52999_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [826]),
    .B(_22573_),
    .S(_22575_),
    .Z(_03764_));
 MUX2_X1 _53000_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [827]),
    .B(_22492_),
    .S(_22575_),
    .Z(_03765_));
 MUX2_X1 _53001_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [828]),
    .B(_22493_),
    .S(_22575_),
    .Z(_03766_));
 MUX2_X1 _53002_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [829]),
    .B(_22455_),
    .S(_22575_),
    .Z(_03767_));
 MUX2_X1 _53003_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [830]),
    .B(_22456_),
    .S(_22575_),
    .Z(_03769_));
 MUX2_X1 _53004_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [831]),
    .B(_22517_),
    .S(_22575_),
    .Z(_03770_));
 MUX2_X1 _53005_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [832]),
    .B(_22494_),
    .S(_22575_),
    .Z(_03771_));
 BUF_X8 _53006_ (.A(_11120_),
    .Z(_22597_));
 AND2_X4 _53007_ (.A1(_22597_),
    .A2(_21412_),
    .ZN(_22598_));
 BUF_X8 _53008_ (.A(_22598_),
    .Z(_22599_));
 BUF_X8 _53009_ (.A(_22599_),
    .Z(_22600_));
 MUX2_X1 _53010_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [735]),
    .B(_22384_),
    .S(_22600_),
    .Z(_03663_));
 MUX2_X1 _53011_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [736]),
    .B(_22358_),
    .S(_22600_),
    .Z(_03664_));
 BUF_X4 _53012_ (.A(_21294_),
    .Z(_22601_));
 MUX2_X1 _53013_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [737]),
    .B(_22601_),
    .S(_22600_),
    .Z(_03665_));
 MUX2_X1 _53014_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [738]),
    .B(_22364_),
    .S(_22600_),
    .Z(_03666_));
 BUF_X4 _53015_ (.A(_11127_),
    .Z(_22602_));
 NAND4_X1 _53016_ (.A1(_22399_),
    .A2(_21297_),
    .A3(_22589_),
    .A4(_22602_),
    .ZN(_22603_));
 INV_X1 _53017_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [739]),
    .ZN(_22604_));
 OAI21_X1 _53018_ (.A(_22603_),
    .B1(_22600_),
    .B2(_22604_),
    .ZN(_03667_));
 MUX2_X1 _53019_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [740]),
    .B(_22392_),
    .S(_22600_),
    .Z(_03669_));
 BUF_X8 _53020_ (.A(_21301_),
    .Z(_22605_));
 BUF_X4 _53021_ (.A(_22598_),
    .Z(_22606_));
 MUX2_X1 _53022_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [741]),
    .B(_22605_),
    .S(_22606_),
    .Z(_03670_));
 MUX2_X1 _53023_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [742]),
    .B(_22529_),
    .S(_22606_),
    .Z(_03671_));
 MUX2_X1 _53024_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [743]),
    .B(_22337_),
    .S(_22606_),
    .Z(_03672_));
 MUX2_X1 _53025_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [744]),
    .B(_22503_),
    .S(_22606_),
    .Z(_03673_));
 MUX2_X1 _53026_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [745]),
    .B(_22582_),
    .S(_22606_),
    .Z(_03674_));
 NAND4_X1 _53027_ (.A1(_22399_),
    .A2(_21311_),
    .A3(_22589_),
    .A4(_22602_),
    .ZN(_22607_));
 INV_X1 _53028_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [746]),
    .ZN(_22608_));
 OAI21_X1 _53029_ (.A(_22607_),
    .B1(_22600_),
    .B2(_22608_),
    .ZN(_03675_));
 MUX2_X1 _53030_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [747]),
    .B(_22370_),
    .S(_22606_),
    .Z(_03676_));
 MUX2_X1 _53031_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [748]),
    .B(_22397_),
    .S(_22606_),
    .Z(_03677_));
 MUX2_X1 _53032_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [749]),
    .B(_22556_),
    .S(_22606_),
    .Z(_03678_));
 BUF_X8 _53033_ (.A(_08561_),
    .Z(_22609_));
 MUX2_X1 _53034_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [750]),
    .B(_22609_),
    .S(_22606_),
    .Z(_03680_));
 MUX2_X1 _53035_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [751]),
    .B(_22583_),
    .S(_22606_),
    .Z(_03681_));
 BUF_X16 _53036_ (.A(_22598_),
    .Z(_22610_));
 MUX2_X1 _53037_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [752]),
    .B(_22470_),
    .S(_22610_),
    .Z(_03682_));
 MUX2_X1 _53038_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [753]),
    .B(_22560_),
    .S(_22610_),
    .Z(_03683_));
 MUX2_X1 _53039_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [754]),
    .B(_22533_),
    .S(_22610_),
    .Z(_03684_));
 NAND4_X1 _53040_ (.A1(_22399_),
    .A2(_08578_),
    .A3(_22589_),
    .A4(_22602_),
    .ZN(_22611_));
 INV_X1 _53041_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [755]),
    .ZN(_22612_));
 OAI21_X1 _53042_ (.A(_22611_),
    .B1(_22600_),
    .B2(_22612_),
    .ZN(_03685_));
 BUF_X8 _53043_ (.A(_08581_),
    .Z(_22613_));
 MUX2_X1 _53044_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [756]),
    .B(_22613_),
    .S(_22610_),
    .Z(_03686_));
 MUX2_X1 _53045_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [757]),
    .B(_22561_),
    .S(_22610_),
    .Z(_03687_));
 MUX2_X1 _53046_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [758]),
    .B(_22511_),
    .S(_22610_),
    .Z(_03688_));
 MUX2_X1 _53047_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [759]),
    .B(_22512_),
    .S(_22610_),
    .Z(_03689_));
 BUF_X16 _53048_ (.A(_08594_),
    .Z(_22614_));
 MUX2_X1 _53049_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [760]),
    .B(_22614_),
    .S(_22610_),
    .Z(_03691_));
 MUX2_X1 _53050_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [761]),
    .B(_22426_),
    .S(_22610_),
    .Z(_03692_));
 BUF_X16 _53051_ (.A(_08600_),
    .Z(_22615_));
 MUX2_X1 _53052_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [762]),
    .B(_22615_),
    .S(_22610_),
    .Z(_03693_));
 BUF_X16 _53053_ (.A(_22598_),
    .Z(_22616_));
 MUX2_X1 _53054_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [763]),
    .B(_22248_),
    .S(_22616_),
    .Z(_03694_));
 MUX2_X1 _53055_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [764]),
    .B(_22479_),
    .S(_22616_),
    .Z(_03695_));
 BUF_X8 _53056_ (.A(_08611_),
    .Z(_22617_));
 MUX2_X1 _53057_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [765]),
    .B(_22617_),
    .S(_22616_),
    .Z(_03696_));
 NAND4_X1 _53058_ (.A1(_22399_),
    .A2(_08614_),
    .A3(_22589_),
    .A4(_22602_),
    .ZN(_22618_));
 INV_X2 _53059_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [766]),
    .ZN(_22619_));
 OAI21_X1 _53060_ (.A(_22618_),
    .B1(_22600_),
    .B2(_22619_),
    .ZN(_03697_));
 BUF_X4 _53061_ (.A(_08617_),
    .Z(_22620_));
 MUX2_X1 _53062_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [767]),
    .B(_22620_),
    .S(_22616_),
    .Z(_03698_));
 MUX2_X1 _53063_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [768]),
    .B(_22570_),
    .S(_22616_),
    .Z(_03699_));
 MUX2_X1 _53064_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [769]),
    .B(_22452_),
    .S(_22616_),
    .Z(_03700_));
 MUX2_X1 _53065_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [770]),
    .B(_22541_),
    .S(_22616_),
    .Z(_03702_));
 MUX2_X1 _53066_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [771]),
    .B(_22380_),
    .S(_22616_),
    .Z(_03703_));
 MUX2_X1 _53067_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [772]),
    .B(_22428_),
    .S(_22616_),
    .Z(_03704_));
 NAND4_X1 _53068_ (.A1(_22399_),
    .A2(_21591_),
    .A3(_22589_),
    .A4(_22602_),
    .ZN(_22621_));
 INV_X2 _53069_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [773]),
    .ZN(_22622_));
 OAI21_X1 _53070_ (.A(_22621_),
    .B1(_22600_),
    .B2(_22622_),
    .ZN(_03705_));
 MUX2_X1 _53071_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [774]),
    .B(_22329_),
    .S(_22616_),
    .Z(_03706_));
 MUX2_X1 _53072_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [775]),
    .B(_22596_),
    .S(_22599_),
    .Z(_03707_));
 MUX2_X1 _53073_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [776]),
    .B(_22516_),
    .S(_22599_),
    .Z(_03708_));
 MUX2_X1 _53074_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [777]),
    .B(_22573_),
    .S(_22599_),
    .Z(_03709_));
 MUX2_X1 _53075_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [778]),
    .B(_22492_),
    .S(_22599_),
    .Z(_03710_));
 MUX2_X1 _53076_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [779]),
    .B(_22493_),
    .S(_22599_),
    .Z(_03711_));
 MUX2_X1 _53077_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [780]),
    .B(_22455_),
    .S(_22599_),
    .Z(_03713_));
 MUX2_X1 _53078_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [781]),
    .B(_22456_),
    .S(_22599_),
    .Z(_03714_));
 MUX2_X1 _53079_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [782]),
    .B(_22517_),
    .S(_22599_),
    .Z(_03715_));
 MUX2_X1 _53080_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [783]),
    .B(_22494_),
    .S(_22599_),
    .Z(_03716_));
 AND2_X4 _53081_ (.A1(_11131_),
    .A2(_21574_),
    .ZN(_22623_));
 BUF_X8 _53082_ (.A(_22623_),
    .Z(_22624_));
 BUF_X8 _53083_ (.A(_22624_),
    .Z(_22625_));
 MUX2_X1 _53084_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [686]),
    .B(_22384_),
    .S(_22625_),
    .Z(_03608_));
 MUX2_X1 _53085_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [687]),
    .B(_22358_),
    .S(_22625_),
    .Z(_03609_));
 MUX2_X1 _53086_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [688]),
    .B(_22601_),
    .S(_22625_),
    .Z(_03610_));
 BUF_X8 _53087_ (.A(_21608_),
    .Z(_22626_));
 MUX2_X1 _53088_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [689]),
    .B(_22626_),
    .S(_22625_),
    .Z(_03611_));
 MUX2_X1 _53089_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [690]),
    .B(_22316_),
    .S(_22625_),
    .Z(_03613_));
 NAND4_X1 _53090_ (.A1(_22422_),
    .A2(_21299_),
    .A3(_22589_),
    .A4(_22602_),
    .ZN(_22627_));
 INV_X1 _53091_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [691]),
    .ZN(_22628_));
 OAI21_X1 _53092_ (.A(_22627_),
    .B1(_22625_),
    .B2(_22628_),
    .ZN(_03614_));
 MUX2_X1 _53093_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [692]),
    .B(_22605_),
    .S(_22625_),
    .Z(_03615_));
 BUF_X8 _53094_ (.A(_22623_),
    .Z(_22629_));
 MUX2_X1 _53095_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [693]),
    .B(_22529_),
    .S(_22629_),
    .Z(_03616_));
 MUX2_X1 _53096_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [694]),
    .B(_22337_),
    .S(_22629_),
    .Z(_03617_));
 MUX2_X1 _53097_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [695]),
    .B(_22503_),
    .S(_22629_),
    .Z(_03618_));
 MUX2_X1 _53098_ (.A(net1392),
    .B(_22582_),
    .S(_22629_),
    .Z(_03619_));
 MUX2_X1 _53099_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [697]),
    .B(_22504_),
    .S(_22629_),
    .Z(_03620_));
 BUF_X8 _53100_ (.A(_08551_),
    .Z(_22630_));
 MUX2_X1 _53101_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [698]),
    .B(_22630_),
    .S(_22629_),
    .Z(_03621_));
 MUX2_X1 _53102_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [699]),
    .B(_22397_),
    .S(_22629_),
    .Z(_03622_));
 MUX2_X1 _53103_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [700]),
    .B(_22556_),
    .S(_22629_),
    .Z(_03625_));
 MUX2_X1 _53104_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [701]),
    .B(_22609_),
    .S(_22629_),
    .Z(_03626_));
 NAND4_X1 _53105_ (.A1(_22422_),
    .A2(_22371_),
    .A3(_22589_),
    .A4(_22602_),
    .ZN(_22631_));
 INV_X1 _53106_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [702]),
    .ZN(_22632_));
 OAI21_X1 _53107_ (.A(_22631_),
    .B1(_22625_),
    .B2(_22632_),
    .ZN(_03627_));
 MUX2_X1 _53108_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [703]),
    .B(_22470_),
    .S(_22629_),
    .Z(_03628_));
 BUF_X16 _53109_ (.A(_22623_),
    .Z(_22633_));
 MUX2_X1 _53110_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [704]),
    .B(_22560_),
    .S(_22633_),
    .Z(_03629_));
 MUX2_X1 _53111_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [705]),
    .B(_22533_),
    .S(_22633_),
    .Z(_03630_));
 MUX2_X1 _53112_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [706]),
    .B(_22471_),
    .S(_22633_),
    .Z(_03631_));
 MUX2_X1 _53113_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [707]),
    .B(_22613_),
    .S(_22633_),
    .Z(_03632_));
 MUX2_X1 _53114_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [708]),
    .B(_22561_),
    .S(_22633_),
    .Z(_03633_));
 MUX2_X1 _53115_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [709]),
    .B(_22511_),
    .S(_22633_),
    .Z(_03634_));
 MUX2_X1 _53116_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [710]),
    .B(_22512_),
    .S(_22633_),
    .Z(_03636_));
 MUX2_X1 _53117_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [711]),
    .B(_22614_),
    .S(_22633_),
    .Z(_03637_));
 MUX2_X1 _53118_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [712]),
    .B(_22426_),
    .S(_22633_),
    .Z(_03638_));
 MUX2_X1 _53119_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [713]),
    .B(_22615_),
    .S(_22633_),
    .Z(_03639_));
 BUF_X4 _53120_ (.A(_22360_),
    .Z(_22634_));
 NAND4_X1 _53121_ (.A1(_22422_),
    .A2(_21725_),
    .A3(_22634_),
    .A4(_22602_),
    .ZN(_22635_));
 INV_X1 _53122_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [714]),
    .ZN(_22636_));
 OAI21_X1 _53123_ (.A(_22635_),
    .B1(_22625_),
    .B2(_22636_),
    .ZN(_03640_));
 BUF_X16 _53124_ (.A(_22623_),
    .Z(_22637_));
 MUX2_X1 _53125_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [715]),
    .B(_22479_),
    .S(_22637_),
    .Z(_03641_));
 MUX2_X1 _53126_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [716]),
    .B(_22617_),
    .S(_22637_),
    .Z(_03642_));
 BUF_X4 _53127_ (.A(_08614_),
    .Z(_22638_));
 MUX2_X1 _53128_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [717]),
    .B(_22638_),
    .S(_22637_),
    .Z(_03643_));
 MUX2_X1 _53129_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [718]),
    .B(_22620_),
    .S(_22637_),
    .Z(_03644_));
 MUX2_X1 _53130_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [719]),
    .B(_22570_),
    .S(_22637_),
    .Z(_03645_));
 MUX2_X1 _53131_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [720]),
    .B(_22452_),
    .S(_22637_),
    .Z(_03647_));
 MUX2_X1 _53132_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [721]),
    .B(_22541_),
    .S(_22637_),
    .Z(_03648_));
 MUX2_X1 _53133_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [722]),
    .B(_22380_),
    .S(_22637_),
    .Z(_03649_));
 NAND4_X1 _53134_ (.A1(_22422_),
    .A2(_21330_),
    .A3(_22634_),
    .A4(_22602_),
    .ZN(_22639_));
 INV_X1 _53135_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [723]),
    .ZN(_22640_));
 OAI21_X1 _53136_ (.A(_22639_),
    .B1(_22625_),
    .B2(_22640_),
    .ZN(_03650_));
 MUX2_X1 _53137_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [724]),
    .B(_22542_),
    .S(_22637_),
    .Z(_03651_));
 BUF_X8 _53138_ (.A(_21339_),
    .Z(_22641_));
 MUX2_X1 _53139_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [725]),
    .B(_22641_),
    .S(_22637_),
    .Z(_03652_));
 MUX2_X1 _53140_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [726]),
    .B(_22596_),
    .S(_22624_),
    .Z(_03653_));
 MUX2_X1 _53141_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [727]),
    .B(_22516_),
    .S(_22624_),
    .Z(_03654_));
 MUX2_X1 _53142_ (.A(net1391),
    .B(_22573_),
    .S(_22624_),
    .Z(_03655_));
 MUX2_X1 _53143_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [729]),
    .B(_22492_),
    .S(_22624_),
    .Z(_03656_));
 MUX2_X1 _53144_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [730]),
    .B(_22493_),
    .S(_22624_),
    .Z(_03658_));
 MUX2_X1 _53145_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [731]),
    .B(_22455_),
    .S(_22624_),
    .Z(_03659_));
 MUX2_X1 _53146_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [732]),
    .B(_22456_),
    .S(_22624_),
    .Z(_03660_));
 MUX2_X1 _53147_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [733]),
    .B(_22517_),
    .S(_22624_),
    .Z(_03661_));
 MUX2_X1 _53148_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [734]),
    .B(_22494_),
    .S(_22624_),
    .Z(_03662_));
 BUF_X16 _53149_ (.A(_11136_),
    .Z(_22642_));
 AND2_X4 _53150_ (.A1(_22642_),
    .A2(_21679_),
    .ZN(_22643_));
 BUF_X16 _53151_ (.A(_22643_),
    .Z(_22644_));
 BUF_X8 _53152_ (.A(_22644_),
    .Z(_22645_));
 MUX2_X1 _53153_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [637]),
    .B(_22384_),
    .S(_22645_),
    .Z(_03554_));
 MUX2_X1 _53154_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [638]),
    .B(_22358_),
    .S(_22645_),
    .Z(_03555_));
 BUF_X4 _53155_ (.A(_11127_),
    .Z(_22646_));
 NAND4_X1 _53156_ (.A1(_22243_),
    .A2(_21383_),
    .A3(_22634_),
    .A4(_22646_),
    .ZN(_22647_));
 INV_X1 _53157_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [639]),
    .ZN(_22648_));
 OAI21_X1 _53158_ (.A(_22647_),
    .B1(_22645_),
    .B2(_22648_),
    .ZN(_03556_));
 MUX2_X1 _53159_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [640]),
    .B(_22626_),
    .S(_22645_),
    .Z(_03558_));
 MUX2_X1 _53160_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [641]),
    .B(_22316_),
    .S(_22645_),
    .Z(_03559_));
 BUF_X8 _53161_ (.A(_22643_),
    .Z(_22649_));
 MUX2_X1 _53162_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [642]),
    .B(_22392_),
    .S(_22649_),
    .Z(_03560_));
 MUX2_X1 _53163_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [643]),
    .B(_22605_),
    .S(_22649_),
    .Z(_03561_));
 MUX2_X1 _53164_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [644]),
    .B(_22529_),
    .S(_22649_),
    .Z(_03562_));
 MUX2_X1 _53165_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [645]),
    .B(_22337_),
    .S(_22649_),
    .Z(_03563_));
 MUX2_X1 _53166_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [646]),
    .B(_22503_),
    .S(_22649_),
    .Z(_03564_));
 MUX2_X1 _53167_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [647]),
    .B(_22582_),
    .S(_22649_),
    .Z(_03565_));
 MUX2_X1 _53168_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [648]),
    .B(_22504_),
    .S(_22649_),
    .Z(_03566_));
 MUX2_X1 _53169_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [649]),
    .B(_22630_),
    .S(_22649_),
    .Z(_03567_));
 BUF_X8 _53170_ (.A(_08555_),
    .Z(_22650_));
 MUX2_X1 _53171_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [650]),
    .B(_22650_),
    .S(_22649_),
    .Z(_03569_));
 MUX2_X1 _53172_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [651]),
    .B(_22556_),
    .S(_22649_),
    .Z(_03570_));
 BUF_X16 _53173_ (.A(_22643_),
    .Z(_22651_));
 MUX2_X1 _53174_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [652]),
    .B(_22609_),
    .S(_22651_),
    .Z(_03571_));
 MUX2_X1 _53175_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [653]),
    .B(_22583_),
    .S(_22651_),
    .Z(_03572_));
 MUX2_X1 _53176_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [654]),
    .B(_22470_),
    .S(_22651_),
    .Z(_03573_));
 MUX2_X1 _53177_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [655]),
    .B(_22560_),
    .S(_22651_),
    .Z(_03574_));
 MUX2_X1 _53178_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [656]),
    .B(_22533_),
    .S(_22651_),
    .Z(_03575_));
 MUX2_X1 _53179_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [657]),
    .B(_22471_),
    .S(_22651_),
    .Z(_03576_));
 MUX2_X1 _53180_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [658]),
    .B(_22613_),
    .S(_22651_),
    .Z(_03577_));
 NAND4_X1 _53181_ (.A1(_22243_),
    .A2(_10579_),
    .A3(_22634_),
    .A4(_22646_),
    .ZN(_22652_));
 INV_X4 _53182_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [659]),
    .ZN(_22653_));
 OAI21_X1 _53183_ (.A(_22652_),
    .B1(_22645_),
    .B2(_22653_),
    .ZN(_03578_));
 MUX2_X1 _53184_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [660]),
    .B(_22511_),
    .S(_22651_),
    .Z(_03580_));
 MUX2_X1 _53185_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [661]),
    .B(_22512_),
    .S(_22651_),
    .Z(_03581_));
 MUX2_X1 _53186_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [662]),
    .B(_22614_),
    .S(_22651_),
    .Z(_03582_));
 BUF_X16 _53187_ (.A(_22643_),
    .Z(_22654_));
 MUX2_X1 _53188_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [663]),
    .B(_22426_),
    .S(_22654_),
    .Z(_03583_));
 MUX2_X1 _53189_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [664]),
    .B(_22615_),
    .S(_22654_),
    .Z(_03584_));
 NAND4_X1 _53190_ (.A1(_10832_),
    .A2(_08604_),
    .A3(_22634_),
    .A4(_22646_),
    .ZN(_22655_));
 INV_X1 _53191_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [665]),
    .ZN(_22656_));
 OAI21_X1 _53192_ (.A(_22655_),
    .B1(_22645_),
    .B2(_22656_),
    .ZN(_03585_));
 NAND4_X1 _53193_ (.A1(_10832_),
    .A2(_08608_),
    .A3(_22634_),
    .A4(_22646_),
    .ZN(_22657_));
 INV_X1 _53194_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [666]),
    .ZN(_22658_));
 OAI21_X1 _53195_ (.A(_22657_),
    .B1(_22645_),
    .B2(_22658_),
    .ZN(_03586_));
 MUX2_X1 _53196_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [667]),
    .B(_22617_),
    .S(_22654_),
    .Z(_03587_));
 MUX2_X1 _53197_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [668]),
    .B(_22638_),
    .S(_22654_),
    .Z(_03588_));
 MUX2_X1 _53198_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [669]),
    .B(_22620_),
    .S(_22654_),
    .Z(_03589_));
 MUX2_X1 _53199_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [670]),
    .B(_22570_),
    .S(_22654_),
    .Z(_03591_));
 MUX2_X1 _53200_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [671]),
    .B(_22452_),
    .S(_22654_),
    .Z(_03592_));
 MUX2_X1 _53201_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [672]),
    .B(_22541_),
    .S(_22654_),
    .Z(_03593_));
 BUF_X8 _53202_ (.A(_08629_),
    .Z(_22659_));
 MUX2_X1 _53203_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [673]),
    .B(_22659_),
    .S(_22654_),
    .Z(_03594_));
 NAND4_X1 _53204_ (.A1(_10832_),
    .A2(_21330_),
    .A3(_22634_),
    .A4(_22646_),
    .ZN(_22660_));
 INV_X2 _53205_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [674]),
    .ZN(_22661_));
 OAI21_X1 _53206_ (.A(_22660_),
    .B1(_22645_),
    .B2(_22661_),
    .ZN(_03595_));
 MUX2_X1 _53207_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [675]),
    .B(_22542_),
    .S(_22654_),
    .Z(_03596_));
 MUX2_X1 _53208_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [676]),
    .B(_22641_),
    .S(_22644_),
    .Z(_03597_));
 MUX2_X1 _53209_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [677]),
    .B(_22596_),
    .S(_22644_),
    .Z(_03598_));
 MUX2_X1 _53210_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [678]),
    .B(_22516_),
    .S(_22644_),
    .Z(_03599_));
 MUX2_X1 _53211_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [679]),
    .B(_22573_),
    .S(_22644_),
    .Z(_03600_));
 MUX2_X1 _53212_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [680]),
    .B(_22492_),
    .S(_22644_),
    .Z(_03602_));
 MUX2_X1 _53213_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [681]),
    .B(_22493_),
    .S(_22644_),
    .Z(_03603_));
 MUX2_X1 _53214_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [682]),
    .B(_22455_),
    .S(_22644_),
    .Z(_03604_));
 MUX2_X1 _53215_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [683]),
    .B(_22456_),
    .S(_22644_),
    .Z(_03605_));
 MUX2_X1 _53216_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [684]),
    .B(_22517_),
    .S(_22644_),
    .Z(_03606_));
 NAND4_X1 _53217_ (.A1(_10832_),
    .A2(_22381_),
    .A3(_11128_),
    .A4(_21377_),
    .ZN(_22662_));
 INV_X1 _53218_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [685]),
    .ZN(_22663_));
 OAI21_X1 _53219_ (.A(_22662_),
    .B1(_22645_),
    .B2(_22663_),
    .ZN(_03607_));
 AND2_X4 _53220_ (.A1(_11141_),
    .A2(_21412_),
    .ZN(_22664_));
 BUF_X8 _53221_ (.A(_22664_),
    .Z(_22665_));
 BUF_X8 _53222_ (.A(_22665_),
    .Z(_22666_));
 MUX2_X1 _53223_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [588]),
    .B(_22384_),
    .S(_22666_),
    .Z(_03499_));
 BUF_X4 _53224_ (.A(_21605_),
    .Z(_22667_));
 MUX2_X1 _53225_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [589]),
    .B(_22667_),
    .S(_22666_),
    .Z(_03500_));
 MUX2_X1 _53226_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [590]),
    .B(_22601_),
    .S(_22666_),
    .Z(_03502_));
 MUX2_X1 _53227_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [591]),
    .B(_22626_),
    .S(_22666_),
    .Z(_03503_));
 NAND4_X1 _53228_ (.A1(_22480_),
    .A2(_21297_),
    .A3(_22634_),
    .A4(_22646_),
    .ZN(_22668_));
 INV_X1 _53229_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [592]),
    .ZN(_22669_));
 OAI21_X1 _53230_ (.A(_22668_),
    .B1(_22666_),
    .B2(_22669_),
    .ZN(_03504_));
 BUF_X8 _53231_ (.A(_21299_),
    .Z(_22670_));
 MUX2_X1 _53232_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [593]),
    .B(_22670_),
    .S(_22666_),
    .Z(_03505_));
 BUF_X8 _53233_ (.A(_22664_),
    .Z(_22671_));
 MUX2_X1 _53234_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [594]),
    .B(_22605_),
    .S(_22671_),
    .Z(_03506_));
 MUX2_X1 _53235_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [595]),
    .B(_22529_),
    .S(_22671_),
    .Z(_03507_));
 MUX2_X1 _53236_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [596]),
    .B(_22337_),
    .S(_22671_),
    .Z(_03508_));
 MUX2_X1 _53237_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [597]),
    .B(_22503_),
    .S(_22671_),
    .Z(_03509_));
 MUX2_X1 _53238_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [598]),
    .B(_22582_),
    .S(_22671_),
    .Z(_03510_));
 NAND4_X1 _53239_ (.A1(_22480_),
    .A2(_21311_),
    .A3(_22634_),
    .A4(_22646_),
    .ZN(_22672_));
 INV_X1 _53240_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [599]),
    .ZN(_22673_));
 OAI21_X1 _53241_ (.A(_22672_),
    .B1(_22666_),
    .B2(_22673_),
    .ZN(_03511_));
 MUX2_X1 _53242_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [600]),
    .B(_22630_),
    .S(_22671_),
    .Z(_03514_));
 MUX2_X1 _53243_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [601]),
    .B(_22650_),
    .S(_22671_),
    .Z(_03515_));
 MUX2_X1 _53244_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [602]),
    .B(_22556_),
    .S(_22671_),
    .Z(_03516_));
 MUX2_X1 _53245_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [603]),
    .B(_22609_),
    .S(_22671_),
    .Z(_03517_));
 MUX2_X1 _53246_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [604]),
    .B(_22583_),
    .S(_22671_),
    .Z(_03518_));
 BUF_X16 _53247_ (.A(_22664_),
    .Z(_22674_));
 MUX2_X1 _53248_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [605]),
    .B(_22470_),
    .S(_22674_),
    .Z(_03519_));
 MUX2_X1 _53249_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [606]),
    .B(_22560_),
    .S(_22674_),
    .Z(_03520_));
 MUX2_X1 _53250_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [607]),
    .B(_22533_),
    .S(_22674_),
    .Z(_03521_));
 NAND4_X1 _53251_ (.A1(_22480_),
    .A2(_08578_),
    .A3(_22634_),
    .A4(_22646_),
    .ZN(_22675_));
 INV_X1 _53252_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [608]),
    .ZN(_22676_));
 OAI21_X1 _53253_ (.A(_22675_),
    .B1(_22666_),
    .B2(_22676_),
    .ZN(_03522_));
 MUX2_X1 _53254_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [609]),
    .B(_22613_),
    .S(_22674_),
    .Z(_03523_));
 MUX2_X1 _53255_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [610]),
    .B(_22561_),
    .S(_22674_),
    .Z(_03525_));
 MUX2_X1 _53256_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [611]),
    .B(_22511_),
    .S(_22674_),
    .Z(_03526_));
 BUF_X4 _53257_ (.A(_22360_),
    .Z(_22677_));
 NAND4_X1 _53258_ (.A1(_22480_),
    .A2(_22025_),
    .A3(_22677_),
    .A4(_22646_),
    .ZN(_22678_));
 INV_X1 _53259_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [612]),
    .ZN(_22679_));
 OAI21_X1 _53260_ (.A(_22678_),
    .B1(_22666_),
    .B2(_22679_),
    .ZN(_03527_));
 MUX2_X1 _53261_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [613]),
    .B(_22614_),
    .S(_22674_),
    .Z(_03528_));
 BUF_X8 _53262_ (.A(_08597_),
    .Z(_22680_));
 MUX2_X1 _53263_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [614]),
    .B(_22680_),
    .S(_22674_),
    .Z(_03529_));
 MUX2_X1 _53264_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [615]),
    .B(_22615_),
    .S(_22674_),
    .Z(_03530_));
 BUF_X8 _53265_ (.A(_08604_),
    .Z(_22681_));
 MUX2_X1 _53266_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [616]),
    .B(_22681_),
    .S(_22674_),
    .Z(_03531_));
 BUF_X16 _53267_ (.A(_22664_),
    .Z(_22682_));
 MUX2_X1 _53268_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [617]),
    .B(_22479_),
    .S(_22682_),
    .Z(_03532_));
 MUX2_X1 _53269_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [618]),
    .B(_22617_),
    .S(_22682_),
    .Z(_03533_));
 MUX2_X1 _53270_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [619]),
    .B(_22638_),
    .S(_22682_),
    .Z(_03534_));
 MUX2_X1 _53271_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [620]),
    .B(_22620_),
    .S(_22682_),
    .Z(_03536_));
 MUX2_X1 _53272_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [621]),
    .B(_22570_),
    .S(_22682_),
    .Z(_03537_));
 MUX2_X1 _53273_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [622]),
    .B(_22452_),
    .S(_22682_),
    .Z(_03538_));
 MUX2_X1 _53274_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [623]),
    .B(_22541_),
    .S(_22682_),
    .Z(_03539_));
 MUX2_X1 _53275_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [624]),
    .B(_22659_),
    .S(_22682_),
    .Z(_03540_));
 NAND4_X1 _53276_ (.A1(_22480_),
    .A2(_21330_),
    .A3(_22677_),
    .A4(_22646_),
    .ZN(_22683_));
 INV_X1 _53277_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [625]),
    .ZN(_22684_));
 OAI21_X1 _53278_ (.A(_22683_),
    .B1(_22666_),
    .B2(_22684_),
    .ZN(_03541_));
 MUX2_X1 _53279_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [626]),
    .B(_22542_),
    .S(_22682_),
    .Z(_03542_));
 MUX2_X1 _53280_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [627]),
    .B(_22641_),
    .S(_22682_),
    .Z(_03543_));
 MUX2_X1 _53281_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [628]),
    .B(_22596_),
    .S(_22665_),
    .Z(_03544_));
 MUX2_X1 _53282_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [629]),
    .B(_22516_),
    .S(_22665_),
    .Z(_03545_));
 MUX2_X1 _53283_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [630]),
    .B(_22573_),
    .S(_22665_),
    .Z(_03547_));
 MUX2_X1 _53284_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [631]),
    .B(_22492_),
    .S(_22665_),
    .Z(_03548_));
 MUX2_X1 _53285_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [632]),
    .B(_22493_),
    .S(_22665_),
    .Z(_03549_));
 MUX2_X1 _53286_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [633]),
    .B(_22455_),
    .S(_22665_),
    .Z(_03550_));
 MUX2_X1 _53287_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [634]),
    .B(_22456_),
    .S(_22665_),
    .Z(_03551_));
 MUX2_X1 _53288_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [635]),
    .B(_22517_),
    .S(_22665_),
    .Z(_03552_));
 MUX2_X1 _53289_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [636]),
    .B(_22494_),
    .S(_22665_),
    .Z(_03553_));
 BUF_X4 _53290_ (.A(_21598_),
    .Z(_22685_));
 AND2_X4 _53291_ (.A1(_11146_),
    .A2(_21432_),
    .ZN(_22686_));
 BUF_X16 _53292_ (.A(_22686_),
    .Z(_22687_));
 BUF_X8 _53293_ (.A(_22687_),
    .Z(_22688_));
 MUX2_X1 _53294_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [539]),
    .B(_22685_),
    .S(_22688_),
    .Z(_03445_));
 MUX2_X1 _53295_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [540]),
    .B(_22667_),
    .S(_22688_),
    .Z(_03447_));
 MUX2_X1 _53296_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [541]),
    .B(_22601_),
    .S(_22688_),
    .Z(_03448_));
 MUX2_X1 _53297_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [542]),
    .B(_22626_),
    .S(_22688_),
    .Z(_03449_));
 MUX2_X1 _53298_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [543]),
    .B(_22316_),
    .S(_22688_),
    .Z(_03450_));
 MUX2_X1 _53299_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [544]),
    .B(_22670_),
    .S(_22688_),
    .Z(_03451_));
 MUX2_X1 _53300_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [545]),
    .B(_22605_),
    .S(_22688_),
    .Z(_03452_));
 MUX2_X1 _53301_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [546]),
    .B(_22529_),
    .S(_22688_),
    .Z(_03453_));
 BUF_X8 _53302_ (.A(_22686_),
    .Z(_22689_));
 MUX2_X1 _53303_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [547]),
    .B(_22337_),
    .S(_22689_),
    .Z(_03454_));
 MUX2_X1 _53304_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [548]),
    .B(_22503_),
    .S(_22689_),
    .Z(_03455_));
 MUX2_X1 _53305_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [549]),
    .B(_22582_),
    .S(_22689_),
    .Z(_03456_));
 MUX2_X1 _53306_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [550]),
    .B(_22504_),
    .S(_22689_),
    .Z(_03458_));
 MUX2_X1 _53307_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [551]),
    .B(_22630_),
    .S(_22689_),
    .Z(_03459_));
 MUX2_X1 _53308_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [552]),
    .B(_22650_),
    .S(_22689_),
    .Z(_03460_));
 MUX2_X1 _53309_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [553]),
    .B(_22556_),
    .S(_22689_),
    .Z(_03461_));
 MUX2_X1 _53310_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [554]),
    .B(_22609_),
    .S(_22689_),
    .Z(_03462_));
 MUX2_X1 _53311_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [555]),
    .B(_22583_),
    .S(_22689_),
    .Z(_03463_));
 MUX2_X1 _53312_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [556]),
    .B(_22470_),
    .S(_22689_),
    .Z(_03464_));
 BUF_X16 _53313_ (.A(_22686_),
    .Z(_22690_));
 MUX2_X1 _53314_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [557]),
    .B(_22560_),
    .S(_22690_),
    .Z(_03465_));
 MUX2_X1 _53315_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [558]),
    .B(_22533_),
    .S(_22690_),
    .Z(_03466_));
 MUX2_X1 _53316_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [559]),
    .B(_22471_),
    .S(_22690_),
    .Z(_03467_));
 BUF_X4 _53317_ (.A(_11127_),
    .Z(_22691_));
 NAND4_X1 _53318_ (.A1(_22498_),
    .A2(_08581_),
    .A3(_22677_),
    .A4(_22691_),
    .ZN(_22692_));
 INV_X1 _53319_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [560]),
    .ZN(_22693_));
 OAI21_X1 _53320_ (.A(_22692_),
    .B1(_22688_),
    .B2(_22693_),
    .ZN(_03469_));
 MUX2_X1 _53321_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [561]),
    .B(_22561_),
    .S(_22690_),
    .Z(_03470_));
 MUX2_X1 _53322_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [562]),
    .B(_22511_),
    .S(_22690_),
    .Z(_03471_));
 MUX2_X1 _53323_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [563]),
    .B(_22512_),
    .S(_22690_),
    .Z(_03472_));
 MUX2_X1 _53324_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [564]),
    .B(_22614_),
    .S(_22690_),
    .Z(_03473_));
 MUX2_X1 _53325_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [565]),
    .B(_22680_),
    .S(_22690_),
    .Z(_03474_));
 MUX2_X1 _53326_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [566]),
    .B(_22615_),
    .S(_22690_),
    .Z(_03475_));
 MUX2_X1 _53327_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [567]),
    .B(_22681_),
    .S(_22690_),
    .Z(_03476_));
 BUF_X16 _53328_ (.A(_22686_),
    .Z(_22694_));
 MUX2_X1 _53329_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [568]),
    .B(_22479_),
    .S(_22694_),
    .Z(_03477_));
 MUX2_X1 _53330_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [569]),
    .B(_22617_),
    .S(_22694_),
    .Z(_03478_));
 MUX2_X1 _53331_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [570]),
    .B(_22638_),
    .S(_22694_),
    .Z(_03480_));
 MUX2_X1 _53332_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [571]),
    .B(_22620_),
    .S(_22694_),
    .Z(_03481_));
 MUX2_X1 _53333_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [572]),
    .B(_22570_),
    .S(_22694_),
    .Z(_03482_));
 MUX2_X1 _53334_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [573]),
    .B(_22452_),
    .S(_22694_),
    .Z(_03483_));
 MUX2_X1 _53335_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [574]),
    .B(_22541_),
    .S(_22694_),
    .Z(_03484_));
 MUX2_X1 _53336_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [575]),
    .B(_22659_),
    .S(_22694_),
    .Z(_03485_));
 MUX2_X1 _53337_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [576]),
    .B(_22428_),
    .S(_22694_),
    .Z(_03486_));
 MUX2_X1 _53338_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [577]),
    .B(_22542_),
    .S(_22694_),
    .Z(_03487_));
 MUX2_X1 _53339_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [578]),
    .B(_22641_),
    .S(_22687_),
    .Z(_03488_));
 MUX2_X1 _53340_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [579]),
    .B(_22596_),
    .S(_22687_),
    .Z(_03489_));
 MUX2_X1 _53341_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [580]),
    .B(_22516_),
    .S(_22687_),
    .Z(_03491_));
 MUX2_X1 _53342_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [581]),
    .B(_22573_),
    .S(_22687_),
    .Z(_03492_));
 NAND4_X1 _53343_ (.A1(_22498_),
    .A2(_22381_),
    .A3(_11128_),
    .A4(_21738_),
    .ZN(_22695_));
 INV_X1 _53344_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [582]),
    .ZN(_22696_));
 OAI21_X1 _53345_ (.A(_22695_),
    .B1(_22688_),
    .B2(_22696_),
    .ZN(_03493_));
 MUX2_X1 _53346_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [583]),
    .B(_22493_),
    .S(_22687_),
    .Z(_03494_));
 BUF_X4 _53347_ (.A(_21365_),
    .Z(_22697_));
 MUX2_X1 _53348_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [584]),
    .B(_22697_),
    .S(_22687_),
    .Z(_03495_));
 BUF_X8 _53349_ (.A(_21369_),
    .Z(_22698_));
 MUX2_X1 _53350_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [585]),
    .B(_22698_),
    .S(_22687_),
    .Z(_03496_));
 MUX2_X1 _53351_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [586]),
    .B(_22517_),
    .S(_22687_),
    .Z(_03497_));
 MUX2_X1 _53352_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [587]),
    .B(_22494_),
    .S(_22687_),
    .Z(_03498_));
 AND2_X4 _53353_ (.A1(_11152_),
    .A2(_21679_),
    .ZN(_22699_));
 BUF_X16 _53354_ (.A(_22699_),
    .Z(_22700_));
 BUF_X8 _53355_ (.A(_22700_),
    .Z(_22701_));
 MUX2_X1 _53356_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [490]),
    .B(_22685_),
    .S(_22701_),
    .Z(_03391_));
 MUX2_X1 _53357_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [491]),
    .B(_22667_),
    .S(_22701_),
    .Z(_03392_));
 MUX2_X1 _53358_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [492]),
    .B(_22601_),
    .S(_22701_),
    .Z(_03393_));
 NAND4_X1 _53359_ (.A1(_22525_),
    .A2(_21608_),
    .A3(_22677_),
    .A4(_22691_),
    .ZN(_22702_));
 INV_X1 _53360_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [493]),
    .ZN(_22703_));
 OAI21_X1 _53361_ (.A(_22702_),
    .B1(_22701_),
    .B2(_22703_),
    .ZN(_03394_));
 BUF_X16 _53362_ (.A(_22699_),
    .Z(_22704_));
 MUX2_X1 _53363_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [494]),
    .B(_21387_),
    .S(_22704_),
    .Z(_03395_));
 MUX2_X1 _53364_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [495]),
    .B(_22670_),
    .S(_22704_),
    .Z(_03396_));
 MUX2_X1 _53365_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [496]),
    .B(_22605_),
    .S(_22704_),
    .Z(_03397_));
 MUX2_X1 _53366_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [497]),
    .B(_22529_),
    .S(_22704_),
    .Z(_03398_));
 BUF_X8 _53367_ (.A(_21305_),
    .Z(_22705_));
 MUX2_X1 _53368_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [498]),
    .B(_22705_),
    .S(_22704_),
    .Z(_03399_));
 MUX2_X1 _53369_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [499]),
    .B(_22503_),
    .S(_22704_),
    .Z(_03400_));
 MUX2_X1 _53370_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [500]),
    .B(_22582_),
    .S(_22704_),
    .Z(_03403_));
 MUX2_X1 _53371_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [501]),
    .B(_22504_),
    .S(_22704_),
    .Z(_03404_));
 NAND4_X1 _53372_ (.A1(_22525_),
    .A2(_10563_),
    .A3(_22677_),
    .A4(_22691_),
    .ZN(_22706_));
 INV_X2 _53373_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [502]),
    .ZN(_22707_));
 OAI21_X1 _53374_ (.A(_22706_),
    .B1(_22701_),
    .B2(_22707_),
    .ZN(_03405_));
 MUX2_X1 _53375_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [503]),
    .B(_22650_),
    .S(_22704_),
    .Z(_03406_));
 MUX2_X1 _53376_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [504]),
    .B(_22556_),
    .S(_22704_),
    .Z(_03407_));
 BUF_X16 _53377_ (.A(_22699_),
    .Z(_22708_));
 MUX2_X1 _53378_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [505]),
    .B(_22609_),
    .S(_22708_),
    .Z(_03408_));
 MUX2_X1 _53379_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [506]),
    .B(_22583_),
    .S(_22708_),
    .Z(_03409_));
 MUX2_X1 _53380_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [507]),
    .B(_10573_),
    .S(_22708_),
    .Z(_03410_));
 MUX2_X1 _53381_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [508]),
    .B(_22560_),
    .S(_22708_),
    .Z(_03411_));
 MUX2_X1 _53382_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [509]),
    .B(_22533_),
    .S(_22708_),
    .Z(_03412_));
 MUX2_X1 _53383_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [510]),
    .B(_22471_),
    .S(_22708_),
    .Z(_03414_));
 NAND4_X1 _53384_ (.A1(_22525_),
    .A2(_08581_),
    .A3(_22677_),
    .A4(_22691_),
    .ZN(_22709_));
 INV_X1 _53385_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [511]),
    .ZN(_22710_));
 OAI21_X1 _53386_ (.A(_22709_),
    .B1(_22701_),
    .B2(_22710_),
    .ZN(_03415_));
 NAND4_X1 _53387_ (.A1(_22525_),
    .A2(_10579_),
    .A3(_22677_),
    .A4(_22691_),
    .ZN(_22711_));
 INV_X4 _53388_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [512]),
    .ZN(_22712_));
 OAI21_X1 _53389_ (.A(_22711_),
    .B1(_22701_),
    .B2(_22712_),
    .ZN(_03416_));
 MUX2_X1 _53390_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [513]),
    .B(_22511_),
    .S(_22708_),
    .Z(_03417_));
 MUX2_X1 _53391_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [514]),
    .B(_22512_),
    .S(_22708_),
    .Z(_03418_));
 MUX2_X1 _53392_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [515]),
    .B(_22614_),
    .S(_22708_),
    .Z(_03419_));
 MUX2_X1 _53393_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [516]),
    .B(_22680_),
    .S(_22708_),
    .Z(_03420_));
 BUF_X16 _53394_ (.A(_22699_),
    .Z(_22713_));
 MUX2_X1 _53395_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [517]),
    .B(_22615_),
    .S(_22713_),
    .Z(_03421_));
 MUX2_X1 _53396_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [518]),
    .B(_22681_),
    .S(_22713_),
    .Z(_03422_));
 MUX2_X1 _53397_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [519]),
    .B(_22479_),
    .S(_22713_),
    .Z(_03423_));
 MUX2_X1 _53398_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [520]),
    .B(_22617_),
    .S(_22713_),
    .Z(_03425_));
 MUX2_X1 _53399_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [521]),
    .B(_22638_),
    .S(_22713_),
    .Z(_03426_));
 MUX2_X1 _53400_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [522]),
    .B(_22620_),
    .S(_22713_),
    .Z(_03427_));
 MUX2_X1 _53401_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [523]),
    .B(_22570_),
    .S(_22713_),
    .Z(_03428_));
 NAND4_X2 _53402_ (.A1(_22525_),
    .A2(_21562_),
    .A3(_22677_),
    .A4(_22691_),
    .ZN(_22714_));
 INV_X1 _53403_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [524]),
    .ZN(_22715_));
 OAI21_X1 _53404_ (.A(_22714_),
    .B1(_22701_),
    .B2(_22715_),
    .ZN(_03429_));
 BUF_X8 _53405_ (.A(_22524_),
    .Z(_22716_));
 NAND4_X2 _53406_ (.A1(_22716_),
    .A2(_08626_),
    .A3(_22677_),
    .A4(_22691_),
    .ZN(_22717_));
 INV_X1 _53407_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [525]),
    .ZN(_22718_));
 OAI21_X1 _53408_ (.A(_22717_),
    .B1(_22701_),
    .B2(_22718_),
    .ZN(_03430_));
 MUX2_X1 _53409_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [526]),
    .B(_22659_),
    .S(_22713_),
    .Z(_03431_));
 MUX2_X1 _53410_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [527]),
    .B(_22428_),
    .S(_22713_),
    .Z(_03432_));
 MUX2_X1 _53411_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [528]),
    .B(_22542_),
    .S(_22713_),
    .Z(_03433_));
 MUX2_X1 _53412_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [529]),
    .B(_22641_),
    .S(_22700_),
    .Z(_03434_));
 MUX2_X1 _53413_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [530]),
    .B(_22596_),
    .S(_22700_),
    .Z(_03436_));
 MUX2_X1 _53414_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [531]),
    .B(_22516_),
    .S(_22700_),
    .Z(_03437_));
 MUX2_X1 _53415_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [532]),
    .B(_22573_),
    .S(_22700_),
    .Z(_03438_));
 MUX2_X1 _53416_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [533]),
    .B(_22492_),
    .S(_22700_),
    .Z(_03439_));
 BUF_X8 _53417_ (.A(_11015_),
    .Z(_22719_));
 NAND4_X1 _53418_ (.A1(_22716_),
    .A2(_22719_),
    .A3(_22602_),
    .A4(_21359_),
    .ZN(_22720_));
 INV_X2 _53419_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [534]),
    .ZN(_22721_));
 OAI21_X1 _53420_ (.A(_22720_),
    .B1(_22701_),
    .B2(_22721_),
    .ZN(_03440_));
 MUX2_X1 _53421_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [535]),
    .B(_22697_),
    .S(_22700_),
    .Z(_03441_));
 MUX2_X1 _53422_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [536]),
    .B(_22698_),
    .S(_22700_),
    .Z(_03442_));
 MUX2_X1 _53423_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [537]),
    .B(_22517_),
    .S(_22700_),
    .Z(_03443_));
 MUX2_X1 _53424_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [538]),
    .B(_22494_),
    .S(_22700_),
    .Z(_03444_));
 AND2_X4 _53425_ (.A1(_11158_),
    .A2(_21432_),
    .ZN(_22722_));
 BUF_X8 _53426_ (.A(_22722_),
    .Z(_22723_));
 BUF_X8 _53427_ (.A(_22723_),
    .Z(_22724_));
 MUX2_X1 _53428_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [441]),
    .B(_22685_),
    .S(_22724_),
    .Z(_03337_));
 MUX2_X1 _53429_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [442]),
    .B(_22667_),
    .S(_22724_),
    .Z(_03338_));
 NAND4_X1 _53430_ (.A1(_22563_),
    .A2(_21294_),
    .A3(_22677_),
    .A4(_22691_),
    .ZN(_22725_));
 INV_X1 _53431_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [443]),
    .ZN(_22726_));
 OAI21_X1 _53432_ (.A(_22725_),
    .B1(_22724_),
    .B2(_22726_),
    .ZN(_03339_));
 MUX2_X1 _53433_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [444]),
    .B(_22626_),
    .S(_22724_),
    .Z(_03340_));
 MUX2_X1 _53434_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [445]),
    .B(_21387_),
    .S(_22724_),
    .Z(_03341_));
 MUX2_X1 _53435_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [446]),
    .B(_22670_),
    .S(_22724_),
    .Z(_03342_));
 MUX2_X1 _53436_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [447]),
    .B(_22605_),
    .S(_22724_),
    .Z(_03343_));
 MUX2_X1 _53437_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [448]),
    .B(_22529_),
    .S(_22724_),
    .Z(_03344_));
 MUX2_X1 _53438_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [449]),
    .B(_22705_),
    .S(_22724_),
    .Z(_03345_));
 MUX2_X1 _53439_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [450]),
    .B(_21395_),
    .S(_22724_),
    .Z(_03347_));
 BUF_X8 _53440_ (.A(_22722_),
    .Z(_22727_));
 MUX2_X1 _53441_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [451]),
    .B(_22582_),
    .S(_22727_),
    .Z(_03348_));
 MUX2_X1 _53442_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [452]),
    .B(_22504_),
    .S(_22727_),
    .Z(_03349_));
 MUX2_X1 _53443_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [453]),
    .B(_22630_),
    .S(_22727_),
    .Z(_03350_));
 MUX2_X1 _53444_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [454]),
    .B(_22650_),
    .S(_22727_),
    .Z(_03351_));
 MUX2_X1 _53445_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [455]),
    .B(_22556_),
    .S(_22727_),
    .Z(_03352_));
 MUX2_X1 _53446_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [456]),
    .B(_22609_),
    .S(_22727_),
    .Z(_03353_));
 MUX2_X1 _53447_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [457]),
    .B(_22583_),
    .S(_22727_),
    .Z(_03354_));
 MUX2_X1 _53448_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [458]),
    .B(_10573_),
    .S(_22727_),
    .Z(_03355_));
 MUX2_X1 _53449_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [459]),
    .B(_22560_),
    .S(_22727_),
    .Z(_03356_));
 MUX2_X1 _53450_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [460]),
    .B(_22533_),
    .S(_22727_),
    .Z(_03358_));
 BUF_X16 _53451_ (.A(_22722_),
    .Z(_22728_));
 MUX2_X1 _53452_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [461]),
    .B(_22471_),
    .S(_22728_),
    .Z(_03359_));
 MUX2_X1 _53453_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [462]),
    .B(_22613_),
    .S(_22728_),
    .Z(_03360_));
 MUX2_X1 _53454_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [463]),
    .B(_22561_),
    .S(_22728_),
    .Z(_03361_));
 BUF_X8 _53455_ (.A(_08588_),
    .Z(_22729_));
 MUX2_X1 _53456_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [464]),
    .B(_22729_),
    .S(_22728_),
    .Z(_03362_));
 MUX2_X1 _53457_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [465]),
    .B(_22512_),
    .S(_22728_),
    .Z(_03363_));
 MUX2_X1 _53458_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [466]),
    .B(_22614_),
    .S(_22728_),
    .Z(_03364_));
 MUX2_X1 _53459_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [467]),
    .B(_22680_),
    .S(_22728_),
    .Z(_03365_));
 MUX2_X1 _53460_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [468]),
    .B(_22615_),
    .S(_22728_),
    .Z(_03366_));
 MUX2_X1 _53461_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [469]),
    .B(_22681_),
    .S(_22728_),
    .Z(_03367_));
 MUX2_X1 _53462_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [470]),
    .B(_22479_),
    .S(_22728_),
    .Z(_03369_));
 BUF_X8 _53463_ (.A(_22722_),
    .Z(_22730_));
 MUX2_X1 _53464_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [471]),
    .B(_22617_),
    .S(_22730_),
    .Z(_03370_));
 MUX2_X1 _53465_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [472]),
    .B(_22638_),
    .S(_22730_),
    .Z(_03371_));
 MUX2_X1 _53466_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [473]),
    .B(_22620_),
    .S(_22730_),
    .Z(_03372_));
 MUX2_X1 _53467_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [474]),
    .B(_22570_),
    .S(_22730_),
    .Z(_03373_));
 MUX2_X1 _53468_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [475]),
    .B(_22452_),
    .S(_22730_),
    .Z(_03374_));
 MUX2_X1 _53469_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [476]),
    .B(_22541_),
    .S(_22730_),
    .Z(_03375_));
 MUX2_X1 _53470_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [477]),
    .B(_22659_),
    .S(_22730_),
    .Z(_03376_));
 MUX2_X1 _53471_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [478]),
    .B(_22428_),
    .S(_22730_),
    .Z(_03377_));
 MUX2_X1 _53472_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [479]),
    .B(_22542_),
    .S(_22730_),
    .Z(_03378_));
 MUX2_X1 _53473_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [480]),
    .B(_22641_),
    .S(_22730_),
    .Z(_03380_));
 MUX2_X1 _53474_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [481]),
    .B(_22596_),
    .S(_22723_),
    .Z(_03381_));
 MUX2_X1 _53475_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [482]),
    .B(_21407_),
    .S(_22723_),
    .Z(_03382_));
 MUX2_X1 _53476_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [483]),
    .B(_22573_),
    .S(_22723_),
    .Z(_03383_));
 MUX2_X1 _53477_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [484]),
    .B(_21533_),
    .S(_22723_),
    .Z(_03384_));
 MUX2_X1 _53478_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [485]),
    .B(_21360_),
    .S(_22723_),
    .Z(_03385_));
 MUX2_X1 _53479_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [486]),
    .B(_22697_),
    .S(_22723_),
    .Z(_03386_));
 MUX2_X1 _53480_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [487]),
    .B(_22698_),
    .S(_22723_),
    .Z(_03387_));
 BUF_X4 _53481_ (.A(_21373_),
    .Z(_22731_));
 MUX2_X1 _53482_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [488]),
    .B(_22731_),
    .S(_22723_),
    .Z(_03388_));
 BUF_X2 _53483_ (.A(_21377_),
    .Z(_22732_));
 MUX2_X1 _53484_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [489]),
    .B(_22732_),
    .S(_22723_),
    .Z(_03389_));
 BUF_X16 _53485_ (.A(_11164_),
    .Z(_22733_));
 AND2_X4 _53486_ (.A1(_22733_),
    .A2(_21432_),
    .ZN(_22734_));
 BUF_X16 _53487_ (.A(_22734_),
    .Z(_22735_));
 BUF_X8 _53488_ (.A(_22735_),
    .Z(_22736_));
 MUX2_X1 _53489_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [392]),
    .B(_22685_),
    .S(_22736_),
    .Z(_03282_));
 MUX2_X1 _53490_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [393]),
    .B(_22667_),
    .S(_22736_),
    .Z(_03283_));
 MUX2_X1 _53491_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [394]),
    .B(_22601_),
    .S(_22736_),
    .Z(_03284_));
 MUX2_X1 _53492_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [395]),
    .B(_22626_),
    .S(_22736_),
    .Z(_03285_));
 MUX2_X1 _53493_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [396]),
    .B(_21387_),
    .S(_22736_),
    .Z(_03286_));
 MUX2_X1 _53494_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [397]),
    .B(_22670_),
    .S(_22736_),
    .Z(_03287_));
 MUX2_X1 _53495_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [398]),
    .B(_22605_),
    .S(_22736_),
    .Z(_03288_));
 MUX2_X1 _53496_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [399]),
    .B(_21582_),
    .S(_22736_),
    .Z(_03289_));
 BUF_X8 _53497_ (.A(_22734_),
    .Z(_22737_));
 MUX2_X1 _53498_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [400]),
    .B(_22705_),
    .S(_22737_),
    .Z(_03292_));
 MUX2_X1 _53499_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [401]),
    .B(_21395_),
    .S(_22737_),
    .Z(_03293_));
 MUX2_X1 _53500_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [402]),
    .B(_22582_),
    .S(_22737_),
    .Z(_03294_));
 MUX2_X1 _53501_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [403]),
    .B(_22504_),
    .S(_22737_),
    .Z(_03295_));
 MUX2_X1 _53502_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [404]),
    .B(_22630_),
    .S(_22737_),
    .Z(_03296_));
 MUX2_X1 _53503_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [405]),
    .B(_22650_),
    .S(_22737_),
    .Z(_03297_));
 MUX2_X1 _53504_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [406]),
    .B(_22556_),
    .S(_22737_),
    .Z(_03298_));
 BUF_X8 _53505_ (.A(_22360_),
    .Z(_22738_));
 NAND4_X1 _53506_ (.A1(_22588_),
    .A2(_08561_),
    .A3(_22738_),
    .A4(_22691_),
    .ZN(_22739_));
 INV_X1 _53507_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [407]),
    .ZN(_22740_));
 OAI21_X1 _53508_ (.A(_22739_),
    .B1(_22736_),
    .B2(_22740_),
    .ZN(_03299_));
 MUX2_X1 _53509_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [408]),
    .B(_22583_),
    .S(_22737_),
    .Z(_03300_));
 MUX2_X1 _53510_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [409]),
    .B(_10573_),
    .S(_22737_),
    .Z(_03301_));
 MUX2_X1 _53511_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [410]),
    .B(_22560_),
    .S(_22737_),
    .Z(_03303_));
 BUF_X16 _53512_ (.A(_22734_),
    .Z(_22741_));
 MUX2_X1 _53513_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [411]),
    .B(_10576_),
    .S(_22741_),
    .Z(_03304_));
 MUX2_X1 _53514_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [412]),
    .B(_22471_),
    .S(_22741_),
    .Z(_03305_));
 MUX2_X1 _53515_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [413]),
    .B(_22613_),
    .S(_22741_),
    .Z(_03306_));
 MUX2_X1 _53516_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [414]),
    .B(_22561_),
    .S(_22741_),
    .Z(_03307_));
 MUX2_X1 _53517_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [415]),
    .B(_22729_),
    .S(_22741_),
    .Z(_03308_));
 NAND4_X1 _53518_ (.A1(_22588_),
    .A2(_22025_),
    .A3(_22738_),
    .A4(_22691_),
    .ZN(_22742_));
 INV_X1 _53519_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [416]),
    .ZN(_22743_));
 OAI21_X1 _53520_ (.A(_22742_),
    .B1(_22736_),
    .B2(_22743_),
    .ZN(_03309_));
 MUX2_X1 _53521_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [417]),
    .B(_22614_),
    .S(_22741_),
    .Z(_03310_));
 MUX2_X1 _53522_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [418]),
    .B(_22680_),
    .S(_22741_),
    .Z(_03311_));
 MUX2_X1 _53523_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [419]),
    .B(_22615_),
    .S(_22741_),
    .Z(_03312_));
 MUX2_X1 _53524_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [420]),
    .B(_22681_),
    .S(_22741_),
    .Z(_03314_));
 MUX2_X1 _53525_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [421]),
    .B(_22479_),
    .S(_22741_),
    .Z(_03315_));
 BUF_X8 _53526_ (.A(_22734_),
    .Z(_22744_));
 MUX2_X1 _53527_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [422]),
    .B(_22617_),
    .S(_22744_),
    .Z(_03316_));
 MUX2_X1 _53528_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [423]),
    .B(_22638_),
    .S(_22744_),
    .Z(_03317_));
 MUX2_X1 _53529_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [424]),
    .B(_22620_),
    .S(_22744_),
    .Z(_03318_));
 MUX2_X1 _53530_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [425]),
    .B(_22570_),
    .S(_22744_),
    .Z(_03319_));
 MUX2_X1 _53531_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [426]),
    .B(_22452_),
    .S(_22744_),
    .Z(_03320_));
 MUX2_X1 _53532_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [427]),
    .B(_22541_),
    .S(_22744_),
    .Z(_03321_));
 MUX2_X1 _53533_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [428]),
    .B(_22659_),
    .S(_22744_),
    .Z(_03322_));
 MUX2_X1 _53534_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [429]),
    .B(_10605_),
    .S(_22744_),
    .Z(_03323_));
 MUX2_X1 _53535_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [430]),
    .B(_22542_),
    .S(_22744_),
    .Z(_03325_));
 MUX2_X1 _53536_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [431]),
    .B(_22641_),
    .S(_22744_),
    .Z(_03326_));
 MUX2_X1 _53537_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [432]),
    .B(_22596_),
    .S(_22735_),
    .Z(_03327_));
 MUX2_X1 _53538_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [433]),
    .B(_21407_),
    .S(_22735_),
    .Z(_03328_));
 MUX2_X1 _53539_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [434]),
    .B(_22573_),
    .S(_22735_),
    .Z(_03329_));
 MUX2_X1 _53540_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [435]),
    .B(_21533_),
    .S(_22735_),
    .Z(_03330_));
 MUX2_X1 _53541_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [436]),
    .B(_21360_),
    .S(_22735_),
    .Z(_03331_));
 MUX2_X1 _53542_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [437]),
    .B(_22697_),
    .S(_22735_),
    .Z(_03332_));
 MUX2_X1 _53543_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [438]),
    .B(_22698_),
    .S(_22735_),
    .Z(_03333_));
 MUX2_X1 _53544_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [439]),
    .B(_22731_),
    .S(_22735_),
    .Z(_03334_));
 MUX2_X1 _53545_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [440]),
    .B(_22732_),
    .S(_22735_),
    .Z(_03336_));
 AND2_X4 _53546_ (.A1(_11170_),
    .A2(_21574_),
    .ZN(_22745_));
 BUF_X8 _53547_ (.A(_22745_),
    .Z(_22746_));
 BUF_X8 _53548_ (.A(_22746_),
    .Z(_22747_));
 MUX2_X1 _53549_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [343]),
    .B(_22685_),
    .S(_22747_),
    .Z(_03228_));
 MUX2_X1 _53550_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [344]),
    .B(_22667_),
    .S(_22747_),
    .Z(_03229_));
 MUX2_X1 _53551_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [345]),
    .B(_22601_),
    .S(_22747_),
    .Z(_03230_));
 MUX2_X1 _53552_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [346]),
    .B(_22626_),
    .S(_22747_),
    .Z(_03231_));
 MUX2_X1 _53553_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [347]),
    .B(_21387_),
    .S(_22747_),
    .Z(_03232_));
 MUX2_X1 _53554_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [348]),
    .B(_22670_),
    .S(_22747_),
    .Z(_03233_));
 BUF_X8 _53555_ (.A(_22745_),
    .Z(_22748_));
 MUX2_X1 _53556_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [349]),
    .B(_22605_),
    .S(_22748_),
    .Z(_03234_));
 BUF_X4 _53557_ (.A(_11177_),
    .Z(_22749_));
 NAND4_X1 _53558_ (.A1(_22399_),
    .A2(_21303_),
    .A3(_22738_),
    .A4(_22749_),
    .ZN(_22750_));
 INV_X1 _53559_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [350]),
    .ZN(_22751_));
 OAI21_X1 _53560_ (.A(_22750_),
    .B1(_22747_),
    .B2(_22751_),
    .ZN(_03236_));
 MUX2_X1 _53561_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [351]),
    .B(_22705_),
    .S(_22748_),
    .Z(_03237_));
 MUX2_X1 _53562_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [352]),
    .B(_21395_),
    .S(_22748_),
    .Z(_03238_));
 MUX2_X1 _53563_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [353]),
    .B(_22582_),
    .S(_22748_),
    .Z(_03239_));
 MUX2_X1 _53564_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [354]),
    .B(_21506_),
    .S(_22748_),
    .Z(_03240_));
 MUX2_X1 _53565_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [355]),
    .B(_22630_),
    .S(_22748_),
    .Z(_03241_));
 MUX2_X1 _53566_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [356]),
    .B(_22650_),
    .S(_22748_),
    .Z(_03242_));
 MUX2_X1 _53567_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [357]),
    .B(_10570_),
    .S(_22748_),
    .Z(_03243_));
 MUX2_X1 _53568_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [358]),
    .B(_22609_),
    .S(_22748_),
    .Z(_03244_));
 MUX2_X1 _53569_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [359]),
    .B(_22583_),
    .S(_22748_),
    .Z(_03245_));
 BUF_X8 _53570_ (.A(_22745_),
    .Z(_22752_));
 MUX2_X1 _53571_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [360]),
    .B(_10573_),
    .S(_22752_),
    .Z(_03247_));
 MUX2_X1 _53572_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [361]),
    .B(_10600_),
    .S(_22752_),
    .Z(_03248_));
 MUX2_X1 _53573_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [362]),
    .B(_10576_),
    .S(_22752_),
    .Z(_03249_));
 MUX2_X1 _53574_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [363]),
    .B(_10577_),
    .S(_22752_),
    .Z(_03250_));
 MUX2_X1 _53575_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [364]),
    .B(_22613_),
    .S(_22752_),
    .Z(_03251_));
 MUX2_X1 _53576_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [365]),
    .B(_22561_),
    .S(_22752_),
    .Z(_03252_));
 MUX2_X1 _53577_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [366]),
    .B(_22729_),
    .S(_22752_),
    .Z(_03253_));
 MUX2_X1 _53578_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [367]),
    .B(_10602_),
    .S(_22752_),
    .Z(_03254_));
 MUX2_X1 _53579_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [368]),
    .B(_22614_),
    .S(_22752_),
    .Z(_03255_));
 MUX2_X1 _53580_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [369]),
    .B(_22680_),
    .S(_22752_),
    .Z(_03256_));
 BUF_X8 _53581_ (.A(_22745_),
    .Z(_22753_));
 MUX2_X1 _53582_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [370]),
    .B(_22615_),
    .S(_22753_),
    .Z(_03258_));
 MUX2_X1 _53583_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [371]),
    .B(_22681_),
    .S(_22753_),
    .Z(_03259_));
 MUX2_X1 _53584_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [372]),
    .B(_10586_),
    .S(_22753_),
    .Z(_03260_));
 MUX2_X1 _53585_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [373]),
    .B(_22617_),
    .S(_22753_),
    .Z(_03261_));
 MUX2_X1 _53586_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [374]),
    .B(_22638_),
    .S(_22753_),
    .Z(_03262_));
 MUX2_X1 _53587_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [375]),
    .B(_22620_),
    .S(_22753_),
    .Z(_03263_));
 MUX2_X1 _53588_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [376]),
    .B(_22570_),
    .S(_22753_),
    .Z(_03264_));
 MUX2_X1 _53589_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [377]),
    .B(_22452_),
    .S(_22753_),
    .Z(_03265_));
 MUX2_X1 _53590_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [378]),
    .B(_10592_),
    .S(_22753_),
    .Z(_03266_));
 MUX2_X1 _53591_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [379]),
    .B(_22659_),
    .S(_22753_),
    .Z(_03267_));
 MUX2_X1 _53592_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [380]),
    .B(_10605_),
    .S(_22746_),
    .Z(_03269_));
 NAND4_X1 _53593_ (.A1(_10805_),
    .A2(_08635_),
    .A3(_22738_),
    .A4(_22749_),
    .ZN(_22754_));
 INV_X1 _53594_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [381]),
    .ZN(_22755_));
 OAI21_X1 _53595_ (.A(_22754_),
    .B1(_22747_),
    .B2(_22755_),
    .ZN(_03270_));
 MUX2_X1 _53596_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [382]),
    .B(_22641_),
    .S(_22746_),
    .Z(_03271_));
 MUX2_X1 _53597_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [383]),
    .B(_22596_),
    .S(_22746_),
    .Z(_03272_));
 MUX2_X1 _53598_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [384]),
    .B(_21407_),
    .S(_22746_),
    .Z(_03273_));
 MUX2_X1 _53599_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [385]),
    .B(_21461_),
    .S(_22746_),
    .Z(_03274_));
 NAND4_X1 _53600_ (.A1(_10805_),
    .A2(_22719_),
    .A3(_11178_),
    .A4(_21738_),
    .ZN(_22756_));
 INV_X1 _53601_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [386]),
    .ZN(_22757_));
 OAI21_X1 _53602_ (.A(_22756_),
    .B1(_22747_),
    .B2(_22757_),
    .ZN(_03275_));
 NAND4_X1 _53603_ (.A1(_10805_),
    .A2(_22719_),
    .A3(_11178_),
    .A4(_21359_),
    .ZN(_22758_));
 INV_X1 _53604_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [387]),
    .ZN(_22759_));
 OAI21_X1 _53605_ (.A(_22758_),
    .B1(_22747_),
    .B2(_22759_),
    .ZN(_03276_));
 MUX2_X1 _53606_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [388]),
    .B(_22697_),
    .S(_22746_),
    .Z(_03277_));
 MUX2_X1 _53607_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [389]),
    .B(_22698_),
    .S(_22746_),
    .Z(_03278_));
 MUX2_X1 _53608_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [390]),
    .B(_22731_),
    .S(_22746_),
    .Z(_03280_));
 MUX2_X1 _53609_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [391]),
    .B(_22732_),
    .S(_22746_),
    .Z(_03281_));
 AND2_X4 _53610_ (.A1(_11181_),
    .A2(_21412_),
    .ZN(_22760_));
 BUF_X8 _53611_ (.A(_22760_),
    .Z(_22761_));
 BUF_X8 _53612_ (.A(_22761_),
    .Z(_22762_));
 MUX2_X1 _53613_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [294]),
    .B(_22685_),
    .S(_22762_),
    .Z(_02987_));
 MUX2_X1 _53614_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [295]),
    .B(_22667_),
    .S(_22762_),
    .Z(_02998_));
 MUX2_X1 _53615_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [296]),
    .B(_22601_),
    .S(_22762_),
    .Z(_03009_));
 MUX2_X1 _53616_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [297]),
    .B(_22626_),
    .S(_22762_),
    .Z(_03020_));
 MUX2_X1 _53617_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [298]),
    .B(_21387_),
    .S(_22762_),
    .Z(_03031_));
 BUF_X8 _53618_ (.A(_22760_),
    .Z(_22763_));
 MUX2_X1 _53619_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [299]),
    .B(_22670_),
    .S(_22763_),
    .Z(_03042_));
 MUX2_X1 _53620_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [300]),
    .B(_22605_),
    .S(_22763_),
    .Z(_03055_));
 NAND4_X1 _53621_ (.A1(_22422_),
    .A2(_21303_),
    .A3(_22738_),
    .A4(_22749_),
    .ZN(_22764_));
 INV_X1 _53622_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [301]),
    .ZN(_22765_));
 OAI21_X1 _53623_ (.A(_22764_),
    .B1(_22762_),
    .B2(_22765_),
    .ZN(_03066_));
 MUX2_X1 _53624_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [302]),
    .B(_22705_),
    .S(_22763_),
    .Z(_03077_));
 MUX2_X1 _53625_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [303]),
    .B(_21395_),
    .S(_22763_),
    .Z(_03088_));
 MUX2_X1 _53626_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [304]),
    .B(_21446_),
    .S(_22763_),
    .Z(_03099_));
 MUX2_X1 _53627_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [305]),
    .B(_21506_),
    .S(_22763_),
    .Z(_03110_));
 MUX2_X1 _53628_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [306]),
    .B(_22630_),
    .S(_22763_),
    .Z(_03121_));
 MUX2_X1 _53629_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [307]),
    .B(_22650_),
    .S(_22763_),
    .Z(_03132_));
 MUX2_X1 _53630_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [308]),
    .B(_10570_),
    .S(_22763_),
    .Z(_03143_));
 MUX2_X1 _53631_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [309]),
    .B(_22609_),
    .S(_22763_),
    .Z(_03154_));
 NAND4_X1 _53632_ (.A1(_22422_),
    .A2(_22371_),
    .A3(_22738_),
    .A4(_22749_),
    .ZN(_22766_));
 INV_X1 _53633_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [310]),
    .ZN(_22767_));
 OAI21_X1 _53634_ (.A(_22766_),
    .B1(_22762_),
    .B2(_22767_),
    .ZN(_03166_));
 BUF_X8 _53635_ (.A(_22760_),
    .Z(_22768_));
 MUX2_X1 _53636_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [311]),
    .B(_10573_),
    .S(_22768_),
    .Z(_03177_));
 MUX2_X1 _53637_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [312]),
    .B(_10600_),
    .S(_22768_),
    .Z(_03188_));
 MUX2_X1 _53638_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [313]),
    .B(_10576_),
    .S(_22768_),
    .Z(_03195_));
 MUX2_X1 _53639_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [314]),
    .B(_10577_),
    .S(_22768_),
    .Z(_03196_));
 MUX2_X1 _53640_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [315]),
    .B(_22613_),
    .S(_22768_),
    .Z(_03197_));
 MUX2_X1 _53641_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [316]),
    .B(_22561_),
    .S(_22768_),
    .Z(_03198_));
 MUX2_X1 _53642_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [317]),
    .B(_22729_),
    .S(_22768_),
    .Z(_03199_));
 NAND4_X1 _53643_ (.A1(_10819_),
    .A2(_22025_),
    .A3(_22738_),
    .A4(_22749_),
    .ZN(_22769_));
 INV_X1 _53644_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [318]),
    .ZN(_22770_));
 OAI21_X1 _53645_ (.A(_22769_),
    .B1(_22762_),
    .B2(_22770_),
    .ZN(_03200_));
 NAND4_X4 _53646_ (.A1(_10819_),
    .A2(_21757_),
    .A3(_22738_),
    .A4(_22749_),
    .ZN(_22771_));
 INV_X1 _53647_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [319]),
    .ZN(_22772_));
 OAI21_X1 _53648_ (.A(_22771_),
    .B1(_22762_),
    .B2(_22772_),
    .ZN(_03201_));
 MUX2_X1 _53649_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [320]),
    .B(_22680_),
    .S(_22768_),
    .Z(_03203_));
 MUX2_X1 _53650_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [321]),
    .B(_22615_),
    .S(_22768_),
    .Z(_03204_));
 MUX2_X1 _53651_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [322]),
    .B(_22681_),
    .S(_22768_),
    .Z(_03205_));
 BUF_X16 _53652_ (.A(_22760_),
    .Z(_22773_));
 MUX2_X1 _53653_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [323]),
    .B(_10586_),
    .S(_22773_),
    .Z(_03206_));
 MUX2_X1 _53654_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [324]),
    .B(_22617_),
    .S(_22773_),
    .Z(_03207_));
 MUX2_X1 _53655_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [325]),
    .B(_22638_),
    .S(_22773_),
    .Z(_03208_));
 MUX2_X1 _53656_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [326]),
    .B(_22620_),
    .S(_22773_),
    .Z(_03209_));
 MUX2_X1 _53657_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [327]),
    .B(_10604_),
    .S(_22773_),
    .Z(_03210_));
 MUX2_X1 _53658_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [328]),
    .B(_10591_),
    .S(_22773_),
    .Z(_03211_));
 MUX2_X1 _53659_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [329]),
    .B(_10592_),
    .S(_22773_),
    .Z(_03212_));
 MUX2_X1 _53660_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [330]),
    .B(_22659_),
    .S(_22773_),
    .Z(_03214_));
 MUX2_X1 _53661_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [331]),
    .B(_10605_),
    .S(_22773_),
    .Z(_03215_));
 MUX2_X1 _53662_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [332]),
    .B(_10595_),
    .S(_22773_),
    .Z(_03216_));
 MUX2_X1 _53663_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [333]),
    .B(_22641_),
    .S(_22761_),
    .Z(_03217_));
 MUX2_X1 _53664_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [334]),
    .B(_21763_),
    .S(_22761_),
    .Z(_03218_));
 MUX2_X1 _53665_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [335]),
    .B(_21407_),
    .S(_22761_),
    .Z(_03219_));
 MUX2_X1 _53666_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [336]),
    .B(_21461_),
    .S(_22761_),
    .Z(_03220_));
 BUF_X4 _53667_ (.A(_11177_),
    .Z(_22774_));
 NAND4_X2 _53668_ (.A1(_10819_),
    .A2(_22719_),
    .A3(_22774_),
    .A4(_21355_),
    .ZN(_22775_));
 INV_X1 _53669_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [337]),
    .ZN(_22776_));
 OAI21_X1 _53670_ (.A(_22775_),
    .B1(_22762_),
    .B2(_22776_),
    .ZN(_03221_));
 MUX2_X1 _53671_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [338]),
    .B(_21360_),
    .S(_22761_),
    .Z(_03222_));
 MUX2_X1 _53672_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [339]),
    .B(_22697_),
    .S(_22761_),
    .Z(_03223_));
 MUX2_X1 _53673_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [340]),
    .B(_22698_),
    .S(_22761_),
    .Z(_03225_));
 MUX2_X1 _53674_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [341]),
    .B(_22731_),
    .S(_22761_),
    .Z(_03226_));
 MUX2_X1 _53675_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [342]),
    .B(_22732_),
    .S(_22761_),
    .Z(_03227_));
 BUF_X8 _53676_ (.A(_11186_),
    .Z(_22777_));
 AND2_X4 _53677_ (.A1(_22777_),
    .A2(_21574_),
    .ZN(_22778_));
 BUF_X8 _53678_ (.A(_22778_),
    .Z(_22779_));
 BUF_X8 _53679_ (.A(_22779_),
    .Z(_22780_));
 MUX2_X1 _53680_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [245]),
    .B(_22685_),
    .S(_22780_),
    .Z(_02443_));
 MUX2_X1 _53681_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [246]),
    .B(_22667_),
    .S(_22780_),
    .Z(_02454_));
 MUX2_X1 _53682_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [247]),
    .B(_22601_),
    .S(_22780_),
    .Z(_02465_));
 MUX2_X1 _53683_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [248]),
    .B(_22626_),
    .S(_22780_),
    .Z(_02476_));
 MUX2_X1 _53684_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [249]),
    .B(_21387_),
    .S(_22780_),
    .Z(_02487_));
 MUX2_X1 _53685_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [250]),
    .B(_22670_),
    .S(_22780_),
    .Z(_02499_));
 BUF_X16 _53686_ (.A(_22778_),
    .Z(_22781_));
 MUX2_X1 _53687_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [251]),
    .B(_21578_),
    .S(_22781_),
    .Z(_02510_));
 MUX2_X1 _53688_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [252]),
    .B(_21582_),
    .S(_22781_),
    .Z(_02521_));
 MUX2_X1 _53689_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [253]),
    .B(_22705_),
    .S(_22781_),
    .Z(_02532_));
 MUX2_X1 _53690_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [254]),
    .B(_21395_),
    .S(_22781_),
    .Z(_02543_));
 MUX2_X1 _53691_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [255]),
    .B(_21446_),
    .S(_22781_),
    .Z(_02554_));
 MUX2_X1 _53692_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [256]),
    .B(_21506_),
    .S(_22781_),
    .Z(_02565_));
 MUX2_X1 _53693_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [257]),
    .B(_22630_),
    .S(_22781_),
    .Z(_02576_));
 MUX2_X1 _53694_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [258]),
    .B(_22650_),
    .S(_22781_),
    .Z(_02587_));
 MUX2_X1 _53695_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [259]),
    .B(_10570_),
    .S(_22781_),
    .Z(_02598_));
 MUX2_X1 _53696_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [260]),
    .B(_22609_),
    .S(_22781_),
    .Z(_02610_));
 NAND4_X1 _53697_ (.A1(_10832_),
    .A2(_22371_),
    .A3(_22738_),
    .A4(_22749_),
    .ZN(_22782_));
 INV_X1 _53698_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [261]),
    .ZN(_22783_));
 OAI21_X1 _53699_ (.A(_22782_),
    .B1(_22780_),
    .B2(_22783_),
    .ZN(_02621_));
 BUF_X8 _53700_ (.A(_22778_),
    .Z(_22784_));
 MUX2_X1 _53701_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [262]),
    .B(_10573_),
    .S(_22784_),
    .Z(_02632_));
 MUX2_X1 _53702_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [263]),
    .B(_10600_),
    .S(_22784_),
    .Z(_02643_));
 MUX2_X1 _53703_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [264]),
    .B(_10576_),
    .S(_22784_),
    .Z(_02654_));
 MUX2_X1 _53704_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [265]),
    .B(_10577_),
    .S(_22784_),
    .Z(_02665_));
 MUX2_X1 _53705_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [266]),
    .B(_22613_),
    .S(_22784_),
    .Z(_02676_));
 NAND4_X1 _53706_ (.A1(_10832_),
    .A2(_08584_),
    .A3(_22738_),
    .A4(_22749_),
    .ZN(_22785_));
 INV_X1 _53707_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [267]),
    .ZN(_22786_));
 OAI21_X1 _53708_ (.A(_22785_),
    .B1(_22780_),
    .B2(_22786_),
    .ZN(_02687_));
 MUX2_X1 _53709_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [268]),
    .B(_22729_),
    .S(_22784_),
    .Z(_02698_));
 BUF_X4 _53710_ (.A(_22360_),
    .Z(_22787_));
 NAND4_X1 _53711_ (.A1(_10832_),
    .A2(_08591_),
    .A3(_22787_),
    .A4(_22749_),
    .ZN(_22788_));
 INV_X1 _53712_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [269]),
    .ZN(_22789_));
 OAI21_X1 _53713_ (.A(_22788_),
    .B1(_22780_),
    .B2(_22789_),
    .ZN(_02709_));
 MUX2_X1 _53714_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [270]),
    .B(_22614_),
    .S(_22784_),
    .Z(_02721_));
 MUX2_X1 _53715_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [271]),
    .B(_22680_),
    .S(_22784_),
    .Z(_02732_));
 MUX2_X1 _53716_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [272]),
    .B(_10584_),
    .S(_22784_),
    .Z(_02743_));
 MUX2_X1 _53717_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [273]),
    .B(_22681_),
    .S(_22784_),
    .Z(_02754_));
 BUF_X8 _53718_ (.A(_22778_),
    .Z(_22790_));
 MUX2_X1 _53719_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [274]),
    .B(_10586_),
    .S(_22790_),
    .Z(_02765_));
 MUX2_X1 _53720_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [275]),
    .B(_10587_),
    .S(_22790_),
    .Z(_02776_));
 MUX2_X1 _53721_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [276]),
    .B(_22638_),
    .S(_22790_),
    .Z(_02787_));
 MUX2_X1 _53722_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [277]),
    .B(_10603_),
    .S(_22790_),
    .Z(_02798_));
 MUX2_X1 _53723_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [278]),
    .B(_10604_),
    .S(_22790_),
    .Z(_02809_));
 MUX2_X1 _53724_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [279]),
    .B(_10591_),
    .S(_22790_),
    .Z(_02820_));
 MUX2_X1 _53725_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [280]),
    .B(_10592_),
    .S(_22790_),
    .Z(_02832_));
 MUX2_X1 _53726_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [281]),
    .B(_22659_),
    .S(_22790_),
    .Z(_02843_));
 MUX2_X1 _53727_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [282]),
    .B(_10605_),
    .S(_22790_),
    .Z(_02854_));
 NAND4_X1 _53728_ (.A1(_10832_),
    .A2(_08635_),
    .A3(_22787_),
    .A4(_22749_),
    .ZN(_22791_));
 INV_X4 _53729_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [283]),
    .ZN(_22792_));
 OAI21_X1 _53730_ (.A(_22791_),
    .B1(_22780_),
    .B2(_22792_),
    .ZN(_02865_));
 MUX2_X1 _53731_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [284]),
    .B(_22641_),
    .S(_22790_),
    .Z(_02876_));
 MUX2_X1 _53732_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [285]),
    .B(_21763_),
    .S(_22779_),
    .Z(_02887_));
 MUX2_X1 _53733_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [286]),
    .B(_21407_),
    .S(_22779_),
    .Z(_02898_));
 MUX2_X1 _53734_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [287]),
    .B(_21461_),
    .S(_22779_),
    .Z(_02909_));
 MUX2_X1 _53735_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [288]),
    .B(_21533_),
    .S(_22779_),
    .Z(_02920_));
 MUX2_X1 _53736_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [289]),
    .B(_21360_),
    .S(_22779_),
    .Z(_02931_));
 MUX2_X1 _53737_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [290]),
    .B(_22697_),
    .S(_22779_),
    .Z(_02943_));
 MUX2_X1 _53738_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [291]),
    .B(_22698_),
    .S(_22779_),
    .Z(_02954_));
 MUX2_X1 _53739_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [292]),
    .B(_22731_),
    .S(_22779_),
    .Z(_02965_));
 MUX2_X1 _53740_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [293]),
    .B(_22732_),
    .S(_22779_),
    .Z(_02976_));
 AND2_X4 _53741_ (.A1(_11190_),
    .A2(_21432_),
    .ZN(_22793_));
 BUF_X16 _53742_ (.A(_22793_),
    .Z(_22794_));
 BUF_X8 _53743_ (.A(_22794_),
    .Z(_22795_));
 MUX2_X1 _53744_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [196]),
    .B(_22685_),
    .S(_22795_),
    .Z(_01898_));
 MUX2_X1 _53745_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [197]),
    .B(_22667_),
    .S(_22795_),
    .Z(_01909_));
 BUF_X4 _53746_ (.A(_11177_),
    .Z(_22796_));
 NAND4_X1 _53747_ (.A1(_10845_),
    .A2(_21294_),
    .A3(_22787_),
    .A4(_22796_),
    .ZN(_22797_));
 INV_X1 _53748_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [198]),
    .ZN(_22798_));
 OAI21_X1 _53749_ (.A(_22797_),
    .B1(_22795_),
    .B2(_22798_),
    .ZN(_01920_));
 MUX2_X1 _53750_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [199]),
    .B(_22626_),
    .S(_22795_),
    .Z(_01931_));
 MUX2_X1 _53751_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [200]),
    .B(_21387_),
    .S(_22795_),
    .Z(_01944_));
 MUX2_X1 _53752_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [201]),
    .B(_22670_),
    .S(_22795_),
    .Z(_01955_));
 MUX2_X1 _53753_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [202]),
    .B(_21578_),
    .S(_22795_),
    .Z(_01966_));
 MUX2_X1 _53754_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [203]),
    .B(_21582_),
    .S(_22795_),
    .Z(_01977_));
 BUF_X8 _53755_ (.A(_22793_),
    .Z(_22799_));
 MUX2_X1 _53756_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [204]),
    .B(_22705_),
    .S(_22799_),
    .Z(_01988_));
 MUX2_X1 _53757_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [205]),
    .B(_21395_),
    .S(_22799_),
    .Z(_01999_));
 MUX2_X1 _53758_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [206]),
    .B(_21446_),
    .S(_22799_),
    .Z(_02010_));
 MUX2_X1 _53759_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [207]),
    .B(_21506_),
    .S(_22799_),
    .Z(_02021_));
 MUX2_X1 _53760_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [208]),
    .B(_22630_),
    .S(_22799_),
    .Z(_02032_));
 MUX2_X1 _53761_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [209]),
    .B(_22650_),
    .S(_22799_),
    .Z(_02043_));
 MUX2_X1 _53762_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [210]),
    .B(_10570_),
    .S(_22799_),
    .Z(_02055_));
 MUX2_X1 _53763_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [211]),
    .B(_10571_),
    .S(_22799_),
    .Z(_02066_));
 MUX2_X1 _53764_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [212]),
    .B(_22583_),
    .S(_22799_),
    .Z(_02077_));
 MUX2_X1 _53765_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [213]),
    .B(_10573_),
    .S(_22799_),
    .Z(_02088_));
 BUF_X16 _53766_ (.A(_22793_),
    .Z(_22800_));
 MUX2_X1 _53767_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [214]),
    .B(_10600_),
    .S(_22800_),
    .Z(_02099_));
 MUX2_X1 _53768_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [215]),
    .B(_10576_),
    .S(_22800_),
    .Z(_02110_));
 MUX2_X1 _53769_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [216]),
    .B(_10577_),
    .S(_22800_),
    .Z(_02121_));
 MUX2_X1 _53770_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [217]),
    .B(_22613_),
    .S(_22800_),
    .Z(_02132_));
 MUX2_X1 _53771_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [218]),
    .B(_10579_),
    .S(_22800_),
    .Z(_02143_));
 MUX2_X1 _53772_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [219]),
    .B(_22729_),
    .S(_22800_),
    .Z(_02154_));
 MUX2_X1 _53773_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [220]),
    .B(_10602_),
    .S(_22800_),
    .Z(_02166_));
 MUX2_X1 _53774_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [221]),
    .B(_10582_),
    .S(_22800_),
    .Z(_02177_));
 MUX2_X1 _53775_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [222]),
    .B(_22680_),
    .S(_22800_),
    .Z(_02188_));
 MUX2_X1 _53776_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [223]),
    .B(_10584_),
    .S(_22800_),
    .Z(_02199_));
 BUF_X8 _53777_ (.A(_22793_),
    .Z(_22801_));
 MUX2_X1 _53778_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [224]),
    .B(_22681_),
    .S(_22801_),
    .Z(_02210_));
 MUX2_X1 _53779_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [225]),
    .B(_10586_),
    .S(_22801_),
    .Z(_02221_));
 MUX2_X1 _53780_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [226]),
    .B(_10587_),
    .S(_22801_),
    .Z(_02232_));
 MUX2_X1 _53781_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [227]),
    .B(_10588_),
    .S(_22801_),
    .Z(_02243_));
 MUX2_X1 _53782_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [228]),
    .B(_10603_),
    .S(_22801_),
    .Z(_02254_));
 MUX2_X1 _53783_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [229]),
    .B(_10604_),
    .S(_22801_),
    .Z(_02265_));
 NAND4_X1 _53784_ (.A1(_10845_),
    .A2(_21562_),
    .A3(_22787_),
    .A4(_22796_),
    .ZN(_22802_));
 INV_X1 _53785_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [230]),
    .ZN(_22803_));
 OAI21_X1 _53786_ (.A(_22802_),
    .B1(_22795_),
    .B2(_22803_),
    .ZN(_02277_));
 MUX2_X1 _53787_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [231]),
    .B(_10592_),
    .S(_22801_),
    .Z(_02288_));
 MUX2_X1 _53788_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [232]),
    .B(_22659_),
    .S(_22801_),
    .Z(_02299_));
 MUX2_X1 _53789_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [233]),
    .B(_10605_),
    .S(_22801_),
    .Z(_02310_));
 MUX2_X1 _53790_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [234]),
    .B(_10595_),
    .S(_22801_),
    .Z(_02321_));
 MUX2_X1 _53791_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [235]),
    .B(_21595_),
    .S(_22794_),
    .Z(_02332_));
 MUX2_X1 _53792_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [236]),
    .B(_21763_),
    .S(_22794_),
    .Z(_02343_));
 MUX2_X1 _53793_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [237]),
    .B(_21407_),
    .S(_22794_),
    .Z(_02354_));
 MUX2_X1 _53794_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [238]),
    .B(_21461_),
    .S(_22794_),
    .Z(_02365_));
 NAND4_X1 _53795_ (.A1(_10845_),
    .A2(_22719_),
    .A3(_22774_),
    .A4(_21355_),
    .ZN(_22804_));
 INV_X1 _53796_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [239]),
    .ZN(_22805_));
 OAI21_X1 _53797_ (.A(_22804_),
    .B1(_22795_),
    .B2(_22805_),
    .ZN(_02376_));
 MUX2_X1 _53798_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [240]),
    .B(_21360_),
    .S(_22794_),
    .Z(_02388_));
 MUX2_X1 _53799_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [241]),
    .B(_22697_),
    .S(_22794_),
    .Z(_02399_));
 MUX2_X1 _53800_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [242]),
    .B(_22698_),
    .S(_22794_),
    .Z(_02410_));
 MUX2_X1 _53801_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [243]),
    .B(_22731_),
    .S(_22794_),
    .Z(_02421_));
 MUX2_X1 _53802_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [244]),
    .B(_22732_),
    .S(_22794_),
    .Z(_02432_));
 BUF_X16 _53803_ (.A(_11195_),
    .Z(_22806_));
 AND2_X4 _53804_ (.A1(_22806_),
    .A2(_21679_),
    .ZN(_22807_));
 BUF_X16 _53805_ (.A(_22807_),
    .Z(_22808_));
 BUF_X8 _53806_ (.A(_22808_),
    .Z(_22809_));
 MUX2_X1 _53807_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [147]),
    .B(_22685_),
    .S(_22809_),
    .Z(_01354_));
 MUX2_X1 _53808_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [148]),
    .B(_22667_),
    .S(_22809_),
    .Z(_01365_));
 MUX2_X1 _53809_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [149]),
    .B(_22601_),
    .S(_22809_),
    .Z(_01376_));
 BUF_X16 _53810_ (.A(_22807_),
    .Z(_22810_));
 MUX2_X1 _53811_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [150]),
    .B(_21608_),
    .S(_22810_),
    .Z(_01388_));
 NAND4_X1 _53812_ (.A1(_22498_),
    .A2(_21297_),
    .A3(_22787_),
    .A4(_22796_),
    .ZN(_22811_));
 INV_X1 _53813_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [151]),
    .ZN(_22812_));
 OAI21_X1 _53814_ (.A(_22811_),
    .B1(_22809_),
    .B2(_22812_),
    .ZN(_01399_));
 MUX2_X1 _53815_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [152]),
    .B(_22670_),
    .S(_22810_),
    .Z(_01410_));
 MUX2_X1 _53816_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [153]),
    .B(_21578_),
    .S(_22810_),
    .Z(_01421_));
 MUX2_X1 _53817_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [154]),
    .B(_21582_),
    .S(_22810_),
    .Z(_01432_));
 MUX2_X1 _53818_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [155]),
    .B(_22705_),
    .S(_22810_),
    .Z(_01443_));
 MUX2_X1 _53819_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [156]),
    .B(_21395_),
    .S(_22810_),
    .Z(_01454_));
 NAND4_X1 _53820_ (.A1(_22498_),
    .A2(_21309_),
    .A3(_22787_),
    .A4(_22796_),
    .ZN(_22813_));
 INV_X1 _53821_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [157]),
    .ZN(_22814_));
 OAI21_X1 _53822_ (.A(_22813_),
    .B1(_22809_),
    .B2(_22814_),
    .ZN(_01465_));
 MUX2_X1 _53823_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [158]),
    .B(_21506_),
    .S(_22810_),
    .Z(_01476_));
 MUX2_X1 _53824_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [159]),
    .B(_10563_),
    .S(_22810_),
    .Z(_01487_));
 MUX2_X1 _53825_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [160]),
    .B(_10569_),
    .S(_22810_),
    .Z(_01499_));
 MUX2_X1 _53826_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [161]),
    .B(_10570_),
    .S(_22810_),
    .Z(_01510_));
 BUF_X8 _53827_ (.A(_22807_),
    .Z(_22815_));
 MUX2_X1 _53828_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [162]),
    .B(_10571_),
    .S(_22815_),
    .Z(_01521_));
 NAND4_X2 _53829_ (.A1(_22498_),
    .A2(_08564_),
    .A3(_22787_),
    .A4(_22796_),
    .ZN(_22816_));
 INV_X1 _53830_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [163]),
    .ZN(_22817_));
 OAI21_X1 _53831_ (.A(_22816_),
    .B1(_22809_),
    .B2(_22817_),
    .ZN(_01532_));
 NAND4_X1 _53832_ (.A1(_22498_),
    .A2(_08567_),
    .A3(_22787_),
    .A4(_22796_),
    .ZN(_22818_));
 INV_X1 _53833_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [164]),
    .ZN(_22819_));
 OAI21_X1 _53834_ (.A(_22818_),
    .B1(_22809_),
    .B2(_22819_),
    .ZN(_01543_));
 NAND4_X1 _53835_ (.A1(_10781_),
    .A2(_08571_),
    .A3(_22787_),
    .A4(_22796_),
    .ZN(_22820_));
 INV_X1 _53836_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [165]),
    .ZN(_22821_));
 OAI21_X1 _53837_ (.A(_22820_),
    .B1(_22809_),
    .B2(_22821_),
    .ZN(_01554_));
 MUX2_X1 _53838_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [166]),
    .B(_10576_),
    .S(_22815_),
    .Z(_01565_));
 MUX2_X1 _53839_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [167]),
    .B(_10577_),
    .S(_22815_),
    .Z(_01576_));
 MUX2_X1 _53840_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [168]),
    .B(_10578_),
    .S(_22815_),
    .Z(_01587_));
 MUX2_X1 _53841_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [169]),
    .B(_10579_),
    .S(_22815_),
    .Z(_01598_));
 MUX2_X1 _53842_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [170]),
    .B(_22729_),
    .S(_22815_),
    .Z(_01610_));
 MUX2_X1 _53843_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [171]),
    .B(_10602_),
    .S(_22815_),
    .Z(_01621_));
 NAND4_X1 _53844_ (.A1(_10781_),
    .A2(_08594_),
    .A3(_22787_),
    .A4(_22796_),
    .ZN(_22822_));
 INV_X1 _53845_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [172]),
    .ZN(_22823_));
 OAI21_X1 _53846_ (.A(_22822_),
    .B1(_22809_),
    .B2(_22823_),
    .ZN(_01632_));
 MUX2_X1 _53847_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [173]),
    .B(_22680_),
    .S(_22815_),
    .Z(_01643_));
 MUX2_X1 _53848_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [174]),
    .B(_10584_),
    .S(_22815_),
    .Z(_01654_));
 MUX2_X1 _53849_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [175]),
    .B(_22681_),
    .S(_22815_),
    .Z(_01665_));
 BUF_X8 _53850_ (.A(_22807_),
    .Z(_22824_));
 MUX2_X1 _53851_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [176]),
    .B(_10586_),
    .S(_22824_),
    .Z(_01676_));
 MUX2_X1 _53852_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [177]),
    .B(_10587_),
    .S(_22824_),
    .Z(_01687_));
 MUX2_X1 _53853_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [178]),
    .B(_10588_),
    .S(_22824_),
    .Z(_01698_));
 MUX2_X1 _53854_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [179]),
    .B(_10603_),
    .S(_22824_),
    .Z(_01709_));
 MUX2_X1 _53855_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [180]),
    .B(_10604_),
    .S(_22824_),
    .Z(_01721_));
 MUX2_X1 _53856_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [181]),
    .B(_10591_),
    .S(_22824_),
    .Z(_01732_));
 MUX2_X1 _53857_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [182]),
    .B(_10592_),
    .S(_22824_),
    .Z(_01743_));
 MUX2_X1 _53858_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [183]),
    .B(_10593_),
    .S(_22824_),
    .Z(_01754_));
 MUX2_X1 _53859_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [184]),
    .B(_10605_),
    .S(_22824_),
    .Z(_01765_));
 MUX2_X1 _53860_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [185]),
    .B(_10595_),
    .S(_22824_),
    .Z(_01776_));
 MUX2_X1 _53861_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [186]),
    .B(_21595_),
    .S(_22808_),
    .Z(_01787_));
 MUX2_X1 _53862_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [187]),
    .B(_21763_),
    .S(_22808_),
    .Z(_01798_));
 MUX2_X1 _53863_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [188]),
    .B(_21407_),
    .S(_22808_),
    .Z(_01809_));
 NAND4_X1 _53864_ (.A1(_10781_),
    .A2(_22719_),
    .A3(_22774_),
    .A4(_21351_),
    .ZN(_22825_));
 INV_X1 _53865_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [189]),
    .ZN(_22826_));
 OAI21_X1 _53866_ (.A(_22825_),
    .B1(_22809_),
    .B2(_22826_),
    .ZN(_01820_));
 MUX2_X1 _53867_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [190]),
    .B(_21533_),
    .S(_22808_),
    .Z(_01832_));
 MUX2_X1 _53868_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [191]),
    .B(_21360_),
    .S(_22808_),
    .Z(_01843_));
 MUX2_X1 _53869_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [192]),
    .B(_22697_),
    .S(_22808_),
    .Z(_01854_));
 MUX2_X1 _53870_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [193]),
    .B(_22698_),
    .S(_22808_),
    .Z(_01865_));
 MUX2_X1 _53871_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [194]),
    .B(_22731_),
    .S(_22808_),
    .Z(_01876_));
 MUX2_X1 _53872_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [195]),
    .B(_22732_),
    .S(_22808_),
    .Z(_01887_));
 BUF_X16 _53873_ (.A(_11200_),
    .Z(_22827_));
 AND2_X4 _53874_ (.A1(_22827_),
    .A2(_10784_),
    .ZN(_22828_));
 BUF_X8 _53875_ (.A(_22828_),
    .Z(_22829_));
 MUX2_X1 _53876_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [98]),
    .B(_22685_),
    .S(_22829_),
    .Z(_03945_));
 MUX2_X1 _53877_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [99]),
    .B(_21605_),
    .S(_22829_),
    .Z(_03956_));
 BUF_X4 _53878_ (.A(_10784_),
    .Z(_22830_));
 NAND4_X1 _53879_ (.A1(_22716_),
    .A2(_21294_),
    .A3(_22830_),
    .A4(_22796_),
    .ZN(_22831_));
 BUF_X4 _53880_ (.A(_22829_),
    .Z(_22832_));
 INV_X1 _53881_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [100]),
    .ZN(_22833_));
 OAI21_X1 _53882_ (.A(_22831_),
    .B1(_22832_),
    .B2(_22833_),
    .ZN(_00833_));
 MUX2_X1 _53883_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [101]),
    .B(_21608_),
    .S(_22829_),
    .Z(_00844_));
 NAND4_X1 _53884_ (.A1(_22716_),
    .A2(_21297_),
    .A3(_22830_),
    .A4(_22796_),
    .ZN(_22834_));
 INV_X1 _53885_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [102]),
    .ZN(_22835_));
 OAI21_X1 _53886_ (.A(_22834_),
    .B1(_22832_),
    .B2(_22835_),
    .ZN(_00855_));
 MUX2_X1 _53887_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [103]),
    .B(_21299_),
    .S(_22829_),
    .Z(_00866_));
 MUX2_X1 _53888_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [104]),
    .B(_21578_),
    .S(_22829_),
    .Z(_00877_));
 MUX2_X1 _53889_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [105]),
    .B(_21582_),
    .S(_22829_),
    .Z(_00888_));
 BUF_X8 _53890_ (.A(_22828_),
    .Z(_22836_));
 MUX2_X1 _53891_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [106]),
    .B(_22705_),
    .S(_22836_),
    .Z(_00899_));
 BUF_X4 _53892_ (.A(_11177_),
    .Z(_22837_));
 NAND4_X1 _53893_ (.A1(_22716_),
    .A2(_21307_),
    .A3(_22830_),
    .A4(_22837_),
    .ZN(_22838_));
 INV_X1 _53894_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [107]),
    .ZN(_22839_));
 OAI21_X1 _53895_ (.A(_22838_),
    .B1(_22832_),
    .B2(_22839_),
    .ZN(_00910_));
 MUX2_X1 _53896_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [108]),
    .B(_21446_),
    .S(_22836_),
    .Z(_00921_));
 NAND4_X1 _53897_ (.A1(_22716_),
    .A2(_21311_),
    .A3(_22830_),
    .A4(_22837_),
    .ZN(_22840_));
 INV_X1 _53898_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [109]),
    .ZN(_22841_));
 OAI21_X1 _53899_ (.A(_22840_),
    .B1(_22832_),
    .B2(_22841_),
    .ZN(_00932_));
 MUX2_X1 _53900_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [110]),
    .B(_10563_),
    .S(_22836_),
    .Z(_00944_));
 MUX2_X1 _53901_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [111]),
    .B(_10569_),
    .S(_22836_),
    .Z(_00955_));
 NAND4_X1 _53902_ (.A1(_22716_),
    .A2(_08558_),
    .A3(_22830_),
    .A4(_22837_),
    .ZN(_22842_));
 INV_X2 _53903_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [112]),
    .ZN(_22843_));
 OAI21_X1 _53904_ (.A(_22842_),
    .B1(_22832_),
    .B2(_22843_),
    .ZN(_00966_));
 MUX2_X1 _53905_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [113]),
    .B(_10571_),
    .S(_22836_),
    .Z(_00977_));
 NAND4_X1 _53906_ (.A1(_22716_),
    .A2(_08564_),
    .A3(_22830_),
    .A4(_22837_),
    .ZN(_22844_));
 INV_X1 _53907_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [114]),
    .ZN(_22845_));
 OAI21_X1 _53908_ (.A(_22844_),
    .B1(_22832_),
    .B2(_22845_),
    .ZN(_00988_));
 NAND4_X1 _53909_ (.A1(_22716_),
    .A2(_08567_),
    .A3(_22830_),
    .A4(_22837_),
    .ZN(_22846_));
 INV_X1 _53910_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [115]),
    .ZN(_22847_));
 OAI21_X1 _53911_ (.A(_22846_),
    .B1(_22832_),
    .B2(_22847_),
    .ZN(_00999_));
 MUX2_X1 _53912_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [116]),
    .B(_10600_),
    .S(_22836_),
    .Z(_01010_));
 MUX2_X1 _53913_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [117]),
    .B(_10576_),
    .S(_22836_),
    .Z(_01021_));
 MUX2_X1 _53914_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [118]),
    .B(_10577_),
    .S(_22836_),
    .Z(_01032_));
 MUX2_X1 _53915_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [119]),
    .B(_10578_),
    .S(_22836_),
    .Z(_01043_));
 MUX2_X1 _53916_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [120]),
    .B(_10579_),
    .S(_22836_),
    .Z(_01055_));
 BUF_X16 _53917_ (.A(_22828_),
    .Z(_22848_));
 MUX2_X1 _53918_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [121]),
    .B(_22729_),
    .S(_22848_),
    .Z(_01066_));
 MUX2_X1 _53919_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [122]),
    .B(_10602_),
    .S(_22848_),
    .Z(_01077_));
 NAND4_X1 _53920_ (.A1(_22716_),
    .A2(_08594_),
    .A3(_22830_),
    .A4(_22837_),
    .ZN(_22849_));
 INV_X1 _53921_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [123]),
    .ZN(_22850_));
 OAI21_X1 _53922_ (.A(_22849_),
    .B1(_22832_),
    .B2(_22850_),
    .ZN(_01088_));
 MUX2_X1 _53923_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [124]),
    .B(_10583_),
    .S(_22848_),
    .Z(_01099_));
 MUX2_X1 _53924_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [125]),
    .B(_10584_),
    .S(_22848_),
    .Z(_01110_));
 MUX2_X1 _53925_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [126]),
    .B(_10585_),
    .S(_22848_),
    .Z(_01121_));
 MUX2_X1 _53926_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [127]),
    .B(_10586_),
    .S(_22848_),
    .Z(_01132_));
 MUX2_X1 _53927_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [128]),
    .B(_10587_),
    .S(_22848_),
    .Z(_01143_));
 MUX2_X1 _53928_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [129]),
    .B(_10588_),
    .S(_22848_),
    .Z(_01154_));
 MUX2_X1 _53929_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [130]),
    .B(_10603_),
    .S(_22848_),
    .Z(_01166_));
 MUX2_X1 _53930_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [131]),
    .B(_10604_),
    .S(_22848_),
    .Z(_01177_));
 NAND4_X1 _53931_ (.A1(_10859_),
    .A2(_08623_),
    .A3(_22830_),
    .A4(_22837_),
    .ZN(_22851_));
 INV_X1 _53932_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [132]),
    .ZN(_22852_));
 OAI21_X1 _53933_ (.A(_22851_),
    .B1(_22832_),
    .B2(_22852_),
    .ZN(_01188_));
 BUF_X16 _53934_ (.A(_22828_),
    .Z(_22853_));
 MUX2_X1 _53935_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [133]),
    .B(_10592_),
    .S(_22853_),
    .Z(_01199_));
 MUX2_X1 _53936_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [134]),
    .B(_10593_),
    .S(_22853_),
    .Z(_01210_));
 NAND4_X1 _53937_ (.A1(_10859_),
    .A2(_08632_),
    .A3(_22830_),
    .A4(_22837_),
    .ZN(_22854_));
 INV_X1 _53938_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [135]),
    .ZN(_22855_));
 OAI21_X1 _53939_ (.A(_22854_),
    .B1(_22832_),
    .B2(_22855_),
    .ZN(_01221_));
 MUX2_X1 _53940_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [136]),
    .B(_10595_),
    .S(_22853_),
    .Z(_01232_));
 MUX2_X1 _53941_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [137]),
    .B(_21595_),
    .S(_22853_),
    .Z(_01243_));
 MUX2_X1 _53942_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [138]),
    .B(_21763_),
    .S(_22853_),
    .Z(_01254_));
 NAND4_X1 _53943_ (.A1(_10859_),
    .A2(_22719_),
    .A3(_22774_),
    .A4(_21347_),
    .ZN(_22856_));
 INV_X1 _53944_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [139]),
    .ZN(_22857_));
 OAI21_X1 _53945_ (.A(_22856_),
    .B1(_22829_),
    .B2(_22857_),
    .ZN(_01265_));
 MUX2_X1 _53946_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [140]),
    .B(_21461_),
    .S(_22853_),
    .Z(_01277_));
 NAND4_X1 _53947_ (.A1(_10859_),
    .A2(_22719_),
    .A3(_22774_),
    .A4(_21355_),
    .ZN(_22858_));
 INV_X1 _53948_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [141]),
    .ZN(_22859_));
 OAI21_X1 _53949_ (.A(_22858_),
    .B1(_22829_),
    .B2(_22859_),
    .ZN(_01288_));
 MUX2_X1 _53950_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [142]),
    .B(_21360_),
    .S(_22853_),
    .Z(_01299_));
 MUX2_X1 _53951_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [143]),
    .B(_22697_),
    .S(_22853_),
    .Z(_01310_));
 NAND4_X1 _53952_ (.A1(_10859_),
    .A2(_22719_),
    .A3(_22774_),
    .A4(_21369_),
    .ZN(_22860_));
 INV_X1 _53953_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [144]),
    .ZN(_22861_));
 OAI21_X1 _53954_ (.A(_22860_),
    .B1(_22829_),
    .B2(_22861_),
    .ZN(_01321_));
 MUX2_X1 _53955_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [145]),
    .B(_22731_),
    .S(_22853_),
    .Z(_01332_));
 MUX2_X1 _53956_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [146]),
    .B(_22732_),
    .S(_22853_),
    .Z(_01343_));
 AND2_X4 _53957_ (.A1(_11205_),
    .A2(_21412_),
    .ZN(_22862_));
 BUF_X16 _53958_ (.A(_22862_),
    .Z(_22863_));
 BUF_X8 _53959_ (.A(_22863_),
    .Z(_22864_));
 MUX2_X1 _53960_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [0]),
    .B(_21598_),
    .S(_22864_),
    .Z(_00822_));
 MUX2_X1 _53961_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1]),
    .B(_21605_),
    .S(_22864_),
    .Z(_01933_));
 MUX2_X1 _53962_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2]),
    .B(_21383_),
    .S(_22864_),
    .Z(_03044_));
 MUX2_X1 _53963_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3]),
    .B(_21608_),
    .S(_22864_),
    .Z(_03291_));
 BUF_X16 _53964_ (.A(_22862_),
    .Z(_22865_));
 MUX2_X1 _53965_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [4]),
    .B(_21387_),
    .S(_22865_),
    .Z(_03402_));
 MUX2_X1 _53966_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [5]),
    .B(_21299_),
    .S(_22865_),
    .Z(_03513_));
 MUX2_X1 _53967_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [6]),
    .B(_21578_),
    .S(_22865_),
    .Z(_03624_));
 MUX2_X1 _53968_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [7]),
    .B(_21582_),
    .S(_22865_),
    .Z(_03735_));
 MUX2_X1 _53969_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [8]),
    .B(_22705_),
    .S(_22865_),
    .Z(_03846_));
 MUX2_X1 _53970_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [9]),
    .B(_21395_),
    .S(_22865_),
    .Z(_03957_));
 MUX2_X1 _53971_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [10]),
    .B(_21446_),
    .S(_22865_),
    .Z(_00933_));
 MUX2_X1 _53972_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [11]),
    .B(_21506_),
    .S(_22865_),
    .Z(_01044_));
 NAND4_X2 _53973_ (.A1(_22588_),
    .A2(_08551_),
    .A3(_10785_),
    .A4(_22837_),
    .ZN(_22866_));
 INV_X1 _53974_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [12]),
    .ZN(_22867_));
 OAI21_X1 _53975_ (.A(_22866_),
    .B1(_22864_),
    .B2(_22867_),
    .ZN(_01155_));
 MUX2_X1 _53976_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [13]),
    .B(_10569_),
    .S(_22865_),
    .Z(_01266_));
 NAND4_X1 _53977_ (.A1(_22588_),
    .A2(_08558_),
    .A3(_10785_),
    .A4(_22837_),
    .ZN(_22868_));
 INV_X1 _53978_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [14]),
    .ZN(_22869_));
 OAI21_X1 _53979_ (.A(_22868_),
    .B1(_22864_),
    .B2(_22869_),
    .ZN(_01377_));
 MUX2_X1 _53980_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [15]),
    .B(_10571_),
    .S(_22865_),
    .Z(_01488_));
 BUF_X16 _53981_ (.A(_22862_),
    .Z(_22870_));
 MUX2_X1 _53982_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [16]),
    .B(_10572_),
    .S(_22870_),
    .Z(_01599_));
 MUX2_X1 _53983_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [17]),
    .B(_10573_),
    .S(_22870_),
    .Z(_01710_));
 MUX2_X1 _53984_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [18]),
    .B(_10600_),
    .S(_22870_),
    .Z(_01821_));
 MUX2_X1 _53985_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [19]),
    .B(_10576_),
    .S(_22870_),
    .Z(_01932_));
 MUX2_X1 _53986_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [20]),
    .B(_10577_),
    .S(_22870_),
    .Z(_02044_));
 MUX2_X1 _53987_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [21]),
    .B(_10578_),
    .S(_22870_),
    .Z(_02155_));
 NAND4_X1 _53988_ (.A1(_22588_),
    .A2(_08584_),
    .A3(_10785_),
    .A4(_11177_),
    .ZN(_22871_));
 INV_X1 _53989_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [22]),
    .ZN(_22872_));
 OAI21_X1 _53990_ (.A(_22871_),
    .B1(_22864_),
    .B2(_22872_),
    .ZN(_02266_));
 MUX2_X1 _53991_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [23]),
    .B(_22729_),
    .S(_22870_),
    .Z(_02377_));
 MUX2_X1 _53992_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [24]),
    .B(_10602_),
    .S(_22870_),
    .Z(_02488_));
 MUX2_X1 _53993_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [25]),
    .B(_10582_),
    .S(_22870_),
    .Z(_02599_));
 MUX2_X1 _53994_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [26]),
    .B(_10583_),
    .S(_22870_),
    .Z(_02710_));
 BUF_X8 _53995_ (.A(_22862_),
    .Z(_22873_));
 MUX2_X1 _53996_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [27]),
    .B(_10584_),
    .S(_22873_),
    .Z(_02821_));
 NAND4_X2 _53997_ (.A1(_22588_),
    .A2(_08604_),
    .A3(_10785_),
    .A4(_11177_),
    .ZN(_22874_));
 INV_X1 _53998_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [28]),
    .ZN(_22875_));
 OAI21_X1 _53999_ (.A(_22874_),
    .B1(_22864_),
    .B2(_22875_),
    .ZN(_02932_));
 MUX2_X1 _54000_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [29]),
    .B(_10586_),
    .S(_22873_),
    .Z(_03043_));
 MUX2_X1 _54001_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [30]),
    .B(_10587_),
    .S(_22873_),
    .Z(_03155_));
 MUX2_X1 _54002_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [31]),
    .B(_10588_),
    .S(_22873_),
    .Z(_03202_));
 MUX2_X1 _54003_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [32]),
    .B(_10603_),
    .S(_22873_),
    .Z(_03213_));
 MUX2_X1 _54004_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [33]),
    .B(_10604_),
    .S(_22873_),
    .Z(_03224_));
 MUX2_X1 _54005_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [34]),
    .B(_10591_),
    .S(_22873_),
    .Z(_03235_));
 MUX2_X1 _54006_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [35]),
    .B(_10592_),
    .S(_22873_),
    .Z(_03246_));
 MUX2_X1 _54007_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [36]),
    .B(_10593_),
    .S(_22873_),
    .Z(_03257_));
 MUX2_X1 _54008_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [37]),
    .B(_10605_),
    .S(_22873_),
    .Z(_03268_));
 MUX2_X1 _54009_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [38]),
    .B(_10595_),
    .S(_22863_),
    .Z(_03279_));
 MUX2_X1 _54010_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [39]),
    .B(_21595_),
    .S(_22863_),
    .Z(_03290_));
 MUX2_X1 _54011_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [40]),
    .B(_21763_),
    .S(_22863_),
    .Z(_03302_));
 MUX2_X1 _54012_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [41]),
    .B(_21407_),
    .S(_22863_),
    .Z(_03313_));
 MUX2_X1 _54013_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [42]),
    .B(_21461_),
    .S(_22863_),
    .Z(_03324_));
 MUX2_X1 _54014_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [43]),
    .B(_21533_),
    .S(_22863_),
    .Z(_03335_));
 NAND4_X1 _54015_ (.A1(_22588_),
    .A2(_22719_),
    .A3(_22774_),
    .A4(_21359_),
    .ZN(_22876_));
 INV_X1 _54016_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [44]),
    .ZN(_22877_));
 OAI21_X1 _54017_ (.A(_22876_),
    .B1(_22864_),
    .B2(_22877_),
    .ZN(_03346_));
 MUX2_X1 _54018_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [45]),
    .B(_21365_),
    .S(_22863_),
    .Z(_03357_));
 NAND4_X1 _54019_ (.A1(_10880_),
    .A2(_21315_),
    .A3(_22774_),
    .A4(_21369_),
    .ZN(_22878_));
 INV_X1 _54020_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [46]),
    .ZN(_22879_));
 OAI21_X1 _54021_ (.A(_22878_),
    .B1(_22864_),
    .B2(_22879_),
    .ZN(_03368_));
 MUX2_X1 _54022_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [47]),
    .B(_22731_),
    .S(_22863_),
    .Z(_03379_));
 MUX2_X1 _54023_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [48]),
    .B(_22732_),
    .S(_22863_),
    .Z(_03390_));
 AND2_X4 _54024_ (.A1(_11211_),
    .A2(_21574_),
    .ZN(_22880_));
 BUF_X16 _54025_ (.A(_22880_),
    .Z(_22881_));
 BUF_X8 _54026_ (.A(_22881_),
    .Z(_22882_));
 MUX2_X1 _54027_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [49]),
    .B(_21598_),
    .S(_22882_),
    .Z(_03401_));
 MUX2_X1 _54028_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [50]),
    .B(_21605_),
    .S(_22882_),
    .Z(_03413_));
 NAND4_X1 _54029_ (.A1(_22563_),
    .A2(_21294_),
    .A3(_10785_),
    .A4(_11177_),
    .ZN(_22883_));
 INV_X1 _54030_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [51]),
    .ZN(_22884_));
 OAI21_X1 _54031_ (.A(_22883_),
    .B1(_22882_),
    .B2(_22884_),
    .ZN(_03424_));
 MUX2_X1 _54032_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [52]),
    .B(_21608_),
    .S(_22882_),
    .Z(_03435_));
 MUX2_X1 _54033_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [53]),
    .B(_21387_),
    .S(_22882_),
    .Z(_03446_));
 MUX2_X1 _54034_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [54]),
    .B(_21299_),
    .S(_22882_),
    .Z(_03457_));
 BUF_X16 _54035_ (.A(_22880_),
    .Z(_22885_));
 MUX2_X1 _54036_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [55]),
    .B(_21578_),
    .S(_22885_),
    .Z(_03468_));
 MUX2_X1 _54037_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [56]),
    .B(_21582_),
    .S(_22885_),
    .Z(_03479_));
 MUX2_X1 _54038_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [57]),
    .B(_21392_),
    .S(_22885_),
    .Z(_03490_));
 MUX2_X1 _54039_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [58]),
    .B(_21395_),
    .S(_22885_),
    .Z(_03501_));
 MUX2_X1 _54040_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [59]),
    .B(_21446_),
    .S(_22885_),
    .Z(_03512_));
 MUX2_X1 _54041_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [60]),
    .B(_21506_),
    .S(_22885_),
    .Z(_03524_));
 NAND4_X1 _54042_ (.A1(_22563_),
    .A2(_08551_),
    .A3(_10785_),
    .A4(_11177_),
    .ZN(_22886_));
 INV_X1 _54043_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [61]),
    .ZN(_22887_));
 OAI21_X1 _54044_ (.A(_22886_),
    .B1(_22882_),
    .B2(_22887_),
    .ZN(_03535_));
 MUX2_X1 _54045_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [62]),
    .B(_10569_),
    .S(_22885_),
    .Z(_03546_));
 MUX2_X1 _54046_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [63]),
    .B(_10570_),
    .S(_22885_),
    .Z(_03557_));
 MUX2_X1 _54047_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [64]),
    .B(_10571_),
    .S(_22885_),
    .Z(_03568_));
 MUX2_X1 _54048_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [65]),
    .B(_10572_),
    .S(_22885_),
    .Z(_03579_));
 BUF_X16 _54049_ (.A(_22880_),
    .Z(_22888_));
 MUX2_X1 _54050_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [66]),
    .B(_10573_),
    .S(_22888_),
    .Z(_03590_));
 MUX2_X1 _54051_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [67]),
    .B(_10600_),
    .S(_22888_),
    .Z(_03601_));
 MUX2_X1 _54052_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [68]),
    .B(_10576_),
    .S(_22888_),
    .Z(_03612_));
 MUX2_X1 _54053_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [69]),
    .B(_10577_),
    .S(_22888_),
    .Z(_03623_));
 MUX2_X1 _54054_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [70]),
    .B(_10578_),
    .S(_22888_),
    .Z(_03635_));
 MUX2_X1 _54055_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [71]),
    .B(_10579_),
    .S(_22888_),
    .Z(_03646_));
 MUX2_X1 _54056_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [72]),
    .B(_22729_),
    .S(_22888_),
    .Z(_03657_));
 MUX2_X1 _54057_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [73]),
    .B(_10602_),
    .S(_22888_),
    .Z(_03668_));
 MUX2_X1 _54058_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [74]),
    .B(_10582_),
    .S(_22888_),
    .Z(_03679_));
 MUX2_X1 _54059_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [75]),
    .B(_10583_),
    .S(_22888_),
    .Z(_03690_));
 BUF_X8 _54060_ (.A(_22880_),
    .Z(_22889_));
 MUX2_X1 _54061_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [76]),
    .B(_10584_),
    .S(_22889_),
    .Z(_03701_));
 MUX2_X1 _54062_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [77]),
    .B(_10585_),
    .S(_22889_),
    .Z(_03712_));
 MUX2_X1 _54063_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [78]),
    .B(_10586_),
    .S(_22889_),
    .Z(_03723_));
 MUX2_X1 _54064_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [79]),
    .B(_10587_),
    .S(_22889_),
    .Z(_03734_));
 MUX2_X1 _54065_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [80]),
    .B(_10588_),
    .S(_22889_),
    .Z(_03746_));
 MUX2_X1 _54066_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [81]),
    .B(_10603_),
    .S(_22889_),
    .Z(_03757_));
 MUX2_X1 _54067_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [82]),
    .B(_10604_),
    .S(_22889_),
    .Z(_03768_));
 NAND4_X1 _54068_ (.A1(_22563_),
    .A2(_08623_),
    .A3(_10785_),
    .A4(_11177_),
    .ZN(_22890_));
 INV_X1 _54069_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [83]),
    .ZN(_22891_));
 OAI21_X1 _54070_ (.A(_22890_),
    .B1(_22882_),
    .B2(_22891_),
    .ZN(_03779_));
 MUX2_X1 _54071_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [84]),
    .B(_10592_),
    .S(_22889_),
    .Z(_03790_));
 MUX2_X1 _54072_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [85]),
    .B(_10593_),
    .S(_22889_),
    .Z(_03801_));
 MUX2_X1 _54073_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [86]),
    .B(_10605_),
    .S(_22889_),
    .Z(_03812_));
 MUX2_X1 _54074_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [87]),
    .B(_10595_),
    .S(_22881_),
    .Z(_03823_));
 MUX2_X1 _54075_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [88]),
    .B(_21595_),
    .S(_22881_),
    .Z(_03834_));
 MUX2_X1 _54076_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [89]),
    .B(_21763_),
    .S(_22881_),
    .Z(_03845_));
 MUX2_X1 _54077_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [90]),
    .B(_21407_),
    .S(_22881_),
    .Z(_03857_));
 MUX2_X1 _54078_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [91]),
    .B(_21461_),
    .S(_22881_),
    .Z(_03868_));
 NAND4_X1 _54079_ (.A1(_22563_),
    .A2(_21315_),
    .A3(_22774_),
    .A4(_21355_),
    .ZN(_22892_));
 INV_X1 _54080_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [92]),
    .ZN(_22893_));
 OAI21_X1 _54081_ (.A(_22892_),
    .B1(_22882_),
    .B2(_22893_),
    .ZN(_03879_));
 NAND4_X1 _54082_ (.A1(_22563_),
    .A2(_21315_),
    .A3(_22774_),
    .A4(_21359_),
    .ZN(_22894_));
 INV_X1 _54083_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [93]),
    .ZN(_22895_));
 OAI21_X1 _54084_ (.A(_22894_),
    .B1(_22882_),
    .B2(_22895_),
    .ZN(_03890_));
 MUX2_X1 _54085_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [94]),
    .B(_21365_),
    .S(_22881_),
    .Z(_03901_));
 MUX2_X1 _54086_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [95]),
    .B(_22698_),
    .S(_22881_),
    .Z(_03912_));
 MUX2_X1 _54087_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [96]),
    .B(_22731_),
    .S(_22881_),
    .Z(_03923_));
 MUX2_X1 _54088_ (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [97]),
    .B(_22732_),
    .S(_22881_),
    .Z(_03934_));
 BUF_X32 _54089_ (.A(net91),
    .Z(_22896_));
 BUF_X32 _54090_ (.A(_22896_),
    .Z(_22897_));
 BUF_X8 _54091_ (.A(_11034_),
    .Z(_22898_));
 NAND3_X1 _54092_ (.A1(_22897_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1519]),
    .A3(_22898_),
    .ZN(_22899_));
 BUF_X32 _54093_ (.A(_10842_),
    .Z(_22900_));
 NAND3_X2 _54094_ (.A1(_22900_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1372]),
    .A3(_22898_),
    .ZN(_22901_));
 NAND2_X4 _54095_ (.A1(_22899_),
    .A2(_22901_),
    .ZN(_22902_));
 BUF_X16 _54096_ (.A(_11181_),
    .Z(_22903_));
 AOI221_X4 _54097_ (.A(_22902_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [686]),
    .B2(_11131_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [294]),
    .C2(_22903_),
    .ZN(_22904_));
 BUF_X16 _54098_ (.A(_11079_),
    .Z(_22905_));
 NAND3_X4 _54099_ (.A1(_22897_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1127]),
    .A3(_22905_),
    .ZN(_22906_));
 BUF_X32 _54100_ (.A(_10877_),
    .Z(_22907_));
 NAND3_X2 _54101_ (.A1(_22907_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1176]),
    .A3(_11035_),
    .ZN(_22908_));
 NAND2_X4 _54102_ (.A1(_22906_),
    .A2(_22908_),
    .ZN(_22909_));
 BUF_X16 _54103_ (.A(_10968_),
    .Z(_22910_));
 BUF_X16 _54104_ (.A(_21937_),
    .Z(_22911_));
 AOI221_X4 _54105_ (.A(_22909_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2058]),
    .B2(_22910_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2009]),
    .C2(_22911_),
    .ZN(_22912_));
 BUF_X16 _54106_ (.A(_10935_),
    .Z(_22913_));
 NAND3_X4 _54107_ (.A1(_22900_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2156]),
    .A3(_22913_),
    .ZN(_22914_));
 BUF_X32 _54108_ (.A(_10866_),
    .Z(_22915_));
 NAND3_X1 _54109_ (.A1(_22915_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [49]),
    .A3(_11174_),
    .ZN(_22916_));
 NAND2_X1 _54110_ (.A1(_22914_),
    .A2(_22916_),
    .ZN(_22917_));
 BUF_X16 _54111_ (.A(_10838_),
    .Z(_22918_));
 AOI221_X4 _54112_ (.A(_22917_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2940]),
    .B2(_22918_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [147]),
    .C2(_22806_),
    .ZN(_22919_));
 BUF_X32 _54113_ (.A(_10816_),
    .Z(_22920_));
 BUF_X8 _54114_ (.A(_10987_),
    .Z(_22921_));
 NAND3_X1 _54115_ (.A1(_22920_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1862]),
    .A3(_22921_),
    .ZN(_22922_));
 BUF_X16 _54116_ (.A(_10982_),
    .Z(_22923_));
 NAND3_X1 _54117_ (.A1(_10829_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1813]),
    .A3(_22923_),
    .ZN(_22924_));
 NAND2_X1 _54118_ (.A1(_22922_),
    .A2(_22924_),
    .ZN(_22925_));
 AOI221_X4 _54119_ (.A(_22925_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1617]),
    .B2(_11019_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1911]),
    .C2(_21978_),
    .ZN(_22926_));
 AND4_X1 _54120_ (.A1(_22904_),
    .A2(_22912_),
    .A3(_22919_),
    .A4(_22926_),
    .ZN(_22927_));
 BUF_X16 _54121_ (.A(_10825_),
    .Z(_22928_));
 AND4_X1 _54122_ (.A1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3038]),
    .A2(_10809_),
    .A3(_22928_),
    .A4(_10795_),
    .ZN(_22929_));
 AOI21_X4 _54123_ (.A(_22929_),
    .B1(_10800_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3087]),
    .ZN(_22930_));
 OAI221_X2 _54124_ (.A(_22930_),
    .B1(_22463_),
    .B2(_11096_),
    .C1(_22548_),
    .C2(_11111_),
    .ZN(_22931_));
 BUF_X32 _54125_ (.A(_22900_),
    .Z(_22932_));
 BUF_X16 _54126_ (.A(_22932_),
    .Z(_22933_));
 BUF_X8 _54127_ (.A(_10987_),
    .Z(_22934_));
 BUF_X8 _54128_ (.A(_22934_),
    .Z(_22935_));
 NAND3_X4 _54129_ (.A1(_22933_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1764]),
    .A3(_22935_),
    .ZN(_22936_));
 BUF_X16 _54130_ (.A(_11185_),
    .Z(_22937_));
 BUF_X16 _54131_ (.A(_22937_),
    .Z(_22938_));
 BUF_X8 _54132_ (.A(_22938_),
    .Z(_22939_));
 BUF_X8 _54133_ (.A(_22939_),
    .Z(_22940_));
 NAND3_X2 _54134_ (.A1(_22933_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [196]),
    .A3(_22940_),
    .ZN(_22941_));
 BUF_X32 _54135_ (.A(_10816_),
    .Z(_22942_));
 BUF_X32 _54136_ (.A(_22942_),
    .Z(_22943_));
 BUF_X16 _54137_ (.A(_22943_),
    .Z(_22944_));
 BUF_X16 _54138_ (.A(_11036_),
    .Z(_22945_));
 NAND3_X4 _54139_ (.A1(_22944_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1470]),
    .A3(_22945_),
    .ZN(_22946_));
 NAND3_X1 _54140_ (.A1(_10858_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [98]),
    .A3(_11176_),
    .ZN(_22947_));
 NAND4_X2 _54141_ (.A1(_22936_),
    .A2(_22941_),
    .A3(_22946_),
    .A4(_22947_),
    .ZN(_22948_));
 BUF_X32 _54142_ (.A(_22897_),
    .Z(_22949_));
 BUF_X16 _54143_ (.A(_22949_),
    .Z(_22950_));
 BUF_X8 _54144_ (.A(_11175_),
    .Z(_22951_));
 NAND3_X2 _54145_ (.A1(_22950_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [343]),
    .A3(_22951_),
    .ZN(_22952_));
 BUF_X32 _54146_ (.A(_10778_),
    .Z(_22953_));
 BUF_X32 _54147_ (.A(_22953_),
    .Z(_22954_));
 BUF_X16 _54148_ (.A(_22954_),
    .Z(_22955_));
 BUF_X16 _54149_ (.A(_22934_),
    .Z(_22956_));
 NAND3_X4 _54150_ (.A1(_22955_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1715]),
    .A3(_22956_),
    .ZN(_22957_));
 BUF_X16 _54151_ (.A(_10830_),
    .Z(_22958_));
 BUF_X8 _54152_ (.A(_11175_),
    .Z(_22959_));
 NAND3_X1 _54153_ (.A1(_22958_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [245]),
    .A3(_22959_),
    .ZN(_22960_));
 BUF_X16 _54154_ (.A(_22943_),
    .Z(_22961_));
 BUF_X16 _54155_ (.A(_10935_),
    .Z(_22962_));
 BUF_X8 _54156_ (.A(_22962_),
    .Z(_22963_));
 BUF_X8 _54157_ (.A(_22963_),
    .Z(_22964_));
 NAND3_X4 _54158_ (.A1(_22961_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2254]),
    .A3(_22964_),
    .ZN(_22965_));
 NAND4_X2 _54159_ (.A1(_22952_),
    .A2(_22957_),
    .A3(_22960_),
    .A4(_22965_),
    .ZN(_22966_));
 BUF_X32 _54160_ (.A(_22907_),
    .Z(_22967_));
 BUF_X16 _54161_ (.A(_22967_),
    .Z(_22968_));
 BUF_X16 _54162_ (.A(_22905_),
    .Z(_22969_));
 BUF_X8 _54163_ (.A(_22969_),
    .Z(_22970_));
 NAND3_X2 _54164_ (.A1(_22968_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [784]),
    .A3(_22970_),
    .ZN(_22971_));
 BUF_X16 _54165_ (.A(_22943_),
    .Z(_22972_));
 BUF_X8 _54166_ (.A(_22969_),
    .Z(_22973_));
 NAND3_X1 _54167_ (.A1(_22972_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1078]),
    .A3(_22973_),
    .ZN(_22974_));
 BUF_X16 _54168_ (.A(_10830_),
    .Z(_22975_));
 BUF_X8 _54169_ (.A(_22969_),
    .Z(_22976_));
 NAND3_X1 _54170_ (.A1(_22975_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1029]),
    .A3(_22976_),
    .ZN(_22977_));
 BUF_X16 _54171_ (.A(_10830_),
    .Z(_22978_));
 BUF_X8 _54172_ (.A(_11034_),
    .Z(_22979_));
 BUF_X8 _54173_ (.A(_22979_),
    .Z(_22980_));
 BUF_X8 _54174_ (.A(_22980_),
    .Z(_22981_));
 NAND3_X4 _54175_ (.A1(_22978_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1421]),
    .A3(_22981_),
    .ZN(_22982_));
 NAND4_X4 _54176_ (.A1(_22971_),
    .A2(_22974_),
    .A3(_22977_),
    .A4(_22982_),
    .ZN(_22983_));
 NOR4_X2 _54177_ (.A1(_22931_),
    .A2(_22948_),
    .A3(_22966_),
    .A4(_22983_),
    .ZN(_22984_));
 BUF_X16 _54178_ (.A(_10780_),
    .Z(_22985_));
 NAND3_X4 _54179_ (.A1(_22985_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [539]),
    .A3(_11127_),
    .ZN(_22986_));
 BUF_X32 _54180_ (.A(_10779_),
    .Z(_22987_));
 BUF_X16 _54181_ (.A(_22987_),
    .Z(_22988_));
 BUF_X16 _54182_ (.A(_10787_),
    .Z(_22989_));
 BUF_X8 _54183_ (.A(_22989_),
    .Z(_22990_));
 BUF_X8 _54184_ (.A(_22990_),
    .Z(_22991_));
 NAND3_X4 _54185_ (.A1(_22988_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2891]),
    .A3(_22991_),
    .ZN(_22992_));
 BUF_X32 _54186_ (.A(_10878_),
    .Z(_22993_));
 BUF_X32 _54187_ (.A(_22993_),
    .Z(_22994_));
 BUF_X8 _54188_ (.A(_11126_),
    .Z(_22995_));
 NAND3_X4 _54189_ (.A1(_22994_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [392]),
    .A3(_22995_),
    .ZN(_22996_));
 BUF_X32 _54190_ (.A(_22240_),
    .Z(_22997_));
 BUF_X16 _54191_ (.A(_22997_),
    .Z(_22998_));
 BUF_X16 _54192_ (.A(_22989_),
    .Z(_22999_));
 BUF_X16 _54193_ (.A(_22999_),
    .Z(_23000_));
 NAND3_X4 _54194_ (.A1(_22998_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2989]),
    .A3(_23000_),
    .ZN(_23001_));
 NAND4_X4 _54195_ (.A1(_22986_),
    .A2(_22992_),
    .A3(_22996_),
    .A4(_23001_),
    .ZN(_23002_));
 BUF_X32 _54196_ (.A(_10779_),
    .Z(_23003_));
 BUF_X16 _54197_ (.A(_23003_),
    .Z(_23004_));
 BUF_X8 _54198_ (.A(_10940_),
    .Z(_23005_));
 BUF_X8 _54199_ (.A(_23005_),
    .Z(_23006_));
 NAND3_X1 _54200_ (.A1(_23004_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2107]),
    .A3(_23006_),
    .ZN(_23007_));
 BUF_X16 _54201_ (.A(_22967_),
    .Z(_23008_));
 BUF_X8 _54202_ (.A(_22934_),
    .Z(_23009_));
 NAND3_X2 _54203_ (.A1(_23008_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1568]),
    .A3(_23009_),
    .ZN(_23010_));
 BUF_X32 _54204_ (.A(_22932_),
    .Z(_23011_));
 BUF_X8 _54205_ (.A(_10890_),
    .Z(_23012_));
 BUF_X8 _54206_ (.A(_23012_),
    .Z(_23013_));
 BUF_X8 _54207_ (.A(_23013_),
    .Z(_23014_));
 NAND3_X4 _54208_ (.A1(_23011_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2548]),
    .A3(_23014_),
    .ZN(_23015_));
 BUF_X32 _54209_ (.A(_10857_),
    .Z(_23016_));
 NAND3_X2 _54210_ (.A1(_23016_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1666]),
    .A3(_22956_),
    .ZN(_23017_));
 NAND4_X4 _54211_ (.A1(_23007_),
    .A2(_23010_),
    .A3(_23015_),
    .A4(_23017_),
    .ZN(_23018_));
 BUF_X32 _54212_ (.A(_10779_),
    .Z(_23019_));
 BUF_X16 _54213_ (.A(_23019_),
    .Z(_23020_));
 NAND3_X1 _54214_ (.A1(_23020_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2499]),
    .A3(_23014_),
    .ZN(_23021_));
 BUF_X16 _54215_ (.A(_22967_),
    .Z(_23022_));
 BUF_X8 _54216_ (.A(_23013_),
    .Z(_23023_));
 NAND3_X2 _54217_ (.A1(_23022_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2352]),
    .A3(_23023_),
    .ZN(_23024_));
 BUF_X16 _54218_ (.A(_10857_),
    .Z(_23025_));
 BUF_X8 _54219_ (.A(_23013_),
    .Z(_23026_));
 NAND3_X2 _54220_ (.A1(_23025_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2450]),
    .A3(_23026_),
    .ZN(_23027_));
 BUF_X16 _54221_ (.A(_10817_),
    .Z(_23028_));
 BUF_X8 _54222_ (.A(_23013_),
    .Z(_23029_));
 NAND3_X2 _54223_ (.A1(_23028_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2646]),
    .A3(_23029_),
    .ZN(_23030_));
 NAND4_X4 _54224_ (.A1(_23021_),
    .A2(_23024_),
    .A3(_23027_),
    .A4(_23030_),
    .ZN(_23031_));
 BUF_X16 _54225_ (.A(_22967_),
    .Z(_23032_));
 BUF_X8 _54226_ (.A(_10789_),
    .Z(_23033_));
 NAND3_X2 _54227_ (.A1(_23032_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2744]),
    .A3(_23033_),
    .ZN(_23034_));
 BUF_X32 _54228_ (.A(_22915_),
    .Z(_23035_));
 BUF_X16 _54229_ (.A(_23035_),
    .Z(_23036_));
 BUF_X8 _54230_ (.A(_22928_),
    .Z(_23037_));
 NAND3_X2 _54231_ (.A1(_23036_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2793]),
    .A3(_23037_),
    .ZN(_23038_));
 BUF_X16 _54232_ (.A(_10857_),
    .Z(_23039_));
 NAND3_X1 _54233_ (.A1(_23039_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2842]),
    .A3(_23037_),
    .ZN(_23040_));
 BUF_X32 _54234_ (.A(_10866_),
    .Z(_23041_));
 BUF_X16 _54235_ (.A(_23041_),
    .Z(_23042_));
 BUF_X16 _54236_ (.A(_10891_),
    .Z(_23043_));
 NAND3_X4 _54237_ (.A1(_23042_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2401]),
    .A3(_23043_),
    .ZN(_23044_));
 NAND4_X4 _54238_ (.A1(_23034_),
    .A2(_23038_),
    .A3(_23040_),
    .A4(_23044_),
    .ZN(_23045_));
 NOR4_X4 _54239_ (.A1(_23002_),
    .A2(_23018_),
    .A3(_23031_),
    .A4(_23045_),
    .ZN(_23046_));
 BUF_X16 _54240_ (.A(_11100_),
    .Z(_23047_));
 BUF_X16 _54241_ (.A(_11065_),
    .Z(_23048_));
 AOI22_X4 _54242_ (.A1(_23047_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [931]),
    .B1(_23048_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1225]),
    .ZN(_23049_));
 BUF_X8 _54243_ (.A(_22898_),
    .Z(_23050_));
 BUF_X16 _54244_ (.A(_23050_),
    .Z(_23051_));
 NAND3_X2 _54245_ (.A1(_10858_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1274]),
    .A3(_23051_),
    .ZN(_23052_));
 OAI211_X4 _54246_ (.A(_23049_),
    .B(_23052_),
    .C1(_22286_),
    .C2(_11055_),
    .ZN(_23053_));
 BUF_X16 _54247_ (.A(_22949_),
    .Z(_23054_));
 BUF_X8 _54248_ (.A(_11124_),
    .Z(_23055_));
 BUF_X16 _54249_ (.A(_23055_),
    .Z(_23056_));
 BUF_X8 _54250_ (.A(_23056_),
    .Z(_23057_));
 NAND3_X1 _54251_ (.A1(_23054_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [735]),
    .A3(_23057_),
    .ZN(_23058_));
 BUF_X16 _54252_ (.A(_22932_),
    .Z(_23059_));
 BUF_X8 _54253_ (.A(_23056_),
    .Z(_23060_));
 NAND3_X2 _54254_ (.A1(_23059_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [588]),
    .A3(_23060_),
    .ZN(_23061_));
 BUF_X16 _54255_ (.A(_23035_),
    .Z(_23062_));
 BUF_X8 _54256_ (.A(_23056_),
    .Z(_23063_));
 NAND3_X2 _54257_ (.A1(_23062_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [441]),
    .A3(_23063_),
    .ZN(_23064_));
 NAND3_X2 _54258_ (.A1(_23016_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [882]),
    .A3(_22970_),
    .ZN(_23065_));
 NAND4_X4 _54259_ (.A1(_23058_),
    .A2(_23061_),
    .A3(_23064_),
    .A4(_23065_),
    .ZN(_23066_));
 BUF_X16 _54260_ (.A(_22949_),
    .Z(_23067_));
 BUF_X8 _54261_ (.A(_23013_),
    .Z(_23068_));
 NAND3_X1 _54262_ (.A1(_23067_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2695]),
    .A3(_23068_),
    .ZN(_23069_));
 NAND3_X4 _54263_ (.A1(_23022_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1960]),
    .A3(_22964_),
    .ZN(_23070_));
 BUF_X16 _54264_ (.A(_10830_),
    .Z(_23071_));
 BUF_X8 _54265_ (.A(_11125_),
    .Z(_23072_));
 NAND3_X4 _54266_ (.A1(_23071_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [637]),
    .A3(_23072_),
    .ZN(_23073_));
 NAND3_X1 _54267_ (.A1(_22978_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2597]),
    .A3(_23043_),
    .ZN(_23074_));
 NAND4_X2 _54268_ (.A1(_23069_),
    .A2(_23070_),
    .A3(_23073_),
    .A4(_23074_),
    .ZN(_23075_));
 BUF_X16 _54269_ (.A(_22949_),
    .Z(_23076_));
 NAND3_X4 _54270_ (.A1(_23076_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2303]),
    .A3(_22964_),
    .ZN(_23077_));
 BUF_X16 _54271_ (.A(_10857_),
    .Z(_23078_));
 NAND3_X4 _54272_ (.A1(_23078_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [490]),
    .A3(_23072_),
    .ZN(_23079_));
 BUF_X16 _54273_ (.A(_10830_),
    .Z(_23080_));
 BUF_X8 _54274_ (.A(_22963_),
    .Z(_23081_));
 NAND3_X4 _54275_ (.A1(_23080_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2205]),
    .A3(_23081_),
    .ZN(_23082_));
 BUF_X32 _54276_ (.A(_10873_),
    .Z(_23083_));
 BUF_X32 _54277_ (.A(_23083_),
    .Z(_23084_));
 BUF_X16 _54278_ (.A(_23084_),
    .Z(_23085_));
 BUF_X8 _54279_ (.A(_22938_),
    .Z(_23086_));
 NAND3_X1 _54280_ (.A1(_23085_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [0]),
    .A3(_23086_),
    .ZN(_23087_));
 NAND4_X1 _54281_ (.A1(_23077_),
    .A2(_23079_),
    .A3(_23082_),
    .A4(_23087_),
    .ZN(_23088_));
 NOR4_X1 _54282_ (.A1(_23053_),
    .A2(_23066_),
    .A3(_23075_),
    .A4(_23088_),
    .ZN(_23089_));
 NAND4_X1 _54283_ (.A1(_22927_),
    .A2(_22984_),
    .A3(_23046_),
    .A4(_23089_),
    .ZN(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [0]));
 AND3_X1 _54284_ (.A1(_10803_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1912]),
    .A3(_10988_),
    .ZN(_23090_));
 AOI21_X4 _54285_ (.A(_23090_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1863]),
    .B2(_22003_),
    .ZN(_23091_));
 BUF_X32 _54286_ (.A(_11131_),
    .Z(_23092_));
 AOI22_X4 _54287_ (.A1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [687]),
    .A2(_23092_),
    .B1(_22827_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [99]),
    .ZN(_23093_));
 BUF_X16 _54288_ (.A(_11050_),
    .Z(_23094_));
 BUF_X8 _54289_ (.A(_11041_),
    .Z(_23095_));
 AOI22_X4 _54290_ (.A1(_23094_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1373]),
    .B1(_23095_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1471]),
    .ZN(_23096_));
 BUF_X16 _54291_ (.A(_10936_),
    .Z(_23097_));
 AOI22_X4 _54292_ (.A1(_23097_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2304]),
    .B1(_10976_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1961]),
    .ZN(_23098_));
 AND4_X4 _54293_ (.A1(_23091_),
    .A2(_23093_),
    .A3(_23096_),
    .A4(_23098_),
    .ZN(_23099_));
 AND3_X1 _54294_ (.A1(_22896_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1128]),
    .A3(_11079_),
    .ZN(_23100_));
 AND3_X1 _54295_ (.A1(_10816_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1079]),
    .A3(_11079_),
    .ZN(_23101_));
 OR2_X1 _54296_ (.A1(_23100_),
    .A2(_23101_),
    .ZN(_23102_));
 BUF_X16 _54297_ (.A(_11069_),
    .Z(_23103_));
 BUF_X16 _54298_ (.A(_11094_),
    .Z(_23104_));
 AOI221_X2 _54299_ (.A(_23102_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1177]),
    .B2(_23103_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [981]),
    .C2(_23104_),
    .ZN(_23105_));
 BUF_X16 _54300_ (.A(_11141_),
    .Z(_23106_));
 BUF_X16 _54301_ (.A(_11136_),
    .Z(_23107_));
 AOI22_X4 _54302_ (.A1(_23106_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [589]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [638]),
    .B2(_23107_),
    .ZN(_23108_));
 AOI22_X4 _54303_ (.A1(_10839_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2941]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2990]),
    .B2(_10826_),
    .ZN(_23109_));
 AND4_X1 _54304_ (.A1(_23099_),
    .A2(net56),
    .A3(_23108_),
    .A4(_23109_),
    .ZN(_23110_));
 NAND3_X2 _54305_ (.A1(_22985_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1324]),
    .A3(_23051_),
    .ZN(_23111_));
 NAND3_X4 _54306_ (.A1(_22988_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1716]),
    .A3(_10990_),
    .ZN(_23112_));
 BUF_X32 _54307_ (.A(_10867_),
    .Z(_23113_));
 BUF_X32 _54308_ (.A(_23113_),
    .Z(_23114_));
 NAND3_X4 _54309_ (.A1(_23114_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1226]),
    .A3(_23051_),
    .ZN(_23115_));
 BUF_X8 _54310_ (.A(_10989_),
    .Z(_23116_));
 NAND3_X2 _54311_ (.A1(_22998_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1814]),
    .A3(_23116_),
    .ZN(_23117_));
 NAND4_X4 _54312_ (.A1(_23111_),
    .A2(_23112_),
    .A3(_23115_),
    .A4(_23117_),
    .ZN(_23118_));
 BUF_X8 _54313_ (.A(_10891_),
    .Z(_23119_));
 BUF_X8 _54314_ (.A(_23119_),
    .Z(_23120_));
 NAND3_X4 _54315_ (.A1(_23004_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2500]),
    .A3(_23120_),
    .ZN(_23121_));
 BUF_X8 _54316_ (.A(_10788_),
    .Z(_23122_));
 BUF_X16 _54317_ (.A(_23122_),
    .Z(_23123_));
 NAND3_X4 _54318_ (.A1(_22950_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3088]),
    .A3(_23123_),
    .ZN(_23124_));
 BUF_X16 _54319_ (.A(_23019_),
    .Z(_23125_));
 NAND3_X1 _54320_ (.A1(_23125_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2892]),
    .A3(_23123_),
    .ZN(_23126_));
 BUF_X16 _54321_ (.A(_22943_),
    .Z(_23127_));
 BUF_X16 _54322_ (.A(_10789_),
    .Z(_23128_));
 NAND3_X2 _54323_ (.A1(_23127_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3039]),
    .A3(_23128_),
    .ZN(_23129_));
 NAND4_X4 _54324_ (.A1(_23121_),
    .A2(_23124_),
    .A3(_23126_),
    .A4(_23129_),
    .ZN(_23130_));
 BUF_X8 _54325_ (.A(_23013_),
    .Z(_23131_));
 NAND3_X2 _54326_ (.A1(_22950_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2696]),
    .A3(_23131_),
    .ZN(_23132_));
 BUF_X16 _54327_ (.A(_22967_),
    .Z(_23133_));
 BUF_X8 _54328_ (.A(_23013_),
    .Z(_23134_));
 NAND3_X2 _54329_ (.A1(_23133_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2353]),
    .A3(_23134_),
    .ZN(_23135_));
 NAND3_X2 _54330_ (.A1(_22958_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2598]),
    .A3(_23023_),
    .ZN(_23136_));
 NAND3_X2 _54331_ (.A1(_23025_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2451]),
    .A3(_23026_),
    .ZN(_23137_));
 NAND4_X4 _54332_ (.A1(_23132_),
    .A2(_23135_),
    .A3(_23136_),
    .A4(_23137_),
    .ZN(_23138_));
 NAND3_X2 _54333_ (.A1(_22968_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1569]),
    .A3(_22956_),
    .ZN(_23139_));
 BUF_X8 _54334_ (.A(_10857_),
    .Z(_23140_));
 BUF_X8 _54335_ (.A(_22934_),
    .Z(_23141_));
 NAND3_X2 _54336_ (.A1(_23140_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1667]),
    .A3(_23141_),
    .ZN(_23142_));
 BUF_X8 _54337_ (.A(_23013_),
    .Z(_23143_));
 NAND3_X4 _54338_ (.A1(_22961_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2647]),
    .A3(_23143_),
    .ZN(_23144_));
 BUF_X16 _54339_ (.A(_23035_),
    .Z(_23145_));
 BUF_X16 _54340_ (.A(_22934_),
    .Z(_23146_));
 NAND3_X2 _54341_ (.A1(_23145_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1618]),
    .A3(_23146_),
    .ZN(_23147_));
 NAND4_X4 _54342_ (.A1(_23139_),
    .A2(_23142_),
    .A3(_23144_),
    .A4(_23147_),
    .ZN(_23148_));
 NOR4_X4 _54343_ (.A1(_23118_),
    .A2(_23130_),
    .A3(_23138_),
    .A4(_23148_),
    .ZN(_23149_));
 BUF_X32 _54344_ (.A(_22896_),
    .Z(_23150_));
 BUF_X16 _54345_ (.A(_11145_),
    .Z(_23151_));
 NAND3_X4 _54346_ (.A1(_23150_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [736]),
    .A3(_23151_),
    .ZN(_23152_));
 BUF_X32 _54347_ (.A(_10842_),
    .Z(_23153_));
 NAND3_X2 _54348_ (.A1(_23153_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [197]),
    .A3(_11174_),
    .ZN(_23154_));
 NAND2_X4 _54349_ (.A1(_23152_),
    .A2(_23154_),
    .ZN(_23155_));
 BUF_X16 _54350_ (.A(_21937_),
    .Z(_23156_));
 AOI221_X1 _54351_ (.A(_23155_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2059]),
    .B2(_22910_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2010]),
    .C2(_23156_),
    .ZN(_23157_));
 BUF_X32 _54352_ (.A(_10778_),
    .Z(_23158_));
 BUF_X8 _54353_ (.A(_11173_),
    .Z(_23159_));
 NAND3_X2 _54354_ (.A1(_23158_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [148]),
    .A3(_23159_),
    .ZN(_23160_));
 BUF_X16 _54355_ (.A(_11145_),
    .Z(_23161_));
 NAND3_X4 _54356_ (.A1(_10856_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [491]),
    .A3(_23161_),
    .ZN(_23162_));
 NAND2_X4 _54357_ (.A1(_23160_),
    .A2(_23162_),
    .ZN(_23163_));
 BUF_X16 _54358_ (.A(_11205_),
    .Z(_23164_));
 AOI221_X2 _54359_ (.A(_23163_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1765]),
    .B2(_11002_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1]),
    .C2(_23164_),
    .ZN(_23165_));
 BUF_X32 _54360_ (.A(_10757_),
    .Z(_23166_));
 NAND3_X1 _54361_ (.A1(_23166_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2108]),
    .A3(_22962_),
    .ZN(_23167_));
 BUF_X32 _54362_ (.A(_10901_),
    .Z(_23168_));
 BUF_X8 _54363_ (.A(_10935_),
    .Z(_23169_));
 NAND3_X1 _54364_ (.A1(_23168_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2206]),
    .A3(_23169_),
    .ZN(_23170_));
 NAND2_X1 _54365_ (.A1(_23167_),
    .A2(_23170_),
    .ZN(_23171_));
 AOI221_X4 _54366_ (.A(_23171_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2255]),
    .B2(_21816_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2157]),
    .C2(_10955_),
    .ZN(_23172_));
 BUF_X32 _54367_ (.A(_10855_),
    .Z(_23173_));
 BUF_X8 _54368_ (.A(net107),
    .Z(_23174_));
 NAND3_X1 _54369_ (.A1(_23173_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2843]),
    .A3(_23174_),
    .ZN(_23175_));
 BUF_X32 _54370_ (.A(_10920_),
    .Z(_23176_));
 NAND3_X2 _54371_ (.A1(_23176_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2794]),
    .A3(_10825_),
    .ZN(_23177_));
 NAND2_X4 _54372_ (.A1(_23175_),
    .A2(_23177_),
    .ZN(_23178_));
 BUF_X8 _54373_ (.A(_11031_),
    .Z(_23179_));
 AOI221_X4 _54374_ (.A(_23178_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1422]),
    .B2(_22232_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1520]),
    .C2(_23179_),
    .ZN(_23180_));
 AND4_X2 _54375_ (.A1(_23157_),
    .A2(_23165_),
    .A3(_23172_),
    .A4(_23180_),
    .ZN(_23181_));
 AND3_X1 _54376_ (.A1(_22522_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [883]),
    .A3(_11080_),
    .ZN(_23182_));
 AOI21_X2 _54377_ (.A(_23182_),
    .B1(_23047_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [932]),
    .ZN(_23183_));
 OAI221_X2 _54378_ (.A(_23183_),
    .B1(_22440_),
    .B2(_11091_),
    .C1(_22578_),
    .C2(_11115_),
    .ZN(_23184_));
 NAND3_X1 _54379_ (.A1(_23054_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [344]),
    .A3(_22940_),
    .ZN(_23185_));
 NAND3_X2 _54380_ (.A1(_10831_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [246]),
    .A3(_22951_),
    .ZN(_23186_));
 BUF_X16 _54381_ (.A(_11175_),
    .Z(_23187_));
 NAND3_X2 _54382_ (.A1(_23062_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [50]),
    .A3(_23187_),
    .ZN(_23188_));
 BUF_X16 _54383_ (.A(_23035_),
    .Z(_23189_));
 NAND3_X4 _54384_ (.A1(_23189_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [834]),
    .A3(_22970_),
    .ZN(_23190_));
 NAND4_X4 _54385_ (.A1(_23185_),
    .A2(_23186_),
    .A3(_23188_),
    .A4(_23190_),
    .ZN(_23191_));
 BUF_X16 _54386_ (.A(_10843_),
    .Z(_23192_));
 NAND3_X2 _54387_ (.A1(_23192_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2549]),
    .A3(_23068_),
    .ZN(_23193_));
 BUF_X8 _54388_ (.A(_23084_),
    .Z(_23194_));
 NAND3_X2 _54389_ (.A1(_23194_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2745]),
    .A3(_10790_),
    .ZN(_23195_));
 BUF_X8 _54390_ (.A(_11175_),
    .Z(_23196_));
 NAND3_X4 _54391_ (.A1(_22961_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [295]),
    .A3(_23196_),
    .ZN(_23197_));
 NAND3_X2 _54392_ (.A1(_23145_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2402]),
    .A3(_23043_),
    .ZN(_23198_));
 NAND4_X4 _54393_ (.A1(_23193_),
    .A2(_23195_),
    .A3(_23197_),
    .A4(_23198_),
    .ZN(_23199_));
 BUF_X16 _54394_ (.A(_22954_),
    .Z(_23200_));
 BUF_X16 _54395_ (.A(_11125_),
    .Z(_23201_));
 NAND3_X2 _54396_ (.A1(_23200_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [540]),
    .A3(_23201_),
    .ZN(_23202_));
 NAND3_X1 _54397_ (.A1(_23145_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [442]),
    .A3(_23072_),
    .ZN(_23203_));
 BUF_X32 _54398_ (.A(_22522_),
    .Z(_23204_));
 BUF_X8 _54399_ (.A(_22980_),
    .Z(_23205_));
 NAND3_X4 _54400_ (.A1(_23204_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1275]),
    .A3(_23205_),
    .ZN(_23206_));
 BUF_X32 _54401_ (.A(_10878_),
    .Z(_23207_));
 BUF_X8 _54402_ (.A(_11125_),
    .Z(_23208_));
 NAND3_X2 _54403_ (.A1(_23207_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [393]),
    .A3(_23208_),
    .ZN(_23209_));
 NAND4_X4 _54404_ (.A1(_23202_),
    .A2(_23203_),
    .A3(_23206_),
    .A4(_23209_),
    .ZN(_23210_));
 NOR4_X4 _54405_ (.A1(_23184_),
    .A2(_23191_),
    .A3(_23199_),
    .A4(_23210_),
    .ZN(_23211_));
 NAND4_X1 _54406_ (.A1(_23110_),
    .A2(_23149_),
    .A3(_23181_),
    .A4(_23211_),
    .ZN(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [1]));
 AND3_X1 _54407_ (.A1(_10867_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2795]),
    .A3(_10788_),
    .ZN(_23212_));
 BUF_X8 _54408_ (.A(_10773_),
    .Z(_23213_));
 AOI221_X4 _54409_ (.A(_23212_),
    .B1(_21502_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2844]),
    .C1(_23213_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2893]),
    .ZN(_23214_));
 BUF_X32 _54410_ (.A(_10901_),
    .Z(_23215_));
 NAND3_X2 _54411_ (.A1(_23215_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2207]),
    .A3(_23169_),
    .ZN(_23216_));
 BUF_X32 _54412_ (.A(_10797_),
    .Z(_23217_));
 NAND3_X2 _54413_ (.A1(_23217_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2305]),
    .A3(_10939_),
    .ZN(_23218_));
 OAI211_X4 _54414_ (.A(_23216_),
    .B(_23218_),
    .C1(_10946_),
    .C2(_21823_),
    .ZN(_23219_));
 AOI221_X2 _54415_ (.A(_23219_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2158]),
    .B2(_10955_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2011]),
    .C2(_23156_),
    .ZN(_23220_));
 BUF_X32 _54416_ (.A(_10843_),
    .Z(_23221_));
 BUF_X8 _54417_ (.A(_22989_),
    .Z(_23222_));
 NAND3_X1 _54418_ (.A1(_23221_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2942]),
    .A3(_23222_),
    .ZN(_23223_));
 BUF_X8 _54419_ (.A(_10799_),
    .Z(_23224_));
 BUF_X8 _54420_ (.A(_10812_),
    .Z(_23225_));
 AOI22_X2 _54421_ (.A1(_23224_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3089]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3040]),
    .B2(_23225_),
    .ZN(_23226_));
 NAND3_X1 _54422_ (.A1(_22993_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2746]),
    .A3(_22999_),
    .ZN(_23227_));
 NAND3_X1 _54423_ (.A1(_22997_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2991]),
    .A3(_22999_),
    .ZN(_23228_));
 AND4_X4 _54424_ (.A1(_23223_),
    .A2(_23226_),
    .A3(_23227_),
    .A4(_23228_),
    .ZN(_23229_));
 BUF_X32 _54425_ (.A(_10873_),
    .Z(_23230_));
 BUF_X8 _54426_ (.A(_10935_),
    .Z(_23231_));
 AND3_X1 _54427_ (.A1(_23230_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1962]),
    .A3(_23231_),
    .ZN(_23232_));
 BUF_X16 _54428_ (.A(_10968_),
    .Z(_23233_));
 AOI221_X4 _54429_ (.A(_23232_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2060]),
    .B2(_23233_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2109]),
    .C2(_10962_),
    .ZN(_23234_));
 AND4_X1 _54430_ (.A1(_23214_),
    .A2(net40),
    .A3(_23229_),
    .A4(_23234_),
    .ZN(_23235_));
 BUF_X32 _54431_ (.A(_10803_),
    .Z(_23236_));
 BUF_X8 _54432_ (.A(_11125_),
    .Z(_23237_));
 NAND3_X1 _54433_ (.A1(_23236_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [737]),
    .A3(_23237_),
    .ZN(_23238_));
 AOI22_X4 _54434_ (.A1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [639]),
    .A2(_23107_),
    .B1(_11158_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [443]),
    .ZN(_23239_));
 BUF_X32 _54435_ (.A(_10817_),
    .Z(_23240_));
 NAND3_X1 _54436_ (.A1(_23240_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [688]),
    .A3(_11126_),
    .ZN(_23241_));
 BUF_X32 _54437_ (.A(_22900_),
    .Z(_23242_));
 NAND3_X1 _54438_ (.A1(_23242_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [590]),
    .A3(_11126_),
    .ZN(_23243_));
 AND4_X4 _54439_ (.A1(_23238_),
    .A2(_23239_),
    .A3(_23241_),
    .A4(_23243_),
    .ZN(_23244_));
 BUF_X32 _54440_ (.A(_10803_),
    .Z(_23245_));
 BUF_X8 _54441_ (.A(_22938_),
    .Z(_23246_));
 NAND3_X1 _54442_ (.A1(_23245_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [345]),
    .A3(_23246_),
    .ZN(_23247_));
 BUF_X16 _54443_ (.A(_11190_),
    .Z(_23248_));
 AOI22_X1 _54444_ (.A1(_23248_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [198]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [51]),
    .B2(_11211_),
    .ZN(_23249_));
 BUF_X8 _54445_ (.A(_22938_),
    .Z(_23250_));
 NAND3_X1 _54446_ (.A1(_10818_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [296]),
    .A3(_23250_),
    .ZN(_23251_));
 BUF_X32 _54447_ (.A(_22240_),
    .Z(_23252_));
 NAND3_X1 _54448_ (.A1(_23252_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [247]),
    .A3(_23250_),
    .ZN(_23253_));
 AND4_X1 _54449_ (.A1(_23247_),
    .A2(_23249_),
    .A3(_23251_),
    .A4(_23253_),
    .ZN(_23254_));
 BUF_X16 _54450_ (.A(_11123_),
    .Z(_23255_));
 AND3_X1 _54451_ (.A1(_23166_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [541]),
    .A3(_23255_),
    .ZN(_23256_));
 AOI221_X4 _54452_ (.A(_23256_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [492]),
    .B2(_11152_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [394]),
    .C2(_22733_),
    .ZN(_23257_));
 BUF_X16 _54453_ (.A(_11173_),
    .Z(_23258_));
 AND3_X1 _54454_ (.A1(_22521_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [100]),
    .A3(_23258_),
    .ZN(_23259_));
 AOI221_X4 _54455_ (.A(_23259_),
    .B1(_11205_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2]),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [149]),
    .C2(_22806_),
    .ZN(_23260_));
 AND4_X4 _54456_ (.A1(_23244_),
    .A2(_23254_),
    .A3(_23257_),
    .A4(_23260_),
    .ZN(_23261_));
 BUF_X16 _54457_ (.A(_11059_),
    .Z(_23262_));
 AOI22_X2 _54458_ (.A1(_22282_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1325]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1276]),
    .B2(_23262_),
    .ZN(_23263_));
 OAI221_X2 _54459_ (.A(_23263_),
    .B1(_22334_),
    .B2(_11066_),
    .C1(_22363_),
    .C2(_11070_),
    .ZN(_23264_));
 BUF_X16 _54460_ (.A(_11106_),
    .Z(_23265_));
 AOI22_X4 _54461_ (.A1(_23047_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [933]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [884]),
    .B2(_23265_),
    .ZN(_23266_));
 BUF_X16 _54462_ (.A(_11114_),
    .Z(_23267_));
 BUF_X16 _54463_ (.A(_11110_),
    .Z(_23268_));
 AOI22_X4 _54464_ (.A1(_23267_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [786]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [835]),
    .B2(_23268_),
    .ZN(_23269_));
 OAI211_X4 _54465_ (.A(_23266_),
    .B(_23269_),
    .C1(_22442_),
    .C2(_11091_),
    .ZN(_23270_));
 BUF_X16 _54466_ (.A(_10843_),
    .Z(_23271_));
 NAND3_X1 _54467_ (.A1(_23271_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [982]),
    .A3(_22976_),
    .ZN(_23272_));
 OAI221_X2 _54468_ (.A(_23272_),
    .B1(_11086_),
    .B2(_22416_),
    .C1(_11076_),
    .C2(_22390_),
    .ZN(_23273_));
 BUF_X8 _54469_ (.A(_11036_),
    .Z(_23274_));
 NAND3_X4 _54470_ (.A1(_23076_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1521]),
    .A3(_23274_),
    .ZN(_23275_));
 BUF_X16 _54471_ (.A(_10843_),
    .Z(_23276_));
 BUF_X8 _54472_ (.A(_11036_),
    .Z(_23277_));
 NAND3_X2 _54473_ (.A1(_23276_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1374]),
    .A3(_23277_),
    .ZN(_23278_));
 NAND3_X1 _54474_ (.A1(_23080_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1423]),
    .A3(_23205_),
    .ZN(_23279_));
 BUF_X32 _54475_ (.A(_10817_),
    .Z(_23280_));
 NAND3_X2 _54476_ (.A1(_23280_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1472]),
    .A3(_23205_),
    .ZN(_23281_));
 NAND4_X4 _54477_ (.A1(_23275_),
    .A2(_23278_),
    .A3(_23279_),
    .A4(_23281_),
    .ZN(_23282_));
 NOR4_X4 _54478_ (.A1(_23264_),
    .A2(_23270_),
    .A3(_23273_),
    .A4(_23282_),
    .ZN(_23283_));
 BUF_X32 _54479_ (.A(_22896_),
    .Z(_23284_));
 AND3_X1 _54480_ (.A1(_23284_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1913]),
    .A3(_22923_),
    .ZN(_23285_));
 BUF_X8 _54481_ (.A(_10997_),
    .Z(_23286_));
 AOI221_X2 _54482_ (.A(_23285_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1864]),
    .B2(_22003_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1815]),
    .C2(_23286_),
    .ZN(_23287_));
 BUF_X32 _54483_ (.A(_10855_),
    .Z(_23288_));
 AND3_X1 _54484_ (.A1(_23288_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1668]),
    .A3(_10988_),
    .ZN(_23289_));
 BUF_X16 _54485_ (.A(_22078_),
    .Z(_23290_));
 AOI21_X1 _54486_ (.A(_23289_),
    .B1(_23290_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1717]),
    .ZN(_23291_));
 NAND3_X1 _54487_ (.A1(_10879_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1570]),
    .A3(_10989_),
    .ZN(_23292_));
 BUF_X32 _54488_ (.A(_10867_),
    .Z(_23293_));
 BUF_X4 _54489_ (.A(_10988_),
    .Z(_23294_));
 NAND3_X1 _54490_ (.A1(_23293_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1619]),
    .A3(_23294_),
    .ZN(_23295_));
 BUF_X32 _54491_ (.A(_22900_),
    .Z(_23296_));
 NAND3_X1 _54492_ (.A1(_23296_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1766]),
    .A3(_23294_),
    .ZN(_23297_));
 AND4_X4 _54493_ (.A1(_23291_),
    .A2(_23292_),
    .A3(_23295_),
    .A4(_23297_),
    .ZN(_23298_));
 NAND3_X1 _54494_ (.A1(_22987_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2501]),
    .A3(_10892_),
    .ZN(_23299_));
 BUF_X16 _54495_ (.A(_10928_),
    .Z(_23300_));
 BUF_X8 _54496_ (.A(_10921_),
    .Z(_23301_));
 AOI22_X1 _54497_ (.A1(_23300_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2354]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2403]),
    .B2(_23301_),
    .ZN(_23302_));
 BUF_X32 _54498_ (.A(_22240_),
    .Z(_23303_));
 BUF_X4 _54499_ (.A(_10891_),
    .Z(_23304_));
 NAND3_X1 _54500_ (.A1(_23303_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2599]),
    .A3(_23304_),
    .ZN(_23305_));
 BUF_X32 _54501_ (.A(_22522_),
    .Z(_23306_));
 NAND3_X1 _54502_ (.A1(_23306_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2452]),
    .A3(_23304_),
    .ZN(_23307_));
 AND4_X2 _54503_ (.A1(_23299_),
    .A2(_23302_),
    .A3(_23305_),
    .A4(_23307_),
    .ZN(_23308_));
 BUF_X32 _54504_ (.A(net73),
    .Z(_23309_));
 BUF_X8 _54505_ (.A(_10886_),
    .Z(_23310_));
 AND3_X1 _54506_ (.A1(_23309_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2550]),
    .A3(_23310_),
    .ZN(_23311_));
 AOI221_X4 _54507_ (.A(_23311_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2648]),
    .B2(_21601_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2697]),
    .C2(_21573_),
    .ZN(_23312_));
 AND4_X2 _54508_ (.A1(net55),
    .A2(_23298_),
    .A3(_23308_),
    .A4(_23312_),
    .ZN(_23313_));
 NAND4_X1 _54509_ (.A1(_23235_),
    .A2(_23261_),
    .A3(net11),
    .A4(_23313_),
    .ZN(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [2]));
 AND3_X1 _54510_ (.A1(_22900_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1375]),
    .A3(_22898_),
    .ZN(_23314_));
 BUF_X16 _54511_ (.A(_11031_),
    .Z(_23315_));
 AOI221_X4 _54512_ (.A(_23314_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1473]),
    .B2(_22210_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1522]),
    .C2(_23315_),
    .ZN(_23316_));
 BUF_X16 _54513_ (.A(_11080_),
    .Z(_23317_));
 NAND3_X1 _54514_ (.A1(_23204_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [885]),
    .A3(_23317_),
    .ZN(_23318_));
 AND3_X1 _54515_ (.A1(_10757_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1326]),
    .A3(_11034_),
    .ZN(_23319_));
 AOI221_X2 _54516_ (.A(_23319_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1277]),
    .B2(_11059_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1228]),
    .C2(_11065_),
    .ZN(_23320_));
 BUF_X8 _54517_ (.A(_11080_),
    .Z(_23321_));
 NAND3_X1 _54518_ (.A1(_22993_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [787]),
    .A3(_23321_),
    .ZN(_23322_));
 NAND3_X1 _54519_ (.A1(_22987_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [934]),
    .A3(_23321_),
    .ZN(_23323_));
 AND4_X1 _54520_ (.A1(_23318_),
    .A2(_23320_),
    .A3(_23322_),
    .A4(_23323_),
    .ZN(_23324_));
 BUF_X16 _54521_ (.A(_11069_),
    .Z(_23325_));
 BUF_X16 _54522_ (.A(_22232_),
    .Z(_23326_));
 AOI22_X2 _54523_ (.A1(_23325_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1179]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1424]),
    .B2(_23326_),
    .ZN(_23327_));
 BUF_X32 _54524_ (.A(_10843_),
    .Z(_23328_));
 BUF_X4 _54525_ (.A(_11080_),
    .Z(_23329_));
 NAND3_X1 _54526_ (.A1(_23328_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [983]),
    .A3(_23329_),
    .ZN(_23330_));
 BUF_X16 _54527_ (.A(_11075_),
    .Z(_23331_));
 BUF_X8 _54528_ (.A(_11085_),
    .Z(_23332_));
 BUF_X16 _54529_ (.A(_23332_),
    .Z(_23333_));
 AOI22_X1 _54530_ (.A1(_23331_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1130]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1081]),
    .B2(_23333_),
    .ZN(_23334_));
 NAND3_X1 _54531_ (.A1(_22997_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1032]),
    .A3(_23321_),
    .ZN(_23335_));
 NAND3_X1 _54532_ (.A1(_23293_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [836]),
    .A3(_11081_),
    .ZN(_23336_));
 AND4_X1 _54533_ (.A1(_23330_),
    .A2(_23334_),
    .A3(_23335_),
    .A4(_23336_),
    .ZN(_23337_));
 AND4_X4 _54534_ (.A1(_23316_),
    .A2(_23324_),
    .A3(_23327_),
    .A4(_23337_),
    .ZN(_23338_));
 BUF_X32 _54535_ (.A(_22900_),
    .Z(_23339_));
 BUF_X32 _54536_ (.A(_23339_),
    .Z(_23340_));
 BUF_X16 _54537_ (.A(_23250_),
    .Z(_23341_));
 NAND3_X1 _54538_ (.A1(_23340_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [199]),
    .A3(_23341_),
    .ZN(_23342_));
 NAND3_X1 _54539_ (.A1(_23328_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [591]),
    .A3(_11126_),
    .ZN(_23343_));
 AND3_X1 _54540_ (.A1(_10757_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [542]),
    .A3(_11123_),
    .ZN(_23344_));
 AOI221_X2 _54541_ (.A(_23344_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [493]),
    .B2(_11151_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [395]),
    .C2(_11164_),
    .ZN(_23345_));
 BUF_X8 _54542_ (.A(_11125_),
    .Z(_23346_));
 NAND3_X1 _54543_ (.A1(_23293_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [444]),
    .A3(_23346_),
    .ZN(_23347_));
 AND3_X1 _54544_ (.A1(_10811_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [689]),
    .A3(_11123_),
    .ZN(_23348_));
 AOI221_X2 _54545_ (.A(_23348_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [640]),
    .B2(_11136_),
    .C1(_22597_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [738]),
    .ZN(_23349_));
 AND4_X4 _54546_ (.A1(_23343_),
    .A2(_23345_),
    .A3(_23347_),
    .A4(_23349_),
    .ZN(_23350_));
 AND3_X1 _54547_ (.A1(_23168_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [248]),
    .A3(_23258_),
    .ZN(_23351_));
 AOI221_X4 _54548_ (.A(_23351_),
    .B1(_22903_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [297]),
    .C1(_11170_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [346]),
    .ZN(_23352_));
 AND3_X1 _54549_ (.A1(_10877_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3]),
    .A3(_11173_),
    .ZN(_23353_));
 AND3_X1 _54550_ (.A1(_10920_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [52]),
    .A3(_11173_),
    .ZN(_23354_));
 OR2_X1 _54551_ (.A1(_23353_),
    .A2(_23354_),
    .ZN(_23355_));
 AOI221_X2 _54552_ (.A(_23355_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [101]),
    .B2(_11200_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [150]),
    .C2(_22806_),
    .ZN(_23356_));
 AND4_X4 _54553_ (.A1(_23342_),
    .A2(_23350_),
    .A3(_23352_),
    .A4(_23356_),
    .ZN(_23357_));
 AND3_X1 _54554_ (.A1(_23173_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2453]),
    .A3(_23012_),
    .ZN(_23358_));
 AOI221_X2 _54555_ (.A(_23358_),
    .B1(_23300_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2355]),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2502]),
    .C2(_10912_),
    .ZN(_23359_));
 BUF_X8 _54556_ (.A(_22989_),
    .Z(_23360_));
 BUF_X8 _54557_ (.A(_23360_),
    .Z(_23361_));
 NAND3_X2 _54558_ (.A1(_10869_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2796]),
    .A3(_23361_),
    .ZN(_23362_));
 NAND3_X1 _54559_ (.A1(_22524_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2845]),
    .A3(_23361_),
    .ZN(_23363_));
 NAND3_X2 _54560_ (.A1(_22985_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2894]),
    .A3(_23361_),
    .ZN(_23364_));
 NAND4_X4 _54561_ (.A1(_23359_),
    .A2(_23362_),
    .A3(_23363_),
    .A4(_23364_),
    .ZN(_23365_));
 AOI22_X4 _54562_ (.A1(_10800_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3090]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3041]),
    .B2(_10813_),
    .ZN(_23366_));
 BUF_X32 _54563_ (.A(_22900_),
    .Z(_23367_));
 BUF_X32 _54564_ (.A(_23367_),
    .Z(_23368_));
 NAND3_X1 _54565_ (.A1(_23368_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2943]),
    .A3(_22991_),
    .ZN(_23369_));
 NAND3_X1 _54566_ (.A1(_22998_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2992]),
    .A3(_23000_),
    .ZN(_23370_));
 NAND3_X1 _54567_ (.A1(_22994_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2747]),
    .A3(_23123_),
    .ZN(_23371_));
 NAND4_X1 _54568_ (.A1(_23366_),
    .A2(_23369_),
    .A3(_23370_),
    .A4(_23371_),
    .ZN(_23372_));
 BUF_X16 _54569_ (.A(_10887_),
    .Z(_23373_));
 BUF_X16 _54570_ (.A(_21600_),
    .Z(_23374_));
 AOI22_X4 _54571_ (.A1(_23373_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2698]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2649]),
    .B2(_23374_),
    .ZN(_23375_));
 NAND3_X2 _54572_ (.A1(_22998_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2600]),
    .A3(_23120_),
    .ZN(_23376_));
 BUF_X32 _54573_ (.A(_23035_),
    .Z(_23377_));
 NAND3_X2 _54574_ (.A1(_23377_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2404]),
    .A3(_23120_),
    .ZN(_23378_));
 NAND3_X2 _54575_ (.A1(_22933_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2551]),
    .A3(_23120_),
    .ZN(_23379_));
 NAND4_X4 _54576_ (.A1(_23375_),
    .A2(_23376_),
    .A3(_23378_),
    .A4(_23379_),
    .ZN(_23380_));
 NOR3_X1 _54577_ (.A1(_23365_),
    .A2(_23372_),
    .A3(_23380_),
    .ZN(_23381_));
 BUF_X32 _54578_ (.A(_10877_),
    .Z(_23382_));
 AND3_X1 _54579_ (.A1(_23382_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1963]),
    .A3(_23231_),
    .ZN(_23383_));
 AOI221_X4 _54580_ (.A(_23383_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2061]),
    .B2(_22910_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2110]),
    .C2(_10962_),
    .ZN(_23384_));
 BUF_X32 _54581_ (.A(_22240_),
    .Z(_23385_));
 NAND3_X1 _54582_ (.A1(_23385_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2208]),
    .A3(_10941_),
    .ZN(_23386_));
 AOI22_X1 _54583_ (.A1(_10956_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2159]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2012]),
    .B2(_21937_),
    .ZN(_23387_));
 BUF_X8 _54584_ (.A(_10940_),
    .Z(_23388_));
 NAND3_X1 _54585_ (.A1(_10818_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2257]),
    .A3(_23388_),
    .ZN(_23389_));
 BUF_X32 _54586_ (.A(_10803_),
    .Z(_23390_));
 NAND3_X1 _54587_ (.A1(_23390_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2306]),
    .A3(_23388_),
    .ZN(_23391_));
 AND4_X2 _54588_ (.A1(_23386_),
    .A2(_23387_),
    .A3(_23389_),
    .A4(_23391_),
    .ZN(_23392_));
 BUF_X8 _54589_ (.A(_10988_),
    .Z(_23393_));
 NAND3_X1 _54590_ (.A1(_22987_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1718]),
    .A3(_23393_),
    .ZN(_23394_));
 BUF_X16 _54591_ (.A(_11025_),
    .Z(_23395_));
 BUF_X8 _54592_ (.A(_11019_),
    .Z(_23396_));
 AOI22_X2 _54593_ (.A1(_23395_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1571]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1620]),
    .B2(_23396_),
    .ZN(_23397_));
 BUF_X8 _54594_ (.A(_10988_),
    .Z(_23398_));
 NAND3_X1 _54595_ (.A1(_22932_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1767]),
    .A3(_23398_),
    .ZN(_23399_));
 NAND3_X1 _54596_ (.A1(_23306_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1669]),
    .A3(_23398_),
    .ZN(_23400_));
 AND4_X4 _54597_ (.A1(_23394_),
    .A2(_23397_),
    .A3(_23399_),
    .A4(_23400_),
    .ZN(_23401_));
 BUF_X8 _54598_ (.A(_10982_),
    .Z(_23402_));
 AND3_X1 _54599_ (.A1(_23217_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1914]),
    .A3(_23402_),
    .ZN(_23403_));
 AOI221_X2 _54600_ (.A(_23403_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1865]),
    .B2(_10993_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1816]),
    .C2(_23286_),
    .ZN(_23404_));
 AND4_X4 _54601_ (.A1(_23384_),
    .A2(_23392_),
    .A3(_23401_),
    .A4(_23404_),
    .ZN(_23405_));
 NAND4_X1 _54602_ (.A1(_23338_),
    .A2(_23357_),
    .A3(_23381_),
    .A4(_23405_),
    .ZN(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [3]));
 AND3_X1 _54603_ (.A1(_10867_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1229]),
    .A3(_22898_),
    .ZN(_23406_));
 AOI221_X4 _54604_ (.A(_23406_),
    .B1(_11060_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1278]),
    .C1(_22282_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1327]),
    .ZN(_23407_));
 BUF_X32 _54605_ (.A(_10811_),
    .Z(_23408_));
 NAND3_X1 _54606_ (.A1(_23408_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [690]),
    .A3(_23255_),
    .ZN(_23409_));
 OAI221_X2 _54607_ (.A(_23409_),
    .B1(_11142_),
    .B2(_22669_),
    .C1(_11121_),
    .C2(_22604_),
    .ZN(_23410_));
 AOI221_X2 _54608_ (.A(_23410_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [641]),
    .B2(_23107_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [445]),
    .C2(_11159_),
    .ZN(_23411_));
 BUF_X8 _54609_ (.A(_22980_),
    .Z(_23412_));
 NAND3_X1 _54610_ (.A1(_23328_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1376]),
    .A3(_23412_),
    .ZN(_23413_));
 AOI22_X2 _54611_ (.A1(_23315_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1523]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1474]),
    .B2(_22210_),
    .ZN(_23414_));
 NAND3_X1 _54612_ (.A1(_22997_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1425]),
    .A3(_23050_),
    .ZN(_23415_));
 NAND3_X1 _54613_ (.A1(_10879_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1180]),
    .A3(_23050_),
    .ZN(_23416_));
 AND4_X4 _54614_ (.A1(_23413_),
    .A2(_23414_),
    .A3(_23415_),
    .A4(_23416_),
    .ZN(_23417_));
 AND3_X1 _54615_ (.A1(_23158_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [543]),
    .A3(_23161_),
    .ZN(_23418_));
 AOI221_X4 _54616_ (.A(_23418_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [494]),
    .B2(_11152_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [396]),
    .C2(_22733_),
    .ZN(_23419_));
 AND4_X4 _54617_ (.A1(_23407_),
    .A2(_23411_),
    .A3(_23417_),
    .A4(_23419_),
    .ZN(_23420_));
 BUF_X32 _54618_ (.A(_10779_),
    .Z(_23421_));
 BUF_X16 _54619_ (.A(_10891_),
    .Z(_23422_));
 NAND3_X1 _54620_ (.A1(_23421_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2503]),
    .A3(_23422_),
    .ZN(_23423_));
 AND3_X1 _54621_ (.A1(_10866_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2797]),
    .A3(_10787_),
    .ZN(_23424_));
 AOI221_X2 _54622_ (.A(_23424_),
    .B1(_10851_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2846]),
    .C1(_10773_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2895]),
    .ZN(_23425_));
 BUF_X16 _54623_ (.A(_23041_),
    .Z(_23426_));
 BUF_X4 _54624_ (.A(_10891_),
    .Z(_23427_));
 NAND3_X1 _54625_ (.A1(_23426_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2405]),
    .A3(_23427_),
    .ZN(_23428_));
 NAND3_X1 _54626_ (.A1(_23204_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2454]),
    .A3(_23427_),
    .ZN(_23429_));
 AND4_X1 _54627_ (.A1(_23423_),
    .A2(_23425_),
    .A3(_23428_),
    .A4(_23429_),
    .ZN(_23430_));
 BUF_X16 _54628_ (.A(_22928_),
    .Z(_23431_));
 NAND3_X1 _54629_ (.A1(_23207_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2748]),
    .A3(_23431_),
    .ZN(_23432_));
 AOI22_X2 _54630_ (.A1(_23224_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3091]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3042]),
    .B2(_10813_),
    .ZN(_23433_));
 BUF_X32 _54631_ (.A(_22240_),
    .Z(_23434_));
 NAND3_X1 _54632_ (.A1(_23434_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2993]),
    .A3(_23222_),
    .ZN(_23435_));
 NAND3_X1 _54633_ (.A1(_23328_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2944]),
    .A3(_23222_),
    .ZN(_23436_));
 AND4_X4 _54634_ (.A1(_23432_),
    .A2(_23433_),
    .A3(_23435_),
    .A4(_23436_),
    .ZN(_23437_));
 BUF_X32 _54635_ (.A(_22240_),
    .Z(_23438_));
 NAND3_X1 _54636_ (.A1(_23438_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2601]),
    .A3(_23422_),
    .ZN(_23439_));
 AOI22_X1 _54637_ (.A1(_23373_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2699]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2650]),
    .B2(_23374_),
    .ZN(_23440_));
 NAND3_X1 _54638_ (.A1(_23328_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2552]),
    .A3(_23427_),
    .ZN(_23441_));
 NAND3_X1 _54639_ (.A1(_22993_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2356]),
    .A3(_23427_),
    .ZN(_23442_));
 AND4_X1 _54640_ (.A1(_23439_),
    .A2(_23440_),
    .A3(_23441_),
    .A4(_23442_),
    .ZN(_23443_));
 AND3_X2 _54641_ (.A1(_23430_),
    .A2(_23437_),
    .A3(_23443_),
    .ZN(_23444_));
 AND3_X1 _54642_ (.A1(_23284_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [347]),
    .A3(_11174_),
    .ZN(_23445_));
 BUF_X16 _54643_ (.A(_11186_),
    .Z(_23446_));
 AOI221_X2 _54644_ (.A(_23445_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [298]),
    .B2(_11181_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [249]),
    .C2(_23446_),
    .ZN(_23447_));
 OAI22_X1 _54645_ (.A1(_11115_),
    .A2(_22580_),
    .B1(_22552_),
    .B2(_11111_),
    .ZN(_23448_));
 OAI22_X2 _54646_ (.A1(_11101_),
    .A2(_22501_),
    .B1(_22527_),
    .B2(_11107_),
    .ZN(_23449_));
 AOI211_X2 _54647_ (.A(_23448_),
    .B(_23449_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [984]),
    .C2(_22459_),
    .ZN(_23450_));
 BUF_X16 _54648_ (.A(_22938_),
    .Z(_23451_));
 NAND3_X1 _54649_ (.A1(_23113_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [53]),
    .A3(_23451_),
    .ZN(_23452_));
 BUF_X16 _54650_ (.A(_11200_),
    .Z(_23453_));
 AOI22_X1 _54651_ (.A1(_22806_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [151]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [102]),
    .B2(_23453_),
    .ZN(_23454_));
 BUF_X32 _54652_ (.A(_10878_),
    .Z(_23455_));
 NAND3_X1 _54653_ (.A1(_23455_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [4]),
    .A3(_22939_),
    .ZN(_23456_));
 NAND3_X1 _54654_ (.A1(_22932_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [200]),
    .A3(_22939_),
    .ZN(_23457_));
 AND4_X2 _54655_ (.A1(_23452_),
    .A2(_23454_),
    .A3(_23456_),
    .A4(_23457_),
    .ZN(_23458_));
 BUF_X32 _54656_ (.A(_10797_),
    .Z(_23459_));
 BUF_X8 _54657_ (.A(_11089_),
    .Z(_23460_));
 AND3_X1 _54658_ (.A1(_23459_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1131]),
    .A3(_23460_),
    .ZN(_23461_));
 AOI221_X2 _54659_ (.A(_23461_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1082]),
    .B2(_23332_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1033]),
    .C2(_22435_),
    .ZN(_23462_));
 AND4_X4 _54660_ (.A1(_23447_),
    .A2(net16),
    .A3(_23458_),
    .A4(net54),
    .ZN(_23463_));
 AND3_X1 _54661_ (.A1(_23382_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1964]),
    .A3(_23231_),
    .ZN(_23464_));
 AOI221_X4 _54662_ (.A(_23464_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2062]),
    .B2(_23233_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2111]),
    .C2(_10962_),
    .ZN(_23465_));
 NAND3_X1 _54663_ (.A1(_23242_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1768]),
    .A3(_23393_),
    .ZN(_23466_));
 BUF_X16 _54664_ (.A(_22078_),
    .Z(_23467_));
 AOI22_X2 _54665_ (.A1(_23467_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1719]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1670]),
    .B2(_22105_),
    .ZN(_23468_));
 NAND3_X1 _54666_ (.A1(_23293_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1621]),
    .A3(_23294_),
    .ZN(_23469_));
 NAND3_X1 _54667_ (.A1(_23455_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1572]),
    .A3(_23294_),
    .ZN(_23470_));
 AND4_X4 _54668_ (.A1(_23466_),
    .A2(_23468_),
    .A3(_23469_),
    .A4(_23470_),
    .ZN(_23471_));
 NAND3_X1 _54669_ (.A1(_22949_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2307]),
    .A3(_23005_),
    .ZN(_23472_));
 OAI21_X2 _54670_ (.A(_23472_),
    .B1(_10946_),
    .B2(_21825_),
    .ZN(_23473_));
 AND3_X1 _54671_ (.A1(_10843_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2160]),
    .A3(_22963_),
    .ZN(_23474_));
 AND3_X1 _54672_ (.A1(_22240_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2209]),
    .A3(_10940_),
    .ZN(_23475_));
 AND3_X1 _54673_ (.A1(_23041_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2013]),
    .A3(_10940_),
    .ZN(_23476_));
 NOR4_X2 _54674_ (.A1(_23473_),
    .A2(_23474_),
    .A3(_23475_),
    .A4(_23476_),
    .ZN(_23477_));
 AND3_X1 _54675_ (.A1(_23217_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1915]),
    .A3(_23402_),
    .ZN(_23478_));
 AOI221_X2 _54676_ (.A(_23478_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1866]),
    .B2(_10993_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1817]),
    .C2(_23286_),
    .ZN(_23479_));
 AND4_X4 _54677_ (.A1(_23465_),
    .A2(_23471_),
    .A3(_23477_),
    .A4(_23479_),
    .ZN(_23480_));
 NAND4_X1 _54678_ (.A1(_23420_),
    .A2(_23444_),
    .A3(_23463_),
    .A4(_23480_),
    .ZN(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [4]));
 BUF_X8 _54679_ (.A(_10890_),
    .Z(_23481_));
 NAND3_X2 _54680_ (.A1(_22897_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2700]),
    .A3(_23481_),
    .ZN(_23482_));
 NAND3_X1 _54681_ (.A1(_22900_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2553]),
    .A3(_23481_),
    .ZN(_23483_));
 NAND2_X4 _54682_ (.A1(_23482_),
    .A2(_23483_),
    .ZN(_23484_));
 BUF_X16 _54683_ (.A(_10976_),
    .Z(_23485_));
 AOI221_X2 _54684_ (.A(_23484_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2259]),
    .B2(_21816_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1965]),
    .C2(_23485_),
    .ZN(_23486_));
 BUF_X32 _54685_ (.A(_22896_),
    .Z(_23487_));
 NAND3_X2 _54686_ (.A1(_23487_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [740]),
    .A3(_23161_),
    .ZN(_23488_));
 OAI21_X4 _54687_ (.A(_23488_),
    .B1(_11132_),
    .B2(_22628_),
    .ZN(_23489_));
 BUF_X16 _54688_ (.A(_11211_),
    .Z(_23490_));
 AOI221_X2 _54689_ (.A(_23489_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [103]),
    .B2(_23453_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [54]),
    .C2(_23490_),
    .ZN(_23491_));
 BUF_X32 _54690_ (.A(_22896_),
    .Z(_23492_));
 NAND3_X1 _54691_ (.A1(_23492_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1916]),
    .A3(_22921_),
    .ZN(_23493_));
 BUF_X16 _54692_ (.A(_11079_),
    .Z(_23494_));
 NAND3_X4 _54693_ (.A1(_22942_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1083]),
    .A3(_23494_),
    .ZN(_23495_));
 NAND2_X1 _54694_ (.A1(_23493_),
    .A2(_23495_),
    .ZN(_23496_));
 AOI221_X2 _54695_ (.A(_23496_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1867]),
    .B2(_22003_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1720]),
    .C2(_23467_),
    .ZN(_23497_));
 BUF_X16 _54696_ (.A(_10787_),
    .Z(_23498_));
 NAND3_X1 _54697_ (.A1(_22920_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3043]),
    .A3(_23498_),
    .ZN(_23499_));
 NAND3_X1 _54698_ (.A1(_10829_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2994]),
    .A3(_23498_),
    .ZN(_23500_));
 NAND2_X1 _54699_ (.A1(_23499_),
    .A2(_23500_),
    .ZN(_23501_));
 AOI221_X4 _54700_ (.A(_23501_),
    .B1(_21289_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2749]),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3092]),
    .C2(_10799_),
    .ZN(_23502_));
 AND4_X1 _54701_ (.A1(net39),
    .A2(_23491_),
    .A3(net38),
    .A4(_23502_),
    .ZN(_23503_));
 BUF_X16 _54702_ (.A(_11124_),
    .Z(_23504_));
 NAND3_X1 _54703_ (.A1(_22915_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [446]),
    .A3(_23504_),
    .ZN(_23505_));
 NAND3_X1 _54704_ (.A1(_10829_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [642]),
    .A3(_23151_),
    .ZN(_23506_));
 NAND2_X1 _54705_ (.A1(_23505_),
    .A2(_23506_),
    .ZN(_23507_));
 AOI221_X4 _54706_ (.A(_23507_),
    .B1(_23104_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [985]),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1132]),
    .C2(_23331_),
    .ZN(_23508_));
 BUF_X32 _54707_ (.A(_10778_),
    .Z(_23509_));
 BUF_X16 _54708_ (.A(_11124_),
    .Z(_23510_));
 NAND3_X1 _54709_ (.A1(_23509_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [544]),
    .A3(_23510_),
    .ZN(_23511_));
 BUF_X8 _54710_ (.A(_11145_),
    .Z(_23512_));
 NAND3_X1 _54711_ (.A1(_23382_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [397]),
    .A3(_23512_),
    .ZN(_23513_));
 NAND2_X1 _54712_ (.A1(_23511_),
    .A2(_23513_),
    .ZN(_23514_));
 BUF_X16 _54713_ (.A(_11141_),
    .Z(_23515_));
 AOI221_X4 _54714_ (.A(_23514_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [593]),
    .B2(_23515_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [495]),
    .C2(_11153_),
    .ZN(_23516_));
 NAND3_X2 _54715_ (.A1(_23230_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1573]),
    .A3(_22923_),
    .ZN(_23517_));
 BUF_X32 _54716_ (.A(_10842_),
    .Z(_23518_));
 BUF_X8 _54717_ (.A(_10982_),
    .Z(_23519_));
 NAND3_X2 _54718_ (.A1(_23518_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1769]),
    .A3(_23519_),
    .ZN(_23520_));
 NAND2_X4 _54719_ (.A1(_23517_),
    .A2(_23520_),
    .ZN(_23521_));
 AOI221_X2 _54720_ (.A(_23521_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2945]),
    .B2(_10838_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2651]),
    .C2(_23374_),
    .ZN(_23522_));
 NAND3_X2 _54721_ (.A1(_23518_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [201]),
    .A3(_23159_),
    .ZN(_23523_));
 BUF_X32 _54722_ (.A(_10811_),
    .Z(_23524_));
 NAND3_X2 _54723_ (.A1(_23524_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [299]),
    .A3(_23258_),
    .ZN(_23525_));
 NAND2_X4 _54724_ (.A1(_23523_),
    .A2(_23525_),
    .ZN(_23526_));
 AOI221_X4 _54725_ (.A(_23526_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2063]),
    .B2(_23233_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2014]),
    .C2(_23156_),
    .ZN(_23527_));
 AND4_X1 _54726_ (.A1(_23508_),
    .A2(_23516_),
    .A3(_23522_),
    .A4(_23527_),
    .ZN(_23528_));
 NAND3_X2 _54727_ (.A1(_22985_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [936]),
    .A3(_11082_),
    .ZN(_23529_));
 NAND3_X2 _54728_ (.A1(_22242_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1034]),
    .A3(_11082_),
    .ZN(_23530_));
 NAND3_X4 _54729_ (.A1(_22524_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1279]),
    .A3(_23051_),
    .ZN(_23531_));
 NAND3_X4 _54730_ (.A1(_23114_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1230]),
    .A3(_22945_),
    .ZN(_23532_));
 NAND4_X4 _54731_ (.A1(_23529_),
    .A2(_23530_),
    .A3(_23531_),
    .A4(_23532_),
    .ZN(_23533_));
 NAND3_X1 _54732_ (.A1(_23004_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [152]),
    .A3(_22940_),
    .ZN(_23534_));
 NAND3_X1 _54733_ (.A1(_22950_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [348]),
    .A3(_22951_),
    .ZN(_23535_));
 BUF_X32 _54734_ (.A(_10830_),
    .Z(_23536_));
 NAND3_X2 _54735_ (.A1(_23536_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [250]),
    .A3(_11176_),
    .ZN(_23537_));
 NAND3_X4 _54736_ (.A1(_23189_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2406]),
    .A3(_23068_),
    .ZN(_23538_));
 NAND4_X2 _54737_ (.A1(_23534_),
    .A2(_23535_),
    .A3(_23537_),
    .A4(_23538_),
    .ZN(_23539_));
 NAND3_X2 _54738_ (.A1(_23020_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2896]),
    .A3(_23128_),
    .ZN(_23540_));
 NAND3_X1 _54739_ (.A1(_22958_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2602]),
    .A3(_23023_),
    .ZN(_23541_));
 NAND3_X2 _54740_ (.A1(_23194_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2357]),
    .A3(_23026_),
    .ZN(_23542_));
 NAND3_X2 _54741_ (.A1(_23078_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2455]),
    .A3(_23029_),
    .ZN(_23543_));
 NAND4_X4 _54742_ (.A1(_23540_),
    .A2(_23541_),
    .A3(_23542_),
    .A4(_23543_),
    .ZN(_23544_));
 NAND3_X2 _54743_ (.A1(_23032_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [789]),
    .A3(_22970_),
    .ZN(_23545_));
 NAND3_X4 _54744_ (.A1(_23036_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [838]),
    .A3(_22976_),
    .ZN(_23546_));
 BUF_X16 _54745_ (.A(_11080_),
    .Z(_23547_));
 NAND3_X1 _54746_ (.A1(_23039_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [887]),
    .A3(_23547_),
    .ZN(_23548_));
 NAND3_X4 _54747_ (.A1(_23042_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2798]),
    .A3(_23431_),
    .ZN(_23549_));
 NAND4_X4 _54748_ (.A1(_23545_),
    .A2(_23546_),
    .A3(_23548_),
    .A4(_23549_),
    .ZN(_23550_));
 NOR4_X1 _54749_ (.A1(_23533_),
    .A2(_23539_),
    .A3(_23544_),
    .A4(_23550_),
    .ZN(_23551_));
 NAND3_X4 _54750_ (.A1(_10805_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1524]),
    .A3(_23051_),
    .ZN(_23552_));
 BUF_X16 _54751_ (.A(_10940_),
    .Z(_23553_));
 BUF_X8 _54752_ (.A(_23553_),
    .Z(_23554_));
 NAND3_X2 _54753_ (.A1(_22988_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2112]),
    .A3(_23554_),
    .ZN(_23555_));
 NAND3_X2 _54754_ (.A1(_23368_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2161]),
    .A3(_23554_),
    .ZN(_23556_));
 NAND3_X2 _54755_ (.A1(_10831_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2210]),
    .A3(_23006_),
    .ZN(_23557_));
 NAND4_X4 _54756_ (.A1(_23552_),
    .A2(_23555_),
    .A3(_23556_),
    .A4(_23557_),
    .ZN(_23558_));
 NAND3_X2 _54757_ (.A1(_23125_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2504]),
    .A3(_23131_),
    .ZN(_23559_));
 BUF_X32 _54758_ (.A(_22949_),
    .Z(_23560_));
 BUF_X8 _54759_ (.A(_22963_),
    .Z(_23561_));
 NAND3_X4 _54760_ (.A1(_23560_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2308]),
    .A3(_23561_),
    .ZN(_23562_));
 NAND3_X2 _54761_ (.A1(_22968_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [5]),
    .A3(_23187_),
    .ZN(_23563_));
 NAND3_X4 _54762_ (.A1(_23016_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2847]),
    .A3(_23033_),
    .ZN(_23564_));
 NAND4_X4 _54763_ (.A1(_23559_),
    .A2(_23562_),
    .A3(_23563_),
    .A4(_23564_),
    .ZN(_23565_));
 BUF_X8 _54764_ (.A(_11036_),
    .Z(_23566_));
 NAND3_X2 _54765_ (.A1(_23020_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1328]),
    .A3(_23566_),
    .ZN(_23567_));
 NAND3_X2 _54766_ (.A1(_22972_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1475]),
    .A3(_23274_),
    .ZN(_23568_));
 NAND3_X2 _54767_ (.A1(_23271_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1377]),
    .A3(_22981_),
    .ZN(_23569_));
 NAND3_X2 _54768_ (.A1(_22978_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1426]),
    .A3(_22981_),
    .ZN(_23570_));
 NAND4_X4 _54769_ (.A1(_23567_),
    .A2(_23568_),
    .A3(_23569_),
    .A4(_23570_),
    .ZN(_23571_));
 NAND3_X2 _54770_ (.A1(_23032_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1181]),
    .A3(_23274_),
    .ZN(_23572_));
 NAND3_X2 _54771_ (.A1(_23078_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1671]),
    .A3(_23146_),
    .ZN(_23573_));
 NAND3_X2 _54772_ (.A1(_23042_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1622]),
    .A3(_23146_),
    .ZN(_23574_));
 BUF_X16 _54773_ (.A(_10830_),
    .Z(_23575_));
 BUF_X16 _54774_ (.A(_22934_),
    .Z(_23576_));
 NAND3_X2 _54775_ (.A1(_23575_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1818]),
    .A3(_23576_),
    .ZN(_23577_));
 NAND4_X4 _54776_ (.A1(_23572_),
    .A2(_23573_),
    .A3(_23574_),
    .A4(_23577_),
    .ZN(_23578_));
 NOR4_X4 _54777_ (.A1(_23558_),
    .A2(_23565_),
    .A3(_23571_),
    .A4(_23578_),
    .ZN(_23579_));
 NAND4_X1 _54778_ (.A1(_23503_),
    .A2(_23528_),
    .A3(_23551_),
    .A4(_23579_),
    .ZN(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [5]));
 AND3_X4 _54779_ (.A1(_10778_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2897]),
    .A3(_10787_),
    .ZN(_23580_));
 AND3_X1 _54780_ (.A1(_10855_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2064]),
    .A3(_10939_),
    .ZN(_23581_));
 OR2_X1 _54781_ (.A1(_23580_),
    .A2(_23581_),
    .ZN(_23582_));
 AOI221_X2 _54782_ (.A(_23582_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2260]),
    .B2(_21816_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1770]),
    .C2(_11003_),
    .ZN(_23583_));
 BUF_X8 _54783_ (.A(_21978_),
    .Z(_23584_));
 AOI22_X1 _54784_ (.A1(_23584_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1917]),
    .B1(_23286_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1819]),
    .ZN(_23585_));
 AND3_X2 _54785_ (.A1(_10867_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2799]),
    .A3(_22989_),
    .ZN(_23586_));
 BUF_X16 _54786_ (.A(_10912_),
    .Z(_23587_));
 AOI21_X4 _54787_ (.A(_23586_),
    .B1(_23587_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2505]),
    .ZN(_23588_));
 AND3_X2 _54788_ (.A1(_23288_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2848]),
    .A3(_22989_),
    .ZN(_23589_));
 AOI21_X4 _54789_ (.A(_23589_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2456]),
    .B2(_21705_),
    .ZN(_23590_));
 BUF_X16 _54790_ (.A(_11012_),
    .Z(_23591_));
 AOI22_X4 _54791_ (.A1(_23591_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1672]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2015]),
    .B2(_23156_),
    .ZN(_23592_));
 AND4_X1 _54792_ (.A1(_23585_),
    .A2(_23588_),
    .A3(_23590_),
    .A4(_23592_),
    .ZN(_23593_));
 AOI22_X2 _54793_ (.A1(_10956_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2162]),
    .B1(_22003_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1868]),
    .ZN(_23594_));
 BUF_X16 _54794_ (.A(_11025_),
    .Z(_23595_));
 AOI22_X2 _54795_ (.A1(_23595_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1574]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2211]),
    .B2(_10950_),
    .ZN(_23596_));
 AND4_X4 _54796_ (.A1(_23583_),
    .A2(_23593_),
    .A3(_23594_),
    .A4(_23596_),
    .ZN(_23597_));
 AOI22_X4 _54797_ (.A1(_23265_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [888]),
    .B1(_23268_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [839]),
    .ZN(_23598_));
 AOI22_X4 _54798_ (.A1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2309]),
    .A2(_23097_),
    .B1(_23290_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1721]),
    .ZN(_23599_));
 BUF_X16 _54799_ (.A(_10940_),
    .Z(_23600_));
 AND3_X1 _54800_ (.A1(_10780_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2113]),
    .A3(_23600_),
    .ZN(_23601_));
 AND3_X1 _54801_ (.A1(_23207_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1966]),
    .A3(_10941_),
    .ZN(_23602_));
 NOR2_X2 _54802_ (.A1(_23601_),
    .A2(_23602_),
    .ZN(_23603_));
 BUF_X16 _54803_ (.A(_11019_),
    .Z(_23604_));
 AOI22_X2 _54804_ (.A1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2407]),
    .A2(_10922_),
    .B1(_23604_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1623]),
    .ZN(_23605_));
 AND4_X4 _54805_ (.A1(_23598_),
    .A2(_23599_),
    .A3(_23603_),
    .A4(_23605_),
    .ZN(_23606_));
 AOI22_X4 _54806_ (.A1(_10813_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3044]),
    .B1(_23490_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [55]),
    .ZN(_23607_));
 BUF_X8 _54807_ (.A(_22898_),
    .Z(_23608_));
 AND3_X4 _54808_ (.A1(_23367_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1378]),
    .A3(_23608_),
    .ZN(_23609_));
 BUF_X16 _54809_ (.A(_22733_),
    .Z(_23610_));
 AOI21_X4 _54810_ (.A(_23609_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [398]),
    .B2(_23610_),
    .ZN(_23611_));
 AOI22_X1 _54811_ (.A1(_23374_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2652]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [251]),
    .B2(_23446_),
    .ZN(_23612_));
 AOI22_X4 _54812_ (.A1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1280]),
    .A2(_23262_),
    .B1(_22827_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [104]),
    .ZN(_23613_));
 AND4_X1 _54813_ (.A1(_23607_),
    .A2(_23611_),
    .A3(_23612_),
    .A4(_23613_),
    .ZN(_23614_));
 BUF_X8 _54814_ (.A(_11170_),
    .Z(_23615_));
 AOI22_X4 _54815_ (.A1(_23615_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [349]),
    .B1(_23248_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [202]),
    .ZN(_23616_));
 AND3_X1 _54816_ (.A1(_22943_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1476]),
    .A3(_11036_),
    .ZN(_23617_));
 AOI21_X4 _54817_ (.A(_23617_),
    .B1(_23315_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1525]),
    .ZN(_23618_));
 AOI22_X4 _54818_ (.A1(_23092_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [692]),
    .B1(_23048_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1231]),
    .ZN(_23619_));
 AOI22_X4 _54819_ (.A1(_11206_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [6]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1427]),
    .B2(_23326_),
    .ZN(_23620_));
 NAND4_X4 _54820_ (.A1(_23616_),
    .A2(_23618_),
    .A3(_23619_),
    .A4(_23620_),
    .ZN(_23621_));
 BUF_X16 _54821_ (.A(_11146_),
    .Z(_23622_));
 AOI22_X4 _54822_ (.A1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1329]),
    .A2(_22282_),
    .B1(_23622_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [545]),
    .ZN(_23623_));
 AOI22_X4 _54823_ (.A1(_10839_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2946]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2995]),
    .B2(_10826_),
    .ZN(_23624_));
 BUF_X16 _54824_ (.A(_10874_),
    .Z(_23625_));
 AOI22_X4 _54825_ (.A1(_10800_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3093]),
    .B1(_23625_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2750]),
    .ZN(_23626_));
 BUF_X16 _54826_ (.A(_10902_),
    .Z(_23627_));
 AOI22_X4 _54827_ (.A1(_23373_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2701]),
    .B1(_23627_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2603]),
    .ZN(_23628_));
 NAND4_X2 _54828_ (.A1(_23623_),
    .A2(_23624_),
    .A3(_23626_),
    .A4(_23628_),
    .ZN(_23629_));
 AOI22_X4 _54829_ (.A1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2554]),
    .A2(_21654_),
    .B1(_10929_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2358]),
    .ZN(_23630_));
 AOI22_X4 _54830_ (.A1(_11196_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [153]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [300]),
    .B2(_22903_),
    .ZN(_23631_));
 BUF_X16 _54831_ (.A(_11090_),
    .Z(_23632_));
 AOI22_X4 _54832_ (.A1(_23331_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1133]),
    .B1(_23632_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1035]),
    .ZN(_23633_));
 AOI22_X4 _54833_ (.A1(_23267_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [790]),
    .B1(_23333_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1084]),
    .ZN(_23634_));
 NAND4_X4 _54834_ (.A1(_23630_),
    .A2(_23631_),
    .A3(_23633_),
    .A4(_23634_),
    .ZN(_23635_));
 AOI22_X4 _54835_ (.A1(_23047_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [937]),
    .B1(_22459_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [986]),
    .ZN(_23636_));
 AOI22_X2 _54836_ (.A1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1182]),
    .A2(_23325_),
    .B1(_23106_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [594]),
    .ZN(_23637_));
 BUF_X16 _54837_ (.A(_22597_),
    .Z(_23638_));
 AOI22_X4 _54838_ (.A1(_23638_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [741]),
    .B1(_23107_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [643]),
    .ZN(_23639_));
 AOI22_X4 _54839_ (.A1(_11153_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [496]),
    .B1(_11159_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [447]),
    .ZN(_23640_));
 NAND4_X4 _54840_ (.A1(_23636_),
    .A2(_23637_),
    .A3(_23639_),
    .A4(_23640_),
    .ZN(_23641_));
 NOR4_X2 _54841_ (.A1(_23621_),
    .A2(_23629_),
    .A3(_23635_),
    .A4(_23641_),
    .ZN(_23642_));
 NAND4_X2 _54842_ (.A1(_23597_),
    .A2(_23606_),
    .A3(_23614_),
    .A4(_23642_),
    .ZN(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [6]));
 BUF_X16 _54843_ (.A(_11173_),
    .Z(_23643_));
 AND3_X1 _54844_ (.A1(_23288_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [105]),
    .A3(_23643_),
    .ZN(_23644_));
 AOI221_X4 _54845_ (.A(_23644_),
    .B1(_11205_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [7]),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [154]),
    .C2(_11196_),
    .ZN(_23645_));
 NAND3_X1 _54846_ (.A1(_23215_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [252]),
    .A3(_22937_),
    .ZN(_23646_));
 OAI221_X2 _54847_ (.A(_23646_),
    .B1(_11182_),
    .B2(_22765_),
    .C1(_11171_),
    .C2(_22751_),
    .ZN(_23647_));
 AOI221_X2 _54848_ (.A(_23647_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [203]),
    .B2(_11190_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [56]),
    .C2(_23490_),
    .ZN(_23648_));
 AND3_X1 _54849_ (.A1(_23284_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1134]),
    .A3(_23494_),
    .ZN(_23649_));
 AOI221_X2 _54850_ (.A(_23649_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1085]),
    .B2(_22410_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1036]),
    .C2(_23632_),
    .ZN(_23650_));
 AOI22_X4 _54851_ (.A1(_22459_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [987]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [840]),
    .B2(_23268_),
    .ZN(_23651_));
 AND4_X4 _54852_ (.A1(_23645_),
    .A2(_23648_),
    .A3(net53),
    .A4(_23651_),
    .ZN(_23652_));
 NAND3_X1 _54853_ (.A1(_23215_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1820]),
    .A3(_23402_),
    .ZN(_23653_));
 OAI221_X2 _54854_ (.A(_23653_),
    .B1(_10994_),
    .B2(_22011_),
    .C1(_10984_),
    .C2(_21987_),
    .ZN(_23654_));
 AOI221_X4 _54855_ (.A(_23654_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1771]),
    .B2(_11002_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1624]),
    .C2(_23396_),
    .ZN(_23655_));
 NAND3_X1 _54856_ (.A1(_23284_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2310]),
    .A3(_22913_),
    .ZN(_23656_));
 BUF_X8 _54857_ (.A(_10935_),
    .Z(_23657_));
 NAND3_X1 _54858_ (.A1(_22942_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2261]),
    .A3(_23657_),
    .ZN(_23658_));
 NAND2_X1 _54859_ (.A1(_23656_),
    .A2(_23658_),
    .ZN(_23659_));
 BUF_X16 _54860_ (.A(_10955_),
    .Z(_23660_));
 AOI221_X2 _54861_ (.A(_23659_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2212]),
    .B2(_10950_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2163]),
    .C2(_23660_),
    .ZN(_23661_));
 BUF_X8 _54862_ (.A(_10987_),
    .Z(_23662_));
 AND3_X1 _54863_ (.A1(_23173_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1673]),
    .A3(_23662_),
    .ZN(_23663_));
 AOI221_X4 _54864_ (.A(_23663_),
    .B1(_11025_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1575]),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1722]),
    .C2(_22078_),
    .ZN(_23664_));
 NAND3_X1 _54865_ (.A1(_10877_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1967]),
    .A3(_10939_),
    .ZN(_23665_));
 OAI21_X1 _54866_ (.A(_23665_),
    .B1(_10973_),
    .B2(_21943_),
    .ZN(_23666_));
 AOI221_X4 _54867_ (.A(_23666_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2114]),
    .B2(_10961_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2065]),
    .C2(_21900_),
    .ZN(_23667_));
 AND4_X4 _54868_ (.A1(_23655_),
    .A2(_23661_),
    .A3(_23664_),
    .A4(_23667_),
    .ZN(_23668_));
 BUF_X8 _54869_ (.A(_10886_),
    .Z(_23669_));
 NAND3_X1 _54870_ (.A1(_23309_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2555]),
    .A3(_23669_),
    .ZN(_23670_));
 OAI221_X2 _54871_ (.A(_23670_),
    .B1(_10897_),
    .B2(_21613_),
    .C1(_10888_),
    .C2(_21584_),
    .ZN(_23671_));
 AOI221_X4 _54872_ (.A(_23671_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2604]),
    .B2(_23627_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2408]),
    .C2(_10922_),
    .ZN(_23672_));
 BUF_X16 _54873_ (.A(_22928_),
    .Z(_23673_));
 NAND3_X1 _54874_ (.A1(_23434_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2996]),
    .A3(_23673_),
    .ZN(_23674_));
 AOI22_X2 _54875_ (.A1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2751]),
    .A2(_23625_),
    .B1(_22918_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2947]),
    .ZN(_23675_));
 NAND3_X1 _54876_ (.A1(_23240_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3045]),
    .A3(_23360_),
    .ZN(_23676_));
 NAND3_X1 _54877_ (.A1(_23245_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3094]),
    .A3(_23360_),
    .ZN(_23677_));
 AND4_X4 _54878_ (.A1(_23674_),
    .A2(_23675_),
    .A3(_23676_),
    .A4(_23677_),
    .ZN(_23678_));
 NAND3_X1 _54879_ (.A1(_10868_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2800]),
    .A3(_23673_),
    .ZN(_23679_));
 AND3_X1 _54880_ (.A1(_10855_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2457]),
    .A3(_10886_),
    .ZN(_23680_));
 AOI221_X2 _54881_ (.A(_23680_),
    .B1(_10928_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2359]),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2506]),
    .C2(_10912_),
    .ZN(_23681_));
 NAND3_X1 _54882_ (.A1(_10780_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2898]),
    .A3(_23360_),
    .ZN(_23682_));
 NAND3_X1 _54883_ (.A1(_22523_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2849]),
    .A3(_22990_),
    .ZN(_23683_));
 AND4_X1 _54884_ (.A1(_23679_),
    .A2(_23681_),
    .A3(_23682_),
    .A4(_23683_),
    .ZN(_23684_));
 AND3_X4 _54885_ (.A1(_23672_),
    .A2(_23678_),
    .A3(_23684_),
    .ZN(_23685_));
 NAND3_X1 _54886_ (.A1(_23385_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [644]),
    .A3(_23237_),
    .ZN(_23686_));
 AND3_X1 _54887_ (.A1(_10797_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [742]),
    .A3(_11145_),
    .ZN(_23687_));
 AOI221_X2 _54888_ (.A(_23687_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [693]),
    .B2(_11130_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [595]),
    .C2(_11141_),
    .ZN(_23688_));
 BUF_X8 _54889_ (.A(_11151_),
    .Z(_23689_));
 AOI22_X1 _54890_ (.A1(_11147_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [546]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [497]),
    .B2(_23689_),
    .ZN(_23690_));
 AOI22_X2 _54891_ (.A1(_22733_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [399]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [448]),
    .B2(_11158_),
    .ZN(_23691_));
 AND4_X2 _54892_ (.A1(_23686_),
    .A2(_23688_),
    .A3(_23690_),
    .A4(_23691_),
    .ZN(_23692_));
 BUF_X4 _54893_ (.A(_22898_),
    .Z(_23693_));
 NAND3_X1 _54894_ (.A1(_23385_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1428]),
    .A3(_23693_),
    .ZN(_23694_));
 NAND3_X1 _54895_ (.A1(_10804_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1526]),
    .A3(_23050_),
    .ZN(_23695_));
 NAND3_X1 _54896_ (.A1(_23367_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1379]),
    .A3(_23608_),
    .ZN(_23696_));
 NAND3_X1 _54897_ (.A1(_10818_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1477]),
    .A3(_23608_),
    .ZN(_23697_));
 AND4_X4 _54898_ (.A1(_23694_),
    .A2(_23695_),
    .A3(_23696_),
    .A4(_23697_),
    .ZN(_23698_));
 AND3_X1 _54899_ (.A1(_23083_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [791]),
    .A3(_23460_),
    .ZN(_23699_));
 AOI221_X4 _54900_ (.A(_23699_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [889]),
    .B2(_11106_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [938]),
    .C2(_11100_),
    .ZN(_23700_));
 BUF_X8 _54901_ (.A(_11034_),
    .Z(_23701_));
 NAND3_X1 _54902_ (.A1(_23166_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1330]),
    .A3(_23701_),
    .ZN(_23702_));
 NAND3_X1 _54903_ (.A1(_22521_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1281]),
    .A3(_23701_),
    .ZN(_23703_));
 NAND2_X2 _54904_ (.A1(_23702_),
    .A2(_23703_),
    .ZN(_23704_));
 AOI221_X2 _54905_ (.A(_23704_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1232]),
    .B2(_11065_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1183]),
    .C2(_23103_),
    .ZN(_23705_));
 AND4_X4 _54906_ (.A1(_23692_),
    .A2(_23698_),
    .A3(_23700_),
    .A4(_23705_),
    .ZN(_23706_));
 NAND4_X1 _54907_ (.A1(_23652_),
    .A2(_23668_),
    .A3(_23685_),
    .A4(_23706_),
    .ZN(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [7]));
 AND3_X1 _54908_ (.A1(_23288_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [498]),
    .A3(_23504_),
    .ZN(_23707_));
 AOI221_X4 _54909_ (.A(_23707_),
    .B1(_22733_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [400]),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [547]),
    .C2(_23622_),
    .ZN(_23708_));
 BUF_X8 _54910_ (.A(_22938_),
    .Z(_23709_));
 NAND3_X1 _54911_ (.A1(_23221_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [204]),
    .A3(_23709_),
    .ZN(_23710_));
 AND3_X1 _54912_ (.A1(_10797_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [351]),
    .A3(_11173_),
    .ZN(_23711_));
 AOI221_X2 _54913_ (.A(_23711_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [302]),
    .B2(_11181_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [253]),
    .C2(_11186_),
    .ZN(_23712_));
 AOI22_X2 _54914_ (.A1(_11196_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [155]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [106]),
    .B2(_23453_),
    .ZN(_23713_));
 BUF_X16 _54915_ (.A(_11211_),
    .Z(_23714_));
 AOI22_X2 _54916_ (.A1(_23164_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [8]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [57]),
    .B2(_23714_),
    .ZN(_23715_));
 AND4_X4 _54917_ (.A1(_23710_),
    .A2(_23712_),
    .A3(_23713_),
    .A4(_23715_),
    .ZN(_23716_));
 AND3_X1 _54918_ (.A1(_22942_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [694]),
    .A3(_23512_),
    .ZN(_23717_));
 AOI221_X4 _54919_ (.A(_23717_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [645]),
    .B2(_22642_),
    .C1(_23638_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [743]),
    .ZN(_23718_));
 AOI22_X2 _54920_ (.A1(_23106_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [596]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [449]),
    .B2(_11159_),
    .ZN(_23719_));
 AND4_X4 _54921_ (.A1(_23708_),
    .A2(_23716_),
    .A3(_23718_),
    .A4(_23719_),
    .ZN(_23720_));
 BUF_X32 _54922_ (.A(_10855_),
    .Z(_23721_));
 AND3_X1 _54923_ (.A1(_23721_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2850]),
    .A3(_23498_),
    .ZN(_23722_));
 AOI221_X4 _54924_ (.A(_23722_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2801]),
    .B2(_10863_),
    .C1(_23213_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2899]),
    .ZN(_23723_));
 NAND3_X1 _54925_ (.A1(_23459_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2311]),
    .A3(_23169_),
    .ZN(_23724_));
 OAI21_X1 _54926_ (.A(_23724_),
    .B1(_10946_),
    .B2(_21830_),
    .ZN(_23725_));
 AOI221_X2 _54927_ (.A(_23725_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2213]),
    .B2(_10950_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2164]),
    .C2(_23660_),
    .ZN(_23726_));
 NAND3_X1 _54928_ (.A1(_23339_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2948]),
    .A3(_22990_),
    .ZN(_23727_));
 AOI22_X2 _54929_ (.A1(_23224_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3095]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3046]),
    .B2(_23225_),
    .ZN(_23728_));
 NAND3_X1 _54930_ (.A1(_10879_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2752]),
    .A3(_22999_),
    .ZN(_23729_));
 NAND3_X1 _54931_ (.A1(_23252_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2997]),
    .A3(_23122_),
    .ZN(_23730_));
 AND4_X4 _54932_ (.A1(_23727_),
    .A2(_23728_),
    .A3(_23729_),
    .A4(_23730_),
    .ZN(_23731_));
 NAND3_X1 _54933_ (.A1(_23230_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1968]),
    .A3(_22962_),
    .ZN(_23732_));
 BUF_X32 _54934_ (.A(_10920_),
    .Z(_23733_));
 NAND3_X1 _54935_ (.A1(_23733_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2017]),
    .A3(_23169_),
    .ZN(_23734_));
 NAND2_X1 _54936_ (.A1(_23732_),
    .A2(_23734_),
    .ZN(_23735_));
 BUF_X16 _54937_ (.A(_10961_),
    .Z(_23736_));
 AOI221_X4 _54938_ (.A(_23735_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2066]),
    .B2(_23233_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2115]),
    .C2(_23736_),
    .ZN(_23737_));
 AND4_X1 _54939_ (.A1(_23723_),
    .A2(_23726_),
    .A3(_23731_),
    .A4(_23737_),
    .ZN(_23738_));
 OAI22_X2 _54940_ (.A1(_22259_),
    .A2(_11051_),
    .B1(_11070_),
    .B2(_22367_),
    .ZN(_23739_));
 OAI22_X4 _54941_ (.A1(_11032_),
    .A2(_22193_),
    .B1(_22219_),
    .B2(_11042_),
    .ZN(_23740_));
 AOI211_X2 _54942_ (.A(_23739_),
    .B(_23740_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1429]),
    .C2(_23326_),
    .ZN(_23741_));
 OAI22_X4 _54943_ (.A1(_22445_),
    .A2(_11091_),
    .B1(_11111_),
    .B2(_22555_),
    .ZN(_23742_));
 OAI22_X2 _54944_ (.A1(_11076_),
    .A2(_22394_),
    .B1(_22419_),
    .B2(_11086_),
    .ZN(_23743_));
 AOI211_X2 _54945_ (.A(_23742_),
    .B(_23743_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [988]),
    .C2(_22459_),
    .ZN(_23744_));
 AND3_X1 _54946_ (.A1(_23083_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [792]),
    .A3(_23460_),
    .ZN(_23745_));
 AOI221_X4 _54947_ (.A(_23745_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [890]),
    .B2(_11106_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [939]),
    .C2(_11100_),
    .ZN(_23746_));
 AND3_X1 _54948_ (.A1(_23176_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1233]),
    .A3(_22979_),
    .ZN(_23747_));
 BUF_X8 _54949_ (.A(_11054_),
    .Z(_23748_));
 AOI221_X4 _54950_ (.A(_23747_),
    .B1(_11059_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1282]),
    .C1(_23748_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1331]),
    .ZN(_23749_));
 AND4_X4 _54951_ (.A1(_23741_),
    .A2(_23744_),
    .A3(_23746_),
    .A4(_23749_),
    .ZN(_23750_));
 BUF_X32 _54952_ (.A(_10811_),
    .Z(_23751_));
 AND3_X1 _54953_ (.A1(_23751_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1870]),
    .A3(_22923_),
    .ZN(_23752_));
 AOI221_X4 _54954_ (.A(_23752_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1821]),
    .B2(_23286_),
    .C1(_23584_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1919]),
    .ZN(_23753_));
 NAND3_X1 _54955_ (.A1(_10780_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2507]),
    .A3(_23427_),
    .ZN(_23754_));
 AOI22_X2 _54956_ (.A1(_10929_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2360]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2409]),
    .B2(_23301_),
    .ZN(_23755_));
 NAND3_X1 _54957_ (.A1(_22523_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2458]),
    .A3(_23119_),
    .ZN(_23756_));
 BUF_X32 _54958_ (.A(_22240_),
    .Z(_23757_));
 NAND3_X1 _54959_ (.A1(_23757_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2605]),
    .A3(_23119_),
    .ZN(_23758_));
 AND4_X1 _54960_ (.A1(_23754_),
    .A2(_23755_),
    .A3(_23756_),
    .A4(_23758_),
    .ZN(_23759_));
 AOI22_X4 _54961_ (.A1(_23290_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1723]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1674]),
    .B2(_22105_),
    .ZN(_23760_));
 NAND3_X1 _54962_ (.A1(_23339_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1772]),
    .A3(_23393_),
    .ZN(_23761_));
 AOI22_X2 _54963_ (.A1(_23595_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1576]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1625]),
    .B2(_23396_),
    .ZN(_23762_));
 AND3_X4 _54964_ (.A1(_23760_),
    .A2(_23761_),
    .A3(_23762_),
    .ZN(_23763_));
 AND3_X1 _54965_ (.A1(_23309_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2556]),
    .A3(_23310_),
    .ZN(_23764_));
 AOI221_X2 _54966_ (.A(_23764_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2654]),
    .B2(_21601_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2703]),
    .C2(_21573_),
    .ZN(_23765_));
 AND4_X4 _54967_ (.A1(_23753_),
    .A2(_23759_),
    .A3(_23763_),
    .A4(_23765_),
    .ZN(_23766_));
 NAND4_X2 _54968_ (.A1(_23720_),
    .A2(_23738_),
    .A3(_23750_),
    .A4(_23766_),
    .ZN(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [8]));
 NAND3_X1 _54969_ (.A1(_22897_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [744]),
    .A3(_23055_),
    .ZN(_23767_));
 NAND3_X1 _54970_ (.A1(_10878_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [401]),
    .A3(_23055_),
    .ZN(_23768_));
 NAND2_X1 _54971_ (.A1(_23767_),
    .A2(_23768_),
    .ZN(_23769_));
 AOI221_X4 _54972_ (.A(_23769_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [646]),
    .B2(_23107_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [597]),
    .C2(_23106_),
    .ZN(_23770_));
 NAND3_X4 _54973_ (.A1(_23158_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [548]),
    .A3(_23161_),
    .ZN(_23771_));
 OAI21_X4 _54974_ (.A(_23771_),
    .B1(_10917_),
    .B2(_21713_),
    .ZN(_23772_));
 AOI221_X4 _54975_ (.A(_23772_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2116]),
    .B2(_23736_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2067]),
    .C2(_21900_),
    .ZN(_23773_));
 NAND3_X2 _54976_ (.A1(_22920_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [695]),
    .A3(_23151_),
    .ZN(_23774_));
 BUF_X32 _54977_ (.A(_10866_),
    .Z(_23775_));
 NAND3_X2 _54978_ (.A1(_23775_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [450]),
    .A3(_23510_),
    .ZN(_23776_));
 NAND2_X4 _54979_ (.A1(_23774_),
    .A2(_23776_),
    .ZN(_23777_));
 AOI221_X4 _54980_ (.A(_23777_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2998]),
    .B2(_10826_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [499]),
    .C2(_11153_),
    .ZN(_23778_));
 NAND3_X2 _54981_ (.A1(_22953_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1724]),
    .A3(_22921_),
    .ZN(_23779_));
 NAND3_X1 _54982_ (.A1(_23775_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2018]),
    .A3(_23657_),
    .ZN(_23780_));
 NAND2_X2 _54983_ (.A1(_23779_),
    .A2(_23780_),
    .ZN(_23781_));
 AOI221_X2 _54984_ (.A(_23781_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2361]),
    .B2(_23300_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1577]),
    .C2(_23395_),
    .ZN(_23782_));
 AND4_X1 _54985_ (.A1(_23770_),
    .A2(_23773_),
    .A3(_23778_),
    .A4(net37),
    .ZN(_23783_));
 NAND3_X1 _54986_ (.A1(_23487_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2704]),
    .A3(_23012_),
    .ZN(_23784_));
 OAI21_X1 _54987_ (.A(_23784_),
    .B1(_10897_),
    .B2(_21615_),
    .ZN(_23785_));
 AOI221_X2 _54988_ (.A(_23785_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2606]),
    .B2(_10902_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2214]),
    .C2(_10950_),
    .ZN(_23786_));
 NAND3_X1 _54989_ (.A1(_10778_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [156]),
    .A3(_22937_),
    .ZN(_23787_));
 OAI21_X1 _54990_ (.A(_23787_),
    .B1(_11201_),
    .B2(_22839_),
    .ZN(_23788_));
 AOI221_X4 _54991_ (.A(_23788_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2753]),
    .B2(_21289_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3047]),
    .C2(_10813_),
    .ZN(_23789_));
 NAND3_X2 _54992_ (.A1(_23518_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2165]),
    .A3(_23231_),
    .ZN(_23790_));
 NAND3_X4 _54993_ (.A1(_23518_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2557]),
    .A3(_23012_),
    .ZN(_23791_));
 NAND2_X4 _54994_ (.A1(_23790_),
    .A2(_23791_),
    .ZN(_23792_));
 AOI221_X4 _54995_ (.A(_23792_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1479]),
    .B2(_22210_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1430]),
    .C2(_23326_),
    .ZN(_23793_));
 BUF_X8 _54996_ (.A(_10787_),
    .Z(_23794_));
 NAND3_X1 _54997_ (.A1(_10856_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2851]),
    .A3(_23794_),
    .ZN(_23795_));
 NAND3_X1 _54998_ (.A1(_23733_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2802]),
    .A3(_23174_),
    .ZN(_23796_));
 NAND2_X1 _54999_ (.A1(_23795_),
    .A2(_23796_),
    .ZN(_23797_));
 AOI221_X4 _55000_ (.A(_23797_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1675]),
    .B2(_11012_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2949]),
    .C2(_22918_),
    .ZN(_23798_));
 AND4_X1 _55001_ (.A1(_23786_),
    .A2(_23789_),
    .A3(_23793_),
    .A4(_23798_),
    .ZN(_23799_));
 NAND3_X1 _55002_ (.A1(_22953_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1332]),
    .A3(_11035_),
    .ZN(_23800_));
 NAND3_X2 _55003_ (.A1(_22915_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1234]),
    .A3(_11035_),
    .ZN(_23801_));
 NAND2_X1 _55004_ (.A1(_23800_),
    .A2(_23801_),
    .ZN(_23802_));
 AOI221_X4 _55005_ (.A(_23802_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2312]),
    .B2(_10936_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [891]),
    .C2(_23265_),
    .ZN(_23803_));
 BUF_X8 _55006_ (.A(_11079_),
    .Z(_23804_));
 NAND3_X1 _55007_ (.A1(_23158_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [940]),
    .A3(_23804_),
    .ZN(_23805_));
 BUF_X32 _55008_ (.A(_10920_),
    .Z(_23806_));
 NAND3_X1 _55009_ (.A1(_23806_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [842]),
    .A3(_23804_),
    .ZN(_23807_));
 NAND2_X1 _55010_ (.A1(_23805_),
    .A2(_23807_),
    .ZN(_23808_));
 AOI221_X4 _55011_ (.A(_23808_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1038]),
    .B2(_22435_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [793]),
    .C2(_11114_),
    .ZN(_23809_));
 BUF_X32 _55012_ (.A(_22896_),
    .Z(_23810_));
 NAND3_X2 _55013_ (.A1(_23810_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1920]),
    .A3(_23662_),
    .ZN(_23811_));
 NAND3_X2 _55014_ (.A1(_23168_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1822]),
    .A3(_23662_),
    .ZN(_23812_));
 NAND2_X4 _55015_ (.A1(_23811_),
    .A2(_23812_),
    .ZN(_23813_));
 AOI221_X2 _55016_ (.A(_23813_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1626]),
    .B2(_11019_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1283]),
    .C2(_23262_),
    .ZN(_23814_));
 NAND3_X1 _55017_ (.A1(_23810_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [352]),
    .A3(_23258_),
    .ZN(_23815_));
 NAND3_X4 _55018_ (.A1(_23408_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1871]),
    .A3(_23402_),
    .ZN(_23816_));
 NAND2_X1 _55019_ (.A1(_23815_),
    .A2(_23816_),
    .ZN(_23817_));
 AOI221_X2 _55020_ (.A(_23817_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1185]),
    .B2(_11069_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [254]),
    .C2(_23446_),
    .ZN(_23818_));
 AND4_X4 _55021_ (.A1(_23803_),
    .A2(_23809_),
    .A3(_23814_),
    .A4(_23818_),
    .ZN(_23819_));
 AND3_X1 _55022_ (.A1(_10803_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1136]),
    .A3(_11080_),
    .ZN(_23820_));
 AOI21_X4 _55023_ (.A(_23820_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1087]),
    .B2(_23333_),
    .ZN(_23821_));
 OAI221_X2 _55024_ (.A(_23821_),
    .B1(_21397_),
    .B2(_10801_),
    .C1(_21472_),
    .C2(_10774_),
    .ZN(_23822_));
 NAND3_X4 _55025_ (.A1(_23054_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1528]),
    .A3(_22945_),
    .ZN(_23823_));
 NAND3_X4 _55026_ (.A1(_22944_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [303]),
    .A3(_22951_),
    .ZN(_23824_));
 NAND3_X2 _55027_ (.A1(_23062_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2410]),
    .A3(_23014_),
    .ZN(_23825_));
 NAND3_X4 _55028_ (.A1(_23192_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1381]),
    .A3(_23566_),
    .ZN(_23826_));
 NAND4_X4 _55029_ (.A1(_23823_),
    .A2(_23824_),
    .A3(_23825_),
    .A4(_23826_),
    .ZN(_23827_));
 NAND3_X2 _55030_ (.A1(_22955_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2508]),
    .A3(_23068_),
    .ZN(_23828_));
 NAND3_X2 _55031_ (.A1(_22972_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2263]),
    .A3(_22964_),
    .ZN(_23829_));
 BUF_X16 _55032_ (.A(_22934_),
    .Z(_23830_));
 NAND3_X2 _55033_ (.A1(_23271_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1773]),
    .A3(_23830_),
    .ZN(_23831_));
 BUF_X8 _55034_ (.A(_22963_),
    .Z(_23832_));
 NAND3_X2 _55035_ (.A1(_23085_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1969]),
    .A3(_23832_),
    .ZN(_23833_));
 NAND4_X4 _55036_ (.A1(_23828_),
    .A2(_23829_),
    .A3(_23831_),
    .A4(_23833_),
    .ZN(_23834_));
 BUF_X8 _55037_ (.A(_11175_),
    .Z(_23835_));
 NAND3_X1 _55038_ (.A1(_10844_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [205]),
    .A3(_23835_),
    .ZN(_23836_));
 BUF_X16 _55039_ (.A(_23084_),
    .Z(_23837_));
 NAND3_X2 _55040_ (.A1(_23837_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [9]),
    .A3(_23196_),
    .ZN(_23838_));
 BUF_X32 _55041_ (.A(_10843_),
    .Z(_23839_));
 NAND3_X4 _55042_ (.A1(_23839_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [989]),
    .A3(_23547_),
    .ZN(_23840_));
 NAND3_X2 _55043_ (.A1(_23426_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [58]),
    .A3(_23086_),
    .ZN(_23841_));
 NAND4_X4 _55044_ (.A1(_23836_),
    .A2(_23838_),
    .A3(_23840_),
    .A4(_23841_),
    .ZN(_23842_));
 NOR4_X2 _55045_ (.A1(_23822_),
    .A2(_23827_),
    .A3(_23834_),
    .A4(_23842_),
    .ZN(_23843_));
 NAND4_X1 _55046_ (.A1(_23783_),
    .A2(_23799_),
    .A3(_23819_),
    .A4(_23843_),
    .ZN(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [9]));
 NAND3_X1 _55047_ (.A1(_10878_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1186]),
    .A3(_22898_),
    .ZN(_23844_));
 NAND3_X4 _55048_ (.A1(_22240_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1431]),
    .A3(_22898_),
    .ZN(_23845_));
 NAND2_X4 _55049_ (.A1(_23844_),
    .A2(_23845_),
    .ZN(_23846_));
 AOI221_X4 _55050_ (.A(_23846_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [647]),
    .B2(_23107_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [745]),
    .C2(_23638_),
    .ZN(_23847_));
 BUF_X16 _55051_ (.A(_11034_),
    .Z(_23848_));
 NAND3_X1 _55052_ (.A1(_23166_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1333]),
    .A3(_23848_),
    .ZN(_23849_));
 OAI21_X2 _55053_ (.A(_23849_),
    .B1(_11051_),
    .B2(_22263_),
    .ZN(_23850_));
 AOI221_X4 _55054_ (.A(_23850_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1529]),
    .B2(_23179_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1480]),
    .C2(_23095_),
    .ZN(_23851_));
 NAND3_X1 _55055_ (.A1(_23733_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2411]),
    .A3(_23669_),
    .ZN(_23852_));
 OAI21_X1 _55056_ (.A(_23852_),
    .B1(_10903_),
    .B2(_21638_),
    .ZN(_23853_));
 AOI221_X4 _55057_ (.A(_23853_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2460]),
    .B2(_21705_),
    .C1(net1392),
    .C2(_23092_),
    .ZN(_23854_));
 NAND3_X4 _55058_ (.A1(_22915_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [451]),
    .A3(_23151_),
    .ZN(_23855_));
 NAND3_X1 _55059_ (.A1(_23775_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2803]),
    .A3(_23498_),
    .ZN(_23856_));
 NAND2_X1 _55060_ (.A1(_23855_),
    .A2(_23856_),
    .ZN(_23857_));
 AOI221_X4 _55061_ (.A(_23857_),
    .B1(_23300_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2362]),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2901]),
    .C2(_21466_),
    .ZN(_23858_));
 AND4_X1 _55062_ (.A1(_23847_),
    .A2(_23851_),
    .A3(_23854_),
    .A4(_23858_),
    .ZN(_23859_));
 NAND3_X1 _55063_ (.A1(_23487_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1921]),
    .A3(_23519_),
    .ZN(_23860_));
 OAI21_X4 _55064_ (.A(_23860_),
    .B1(_10994_),
    .B2(_22015_),
    .ZN(_23861_));
 AOI221_X2 _55065_ (.A(_23861_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1774]),
    .B2(_11002_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1235]),
    .C2(_23048_),
    .ZN(_23862_));
 NAND3_X1 _55066_ (.A1(_23509_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [549]),
    .A3(_23510_),
    .ZN(_23863_));
 NAND3_X2 _55067_ (.A1(_23153_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [598]),
    .A3(_23512_),
    .ZN(_23864_));
 NAND2_X4 _55068_ (.A1(_23863_),
    .A2(_23864_),
    .ZN(_23865_));
 AOI221_X4 _55069_ (.A(_23865_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1823]),
    .B2(_22044_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1284]),
    .C2(_23262_),
    .ZN(_23866_));
 NAND3_X1 _55070_ (.A1(_23487_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2705]),
    .A3(_23481_),
    .ZN(_23867_));
 NAND3_X4 _55071_ (.A1(_23230_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2754]),
    .A3(_23794_),
    .ZN(_23868_));
 NAND2_X1 _55072_ (.A1(_23867_),
    .A2(_23868_),
    .ZN(_23869_));
 AOI221_X2 _55073_ (.A(_23869_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2656]),
    .B2(_21601_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2068]),
    .C2(_21900_),
    .ZN(_23870_));
 NAND3_X4 _55074_ (.A1(_23810_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [353]),
    .A3(_23258_),
    .ZN(_23871_));
 NAND3_X2 _55075_ (.A1(_23518_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [206]),
    .A3(_23258_),
    .ZN(_23872_));
 NAND2_X4 _55076_ (.A1(_23871_),
    .A2(_23872_),
    .ZN(_23873_));
 AOI221_X2 _55077_ (.A(_23873_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3048]),
    .B2(_10812_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2999]),
    .C2(_10826_),
    .ZN(_23874_));
 AND4_X2 _55078_ (.A1(_23862_),
    .A2(_23866_),
    .A3(_23870_),
    .A4(net36),
    .ZN(_23875_));
 AND3_X1 _55079_ (.A1(_10817_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2264]),
    .A3(_22963_),
    .ZN(_23876_));
 AOI21_X4 _55080_ (.A(_23876_),
    .B1(_23097_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2313]),
    .ZN(_23877_));
 OAI221_X2 _55081_ (.A(_23877_),
    .B1(_22117_),
    .B2(_11013_),
    .C1(_22396_),
    .C2(_11076_),
    .ZN(_23878_));
 BUF_X8 _55082_ (.A(_11080_),
    .Z(_23879_));
 BUF_X8 _55083_ (.A(_23879_),
    .Z(_23880_));
 NAND3_X1 _55084_ (.A1(_23004_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [941]),
    .A3(_23880_),
    .ZN(_23881_));
 BUF_X8 _55085_ (.A(_22969_),
    .Z(_23882_));
 NAND3_X2 _55086_ (.A1(_23377_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [843]),
    .A3(_23882_),
    .ZN(_23883_));
 NAND3_X2 _55087_ (.A1(_10858_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [892]),
    .A3(_23882_),
    .ZN(_23884_));
 NAND3_X2 _55088_ (.A1(_22968_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [794]),
    .A3(_22970_),
    .ZN(_23885_));
 NAND4_X4 _55089_ (.A1(_23881_),
    .A2(_23883_),
    .A3(_23884_),
    .A4(_23885_),
    .ZN(_23886_));
 NAND3_X4 _55090_ (.A1(_23560_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3097]),
    .A3(_23128_),
    .ZN(_23887_));
 BUF_X32 _55091_ (.A(_22943_),
    .Z(_23888_));
 NAND3_X2 _55092_ (.A1(_23888_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1088]),
    .A3(_22973_),
    .ZN(_23889_));
 NAND3_X2 _55093_ (.A1(_23276_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [990]),
    .A3(_22976_),
    .ZN(_23890_));
 BUF_X8 _55094_ (.A(_22969_),
    .Z(_23891_));
 NAND3_X2 _55095_ (.A1(_23071_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1039]),
    .A3(_23891_),
    .ZN(_23892_));
 NAND4_X4 _55096_ (.A1(_23887_),
    .A2(_23889_),
    .A3(_23890_),
    .A4(_23892_),
    .ZN(_23893_));
 BUF_X8 _55097_ (.A(_22963_),
    .Z(_23894_));
 NAND3_X2 _55098_ (.A1(_22955_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2117]),
    .A3(_23894_),
    .ZN(_23895_));
 NAND3_X2 _55099_ (.A1(_23276_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2166]),
    .A3(_23832_),
    .ZN(_23896_));
 NAND3_X2 _55100_ (.A1(_23080_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2215]),
    .A3(_23081_),
    .ZN(_23897_));
 NAND3_X4 _55101_ (.A1(_23042_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1627]),
    .A3(_23576_),
    .ZN(_23898_));
 NAND4_X4 _55102_ (.A1(_23895_),
    .A2(_23896_),
    .A3(_23897_),
    .A4(_23898_),
    .ZN(_23899_));
 NOR4_X2 _55103_ (.A1(_23878_),
    .A2(_23886_),
    .A3(_23893_),
    .A4(_23899_),
    .ZN(_23900_));
 AND3_X1 _55104_ (.A1(_23035_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [59]),
    .A3(_22938_),
    .ZN(_23901_));
 AOI21_X4 _55105_ (.A(_23901_),
    .B1(_11206_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [10]),
    .ZN(_23902_));
 OAI221_X2 _55106_ (.A(_23902_),
    .B1(_10840_),
    .B2(_21448_),
    .C1(_21661_),
    .C2(_10908_),
    .ZN(_23903_));
 AOI22_X4 _55107_ (.A1(_22903_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [304]),
    .B1(_23446_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [255]),
    .ZN(_23904_));
 NAND3_X2 _55108_ (.A1(_23016_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [108]),
    .A3(_11176_),
    .ZN(_23905_));
 OAI211_X4 _55109_ (.A(_23904_),
    .B(_23905_),
    .C1(_11197_),
    .C2(_22814_),
    .ZN(_23906_));
 NAND3_X4 _55110_ (.A1(_23133_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1578]),
    .A3(_22956_),
    .ZN(_23907_));
 NAND3_X4 _55111_ (.A1(_23194_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [402]),
    .A3(_23201_),
    .ZN(_23908_));
 NAND3_X1 _55112_ (.A1(_23078_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2852]),
    .A3(_23037_),
    .ZN(_23909_));
 NAND3_X4 _55113_ (.A1(_23039_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [500]),
    .A3(_23072_),
    .ZN(_23910_));
 NAND4_X1 _55114_ (.A1(_23907_),
    .A2(_23908_),
    .A3(_23909_),
    .A4(_23910_),
    .ZN(_23911_));
 NAND3_X2 _55115_ (.A1(_23200_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1725]),
    .A3(_23141_),
    .ZN(_23912_));
 NAND3_X4 _55116_ (.A1(_23421_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2509]),
    .A3(_23029_),
    .ZN(_23913_));
 NAND3_X2 _55117_ (.A1(_23042_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2019]),
    .A3(_23081_),
    .ZN(_23914_));
 NAND3_X2 _55118_ (.A1(_23207_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1970]),
    .A3(_23600_),
    .ZN(_23915_));
 NAND4_X4 _55119_ (.A1(_23912_),
    .A2(_23913_),
    .A3(_23914_),
    .A4(_23915_),
    .ZN(_23916_));
 NOR4_X1 _55120_ (.A1(_23903_),
    .A2(_23906_),
    .A3(_23911_),
    .A4(_23916_),
    .ZN(_23917_));
 NAND4_X1 _55121_ (.A1(_23859_),
    .A2(_23875_),
    .A3(_23900_),
    .A4(_23917_),
    .ZN(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [10]));
 NAND3_X1 _55122_ (.A1(_23524_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [697]),
    .A3(_23255_),
    .ZN(_23918_));
 OAI221_X2 _55123_ (.A(_23918_),
    .B1(_11142_),
    .B2(_22673_),
    .C1(_11121_),
    .C2(_22608_),
    .ZN(_23919_));
 AOI221_X4 _55124_ (.A(_23919_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [648]),
    .B2(_23107_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [403]),
    .C2(_23610_),
    .ZN(_23920_));
 NAND3_X1 _55125_ (.A1(_23434_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [256]),
    .A3(_23709_),
    .ZN(_23921_));
 AOI22_X1 _55126_ (.A1(_23615_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [354]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [305]),
    .B2(_22903_),
    .ZN(_23922_));
 NAND3_X1 _55127_ (.A1(_10868_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [60]),
    .A3(_23246_),
    .ZN(_23923_));
 NAND3_X1 _55128_ (.A1(_23242_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [207]),
    .A3(_23246_),
    .ZN(_23924_));
 AND4_X1 _55129_ (.A1(_23921_),
    .A2(_23922_),
    .A3(_23923_),
    .A4(_23924_),
    .ZN(_23925_));
 AND3_X1 _55130_ (.A1(_23509_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [158]),
    .A3(_11174_),
    .ZN(_23926_));
 AOI221_X4 _55131_ (.A(_23926_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [109]),
    .B2(_23453_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [11]),
    .C2(_23164_),
    .ZN(_23927_));
 AND3_X1 _55132_ (.A1(_23806_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [452]),
    .A3(_23161_),
    .ZN(_23928_));
 AOI221_X4 _55133_ (.A(_23928_),
    .B1(_23689_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [501]),
    .C1(_23622_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [550]),
    .ZN(_23929_));
 AND4_X4 _55134_ (.A1(_23920_),
    .A2(_23925_),
    .A3(_23927_),
    .A4(_23929_),
    .ZN(_23930_));
 BUF_X4 _55135_ (.A(_22980_),
    .Z(_23931_));
 NAND3_X1 _55136_ (.A1(_23434_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1432]),
    .A3(_23931_),
    .ZN(_23932_));
 AOI22_X4 _55137_ (.A1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1383]),
    .A2(_23094_),
    .B1(_23103_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1187]),
    .ZN(_23933_));
 NAND3_X1 _55138_ (.A1(_10804_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1530]),
    .A3(_23693_),
    .ZN(_23934_));
 BUF_X32 _55139_ (.A(_10817_),
    .Z(_23935_));
 NAND3_X1 _55140_ (.A1(_23935_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1481]),
    .A3(_23693_),
    .ZN(_23936_));
 AND4_X4 _55141_ (.A1(_23932_),
    .A2(_23933_),
    .A3(_23934_),
    .A4(_23936_),
    .ZN(_23937_));
 BUF_X8 _55142_ (.A(_11089_),
    .Z(_23938_));
 NAND3_X1 _55143_ (.A1(_10798_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1138]),
    .A3(_23938_),
    .ZN(_23939_));
 OAI221_X2 _55144_ (.A(_23939_),
    .B1(_11086_),
    .B2(_22421_),
    .C1(_11095_),
    .C2(_22467_),
    .ZN(_23940_));
 AOI221_X2 _55145_ (.A(_23940_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1040]),
    .B2(_22435_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [795]),
    .C2(_23267_),
    .ZN(_23941_));
 AND3_X1 _55146_ (.A1(_23173_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [893]),
    .A3(_23804_),
    .ZN(_23942_));
 AOI221_X4 _55147_ (.A(_23942_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [844]),
    .B2(_11110_),
    .C1(_23047_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [942]),
    .ZN(_23943_));
 AND3_X1 _55148_ (.A1(_22521_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1285]),
    .A3(_23701_),
    .ZN(_23944_));
 AOI221_X2 _55149_ (.A(_23944_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1236]),
    .B2(_11065_),
    .C1(_23748_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1334]),
    .ZN(_23945_));
 AND4_X4 _55150_ (.A1(_23937_),
    .A2(_23941_),
    .A3(_23943_),
    .A4(_23945_),
    .ZN(_23946_));
 AND3_X1 _55151_ (.A1(_23509_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2118]),
    .A3(_23657_),
    .ZN(_23947_));
 AOI221_X4 _55152_ (.A(_23947_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2069]),
    .B2(_22910_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2020]),
    .C2(_23156_),
    .ZN(_23948_));
 NAND3_X1 _55153_ (.A1(_10798_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2314]),
    .A3(_10939_),
    .ZN(_23949_));
 OAI221_X2 _55154_ (.A(_23949_),
    .B1(_21851_),
    .B2(_10951_),
    .C1(_10946_),
    .C2(_21832_),
    .ZN(_23950_));
 AOI221_X2 _55155_ (.A(_23950_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2167]),
    .B2(_10955_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1971]),
    .C2(_10976_),
    .ZN(_23951_));
 AND3_X1 _55156_ (.A1(_23309_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2559]),
    .A3(_23669_),
    .ZN(_23952_));
 AOI221_X4 _55157_ (.A(_23952_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2657]),
    .B2(_21601_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2706]),
    .C2(_23373_),
    .ZN(_23953_));
 AOI22_X2 _55158_ (.A1(_10929_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2363]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2608]),
    .B2(_23627_),
    .ZN(_23954_));
 AND4_X4 _55159_ (.A1(_23948_),
    .A2(_23951_),
    .A3(_23953_),
    .A4(_23954_),
    .ZN(_23955_));
 AND3_X1 _55160_ (.A1(_23751_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1873]),
    .A3(_22923_),
    .ZN(_23956_));
 AOI221_X4 _55161_ (.A(_23956_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1824]),
    .B2(_23286_),
    .C1(_23584_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1922]),
    .ZN(_23957_));
 OAI22_X2 _55162_ (.A1(_11026_),
    .A2(_22165_),
    .B1(_22138_),
    .B2(_11020_),
    .ZN(_23958_));
 OAI22_X2 _55163_ (.A1(_11009_),
    .A2(_22087_),
    .B1(_22119_),
    .B2(_11013_),
    .ZN(_23959_));
 AOI211_X2 _55164_ (.A(_23958_),
    .B(_23959_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1775]),
    .C2(_11003_),
    .ZN(_23960_));
 NAND3_X1 _55165_ (.A1(_23245_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3098]),
    .A3(_23360_),
    .ZN(_23961_));
 NAND3_X1 _55166_ (.A1(_23240_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3049]),
    .A3(_22990_),
    .ZN(_23962_));
 NAND2_X2 _55167_ (.A1(_23961_),
    .A2(_23962_),
    .ZN(_23963_));
 AND3_X1 _55168_ (.A1(_22932_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2951]),
    .A3(_23122_),
    .ZN(_23964_));
 AND3_X1 _55169_ (.A1(_23303_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3000]),
    .A3(_23122_),
    .ZN(_23965_));
 NOR3_X4 _55170_ (.A1(_23963_),
    .A2(_23964_),
    .A3(_23965_),
    .ZN(_23966_));
 OAI22_X1 _55171_ (.A1(_10913_),
    .A2(_21691_),
    .B1(_21719_),
    .B2(_10917_),
    .ZN(_23967_));
 NAND3_X1 _55172_ (.A1(_22954_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2902]),
    .A3(_22928_),
    .ZN(_23968_));
 OAI21_X2 _55173_ (.A(_23968_),
    .B1(_10852_),
    .B2(_21509_),
    .ZN(_23969_));
 NAND3_X2 _55174_ (.A1(_23084_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2755]),
    .A3(_22928_),
    .ZN(_23970_));
 OAI21_X4 _55175_ (.A(_23970_),
    .B1(_10864_),
    .B2(_21543_),
    .ZN(_23971_));
 AND3_X1 _55176_ (.A1(_23041_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2412]),
    .A3(_10891_),
    .ZN(_23972_));
 NOR4_X1 _55177_ (.A1(_23967_),
    .A2(_23969_),
    .A3(_23971_),
    .A4(_23972_),
    .ZN(_23973_));
 AND4_X1 _55178_ (.A1(_23957_),
    .A2(net15),
    .A3(_23966_),
    .A4(_23973_),
    .ZN(_23974_));
 NAND4_X2 _55179_ (.A1(_23930_),
    .A2(_23946_),
    .A3(_23955_),
    .A4(_23974_),
    .ZN(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [11]));
 AND3_X1 _55180_ (.A1(_22920_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [306]),
    .A3(_23643_),
    .ZN(_23975_));
 AOI221_X4 _55181_ (.A(_23975_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [257]),
    .B2(_22777_),
    .C1(_23615_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [355]),
    .ZN(_23976_));
 NAND3_X1 _55182_ (.A1(_23207_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [796]),
    .A3(_23317_),
    .ZN(_23977_));
 AOI22_X4 _55183_ (.A1(_23047_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [943]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [894]),
    .B2(_23265_),
    .ZN(_23978_));
 NAND3_X1 _55184_ (.A1(_10868_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [845]),
    .A3(_23321_),
    .ZN(_23979_));
 NAND3_X1 _55185_ (.A1(_22241_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1041]),
    .A3(_23321_),
    .ZN(_23980_));
 AND4_X4 _55186_ (.A1(_23977_),
    .A2(_23978_),
    .A3(_23979_),
    .A4(_23980_),
    .ZN(_23981_));
 BUF_X32 _55187_ (.A(_22522_),
    .Z(_23982_));
 NAND3_X1 _55188_ (.A1(_23982_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [110]),
    .A3(_23709_),
    .ZN(_23983_));
 AOI22_X4 _55189_ (.A1(_11206_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [12]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [61]),
    .B2(_23714_),
    .ZN(_23984_));
 NAND3_X1 _55190_ (.A1(_23242_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [208]),
    .A3(_23451_),
    .ZN(_23985_));
 NAND3_X1 _55191_ (.A1(_23003_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [159]),
    .A3(_23451_),
    .ZN(_23986_));
 AND4_X4 _55192_ (.A1(_23983_),
    .A2(_23984_),
    .A3(_23985_),
    .A4(_23986_),
    .ZN(_23987_));
 AND3_X1 _55193_ (.A1(_23487_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1139]),
    .A3(_23804_),
    .ZN(_23988_));
 AOI221_X2 _55194_ (.A(_23988_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1090]),
    .B2(_22410_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [992]),
    .C2(_23104_),
    .ZN(_23989_));
 AND4_X4 _55195_ (.A1(_23976_),
    .A2(_23981_),
    .A3(_23987_),
    .A4(net52),
    .ZN(_23990_));
 AND3_X4 _55196_ (.A1(_23492_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1923]),
    .A3(_22921_),
    .ZN(_23991_));
 AOI221_X2 _55197_ (.A(_23991_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1874]),
    .B2(_22003_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1825]),
    .C2(_23286_),
    .ZN(_23992_));
 NAND3_X1 _55198_ (.A1(_22993_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1580]),
    .A3(_23576_),
    .ZN(_23993_));
 AOI22_X4 _55199_ (.A1(_23467_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1727]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1678]),
    .B2(_22105_),
    .ZN(_23994_));
 NAND3_X1 _55200_ (.A1(_23367_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1776]),
    .A3(_10989_),
    .ZN(_23995_));
 NAND3_X1 _55201_ (.A1(_23293_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1629]),
    .A3(_10989_),
    .ZN(_23996_));
 AND4_X4 _55202_ (.A1(_23993_),
    .A2(_23994_),
    .A3(_23995_),
    .A4(_23996_),
    .ZN(_23997_));
 AND3_X1 _55203_ (.A1(_23810_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2707]),
    .A3(_23669_),
    .ZN(_23998_));
 AOI221_X2 _55204_ (.A(_23998_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2658]),
    .B2(_21601_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2560]),
    .C2(_21654_),
    .ZN(_23999_));
 NAND3_X1 _55205_ (.A1(_22241_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2609]),
    .A3(_10892_),
    .ZN(_24000_));
 AOI22_X2 _55206_ (.A1(_23300_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2364]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2413]),
    .B2(_23301_),
    .ZN(_24001_));
 NAND3_X1 _55207_ (.A1(_23306_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2462]),
    .A3(_23119_),
    .ZN(_24002_));
 NAND3_X1 _55208_ (.A1(_23019_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2511]),
    .A3(_23304_),
    .ZN(_24003_));
 AND4_X4 _55209_ (.A1(_24000_),
    .A2(_24001_),
    .A3(_24002_),
    .A4(_24003_),
    .ZN(_24004_));
 AND4_X4 _55210_ (.A1(_23992_),
    .A2(_23997_),
    .A3(_23999_),
    .A4(_24004_),
    .ZN(_24005_));
 AND3_X1 _55211_ (.A1(_23775_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2805]),
    .A3(_23498_),
    .ZN(_24006_));
 AOI221_X4 _55212_ (.A(_24006_),
    .B1(_10851_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2854]),
    .C1(_21466_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2903]),
    .ZN(_24007_));
 AOI22_X2 _55213_ (.A1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2756]),
    .A2(_23625_),
    .B1(_10839_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2952]),
    .ZN(_24008_));
 AOI22_X1 _55214_ (.A1(_23224_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3099]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3050]),
    .B2(_23225_),
    .ZN(_24009_));
 NAND3_X1 _55215_ (.A1(_23385_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3001]),
    .A3(_23222_),
    .ZN(_24010_));
 AND3_X4 _55216_ (.A1(_24008_),
    .A2(_24009_),
    .A3(_24010_),
    .ZN(_24011_));
 NAND3_X1 _55217_ (.A1(_23935_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2266]),
    .A3(_23553_),
    .ZN(_24012_));
 AOI22_X2 _55218_ (.A1(_23660_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2168]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2021]),
    .B2(_21937_),
    .ZN(_24013_));
 NAND3_X1 _55219_ (.A1(_23757_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2217]),
    .A3(_23388_),
    .ZN(_24014_));
 NAND3_X1 _55220_ (.A1(_22949_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2315]),
    .A3(_23005_),
    .ZN(_24015_));
 AND4_X4 _55221_ (.A1(_24012_),
    .A2(_24013_),
    .A3(_24014_),
    .A4(_24015_),
    .ZN(_24016_));
 AND3_X1 _55222_ (.A1(_23083_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1972]),
    .A3(_23169_),
    .ZN(_24017_));
 AOI221_X4 _55223_ (.A(_24017_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2070]),
    .B2(_10968_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2119]),
    .C2(_23736_),
    .ZN(_24018_));
 AND4_X2 _55224_ (.A1(_24007_),
    .A2(_24011_),
    .A3(_24016_),
    .A4(_24018_),
    .ZN(_24019_));
 AOI22_X4 _55225_ (.A1(_23638_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [747]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [698]),
    .B2(_23092_),
    .ZN(_24020_));
 NAND3_X2 _55226_ (.A1(_22242_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [649]),
    .A3(_22995_),
    .ZN(_24021_));
 NAND3_X2 _55227_ (.A1(_23368_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [600]),
    .A3(_23057_),
    .ZN(_24022_));
 NAND3_X2 _55228_ (.A1(_23377_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [453]),
    .A3(_23057_),
    .ZN(_24023_));
 NAND4_X4 _55229_ (.A1(_24020_),
    .A2(_24021_),
    .A3(_24022_),
    .A4(_24023_),
    .ZN(_24024_));
 AOI22_X4 _55230_ (.A1(_23315_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1531]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1482]),
    .B2(_23095_),
    .ZN(_24025_));
 BUF_X8 _55231_ (.A(_11036_),
    .Z(_24026_));
 NAND3_X2 _55232_ (.A1(_23059_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1384]),
    .A3(_24026_),
    .ZN(_24027_));
 NAND3_X2 _55233_ (.A1(_22968_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1188]),
    .A3(_11037_),
    .ZN(_24028_));
 BUF_X16 _55234_ (.A(_10830_),
    .Z(_24029_));
 NAND3_X2 _55235_ (.A1(_24029_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1433]),
    .A3(_23566_),
    .ZN(_24030_));
 NAND4_X4 _55236_ (.A1(_24025_),
    .A2(_24027_),
    .A3(_24028_),
    .A4(_24030_),
    .ZN(_24031_));
 NAND3_X2 _55237_ (.A1(_23036_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1237]),
    .A3(_23277_),
    .ZN(_24032_));
 NAND3_X2 _55238_ (.A1(_23078_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1286]),
    .A3(_23277_),
    .ZN(_24033_));
 OAI211_X4 _55239_ (.A(_24032_),
    .B(_24033_),
    .C1(_11055_),
    .C2(_22290_),
    .ZN(_24034_));
 NAND3_X2 _55240_ (.A1(_23421_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [551]),
    .A3(_23072_),
    .ZN(_24035_));
 NAND3_X2 _55241_ (.A1(_23085_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [404]),
    .A3(_23208_),
    .ZN(_24036_));
 OAI211_X4 _55242_ (.A(_24035_),
    .B(_24036_),
    .C1(_11154_),
    .C2(_22707_),
    .ZN(_24037_));
 NOR4_X4 _55243_ (.A1(_24024_),
    .A2(_24031_),
    .A3(_24034_),
    .A4(_24037_),
    .ZN(_24038_));
 NAND4_X1 _55244_ (.A1(_23990_),
    .A2(_24005_),
    .A3(_24019_),
    .A4(net4),
    .ZN(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [12]));
 AND3_X1 _55245_ (.A1(_23168_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3002]),
    .A3(_23174_),
    .ZN(_24039_));
 AOI221_X2 _55246_ (.A(_24039_),
    .B1(_23225_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3051]),
    .C1(_23224_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3100]),
    .ZN(_24040_));
 OAI21_X2 _55247_ (.A(_24040_),
    .B1(_21450_),
    .B2(_10840_),
    .ZN(_24041_));
 AOI22_X4 _55248_ (.A1(_23213_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2904]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2855]),
    .B2(_21502_),
    .ZN(_24042_));
 OAI221_X2 _55249_ (.A(_24042_),
    .B1(_21318_),
    .B2(_10875_),
    .C1(_21548_),
    .C2(_10864_),
    .ZN(_24043_));
 NAND3_X2 _55250_ (.A1(_23008_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1973]),
    .A3(_23561_),
    .ZN(_24044_));
 BUF_X16 _55251_ (.A(_23019_),
    .Z(_24045_));
 BUF_X8 _55252_ (.A(_22963_),
    .Z(_24046_));
 NAND3_X2 _55253_ (.A1(_24045_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2120]),
    .A3(_24046_),
    .ZN(_24047_));
 OAI211_X4 _55254_ (.A(_24044_),
    .B(_24047_),
    .C1(_10969_),
    .C2(_21910_),
    .ZN(_24048_));
 AOI22_X4 _55255_ (.A1(_10956_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2169]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2022]),
    .B2(_22911_),
    .ZN(_24049_));
 BUF_X32 _55256_ (.A(_22943_),
    .Z(_24050_));
 NAND3_X1 _55257_ (.A1(_24050_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2267]),
    .A3(_24046_),
    .ZN(_24051_));
 BUF_X8 _55258_ (.A(_22963_),
    .Z(_24052_));
 NAND3_X2 _55259_ (.A1(_22958_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2218]),
    .A3(_24052_),
    .ZN(_24053_));
 NAND3_X2 _55260_ (.A1(_23076_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2316]),
    .A3(_23894_),
    .ZN(_24054_));
 NAND4_X4 _55261_ (.A1(_24049_),
    .A2(_24051_),
    .A3(_24053_),
    .A4(_24054_),
    .ZN(_24055_));
 NOR4_X2 _55262_ (.A1(_24041_),
    .A2(_24043_),
    .A3(_24048_),
    .A4(_24055_),
    .ZN(_24056_));
 NAND3_X1 _55263_ (.A1(_23434_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1434]),
    .A3(_23931_),
    .ZN(_24057_));
 AOI22_X2 _55264_ (.A1(_23315_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1532]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1483]),
    .B2(_22210_),
    .ZN(_24058_));
 NAND3_X1 _55265_ (.A1(_23339_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1385]),
    .A3(_23693_),
    .ZN(_24059_));
 NAND3_X1 _55266_ (.A1(_22993_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1189]),
    .A3(_23693_),
    .ZN(_24060_));
 AND4_X4 _55267_ (.A1(_24057_),
    .A2(_24058_),
    .A3(_24059_),
    .A4(_24060_),
    .ZN(_24061_));
 NAND3_X1 _55268_ (.A1(_23328_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [993]),
    .A3(_23329_),
    .ZN(_24062_));
 AOI22_X1 _55269_ (.A1(_23331_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1140]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1091]),
    .B2(_22410_),
    .ZN(_24063_));
 NAND3_X1 _55270_ (.A1(_23252_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1042]),
    .A3(_23321_),
    .ZN(_24064_));
 NAND3_X1 _55271_ (.A1(_23293_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [846]),
    .A3(_11081_),
    .ZN(_24065_));
 AND4_X1 _55272_ (.A1(_24062_),
    .A2(_24063_),
    .A3(_24064_),
    .A4(_24065_),
    .ZN(_24066_));
 NAND3_X1 _55273_ (.A1(_10780_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [944]),
    .A3(_23317_),
    .ZN(_24067_));
 NAND3_X1 _55274_ (.A1(_23207_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [797]),
    .A3(_23329_),
    .ZN(_24068_));
 NAND3_X1 _55275_ (.A1(_23982_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [895]),
    .A3(_23329_),
    .ZN(_24069_));
 AND3_X1 _55276_ (.A1(_24067_),
    .A2(_24068_),
    .A3(_24069_),
    .ZN(_24070_));
 AND3_X1 _55277_ (.A1(_23176_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1238]),
    .A3(_23701_),
    .ZN(_24071_));
 AOI221_X4 _55278_ (.A(_24071_),
    .B1(_11060_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1287]),
    .C1(_23748_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1336]),
    .ZN(_24072_));
 AND4_X4 _55279_ (.A1(_24061_),
    .A2(_24066_),
    .A3(_24070_),
    .A4(_24072_),
    .ZN(_24073_));
 AND3_X1 _55280_ (.A1(_23284_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1924]),
    .A3(_22923_),
    .ZN(_24074_));
 AOI221_X2 _55281_ (.A(_24074_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1875]),
    .B2(_22003_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1826]),
    .C2(_23286_),
    .ZN(_24075_));
 NAND3_X1 _55282_ (.A1(_10868_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1630]),
    .A3(_23393_),
    .ZN(_24076_));
 AOI22_X2 _55283_ (.A1(_23467_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1728]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1679]),
    .B2(_22105_),
    .ZN(_24077_));
 NAND3_X1 _55284_ (.A1(_10879_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1581]),
    .A3(_10989_),
    .ZN(_24078_));
 NAND3_X1 _55285_ (.A1(_23296_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1777]),
    .A3(_23294_),
    .ZN(_24079_));
 AND4_X4 _55286_ (.A1(_24076_),
    .A2(_24077_),
    .A3(_24078_),
    .A4(_24079_),
    .ZN(_24080_));
 NAND3_X1 _55287_ (.A1(_23113_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2414]),
    .A3(_10892_),
    .ZN(_24081_));
 AOI22_X4 _55288_ (.A1(_23587_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2512]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2463]),
    .B2(_21705_),
    .ZN(_24082_));
 NAND3_X1 _55289_ (.A1(_23455_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2365]),
    .A3(_23304_),
    .ZN(_24083_));
 NAND3_X1 _55290_ (.A1(_23303_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2610]),
    .A3(_23304_),
    .ZN(_24084_));
 AND4_X2 _55291_ (.A1(_24081_),
    .A2(_24082_),
    .A3(_24083_),
    .A4(_24084_),
    .ZN(_24085_));
 AND3_X1 _55292_ (.A1(_23309_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2561]),
    .A3(_23669_),
    .ZN(_24086_));
 AOI221_X2 _55293_ (.A(_24086_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2659]),
    .B2(_21601_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2708]),
    .C2(_23373_),
    .ZN(_24087_));
 AND4_X4 _55294_ (.A1(net51),
    .A2(_24080_),
    .A3(_24085_),
    .A4(_24087_),
    .ZN(_24088_));
 NAND3_X1 _55295_ (.A1(_23385_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [258]),
    .A3(_23709_),
    .ZN(_24089_));
 AOI22_X1 _55296_ (.A1(_23248_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [209]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [62]),
    .B2(_23714_),
    .ZN(_24090_));
 NAND3_X1 _55297_ (.A1(_23935_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [307]),
    .A3(_23451_),
    .ZN(_24091_));
 NAND3_X1 _55298_ (.A1(_10804_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [356]),
    .A3(_23250_),
    .ZN(_24092_));
 AND4_X1 _55299_ (.A1(_24089_),
    .A2(_24090_),
    .A3(_24091_),
    .A4(_24092_),
    .ZN(_24093_));
 NAND3_X1 _55300_ (.A1(_23230_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [405]),
    .A3(_23161_),
    .ZN(_24094_));
 NAND3_X1 _55301_ (.A1(_23733_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [454]),
    .A3(_23161_),
    .ZN(_24095_));
 NAND2_X1 _55302_ (.A1(_24094_),
    .A2(_24095_),
    .ZN(_24096_));
 AOI221_X4 _55303_ (.A(_24096_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [552]),
    .B2(_11146_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [503]),
    .C2(_23689_),
    .ZN(_24097_));
 NAND3_X1 _55304_ (.A1(_10804_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [748]),
    .A3(_23346_),
    .ZN(_24098_));
 NAND3_X1 _55305_ (.A1(_23296_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [601]),
    .A3(_23346_),
    .ZN(_24099_));
 NAND3_X1 _55306_ (.A1(_23303_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [650]),
    .A3(_23056_),
    .ZN(_24100_));
 NAND3_X1 _55307_ (.A1(_22943_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [699]),
    .A3(_23056_),
    .ZN(_24101_));
 AND4_X4 _55308_ (.A1(_24098_),
    .A2(_24099_),
    .A3(_24100_),
    .A4(_24101_),
    .ZN(_24102_));
 AND3_X1 _55309_ (.A1(_10778_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [160]),
    .A3(_22937_),
    .ZN(_24103_));
 AOI221_X4 _55310_ (.A(_24103_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [111]),
    .B2(_11200_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [13]),
    .C2(_11205_),
    .ZN(_24104_));
 AND4_X4 _55311_ (.A1(_24093_),
    .A2(_24097_),
    .A3(_24102_),
    .A4(_24104_),
    .ZN(_24105_));
 NAND4_X4 _55312_ (.A1(_24056_),
    .A2(_24073_),
    .A3(_24088_),
    .A4(_24105_),
    .ZN(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [13]));
 NAND3_X1 _55313_ (.A1(_23288_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [896]),
    .A3(_11080_),
    .ZN(_24106_));
 NAND3_X4 _55314_ (.A1(_10829_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1827]),
    .A3(_10988_),
    .ZN(_24107_));
 NAND2_X1 _55315_ (.A1(_24106_),
    .A2(_24107_),
    .ZN(_24108_));
 AOI221_X4 _55316_ (.A(_24108_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [504]),
    .B2(_23689_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [994]),
    .C2(_23104_),
    .ZN(_24109_));
 NAND3_X1 _55317_ (.A1(_22897_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1533]),
    .A3(_11035_),
    .ZN(_24110_));
 NAND3_X4 _55318_ (.A1(_23721_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2072]),
    .A3(_22913_),
    .ZN(_24111_));
 NAND2_X2 _55319_ (.A1(_24110_),
    .A2(_24111_),
    .ZN(_24112_));
 AOI221_X2 _55320_ (.A(_24112_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1386]),
    .B2(_23094_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1288]),
    .C2(_23262_),
    .ZN(_24113_));
 NAND3_X1 _55321_ (.A1(_23492_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [749]),
    .A3(_23151_),
    .ZN(_24114_));
 NAND3_X1 _55322_ (.A1(_23153_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [602]),
    .A3(_23510_),
    .ZN(_24115_));
 NAND2_X2 _55323_ (.A1(_24114_),
    .A2(_24115_),
    .ZN(_24116_));
 AOI221_X2 _55324_ (.A(_24116_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1092]),
    .B2(_22410_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1043]),
    .C2(_23632_),
    .ZN(_24117_));
 NAND3_X2 _55325_ (.A1(_23492_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1141]),
    .A3(_23494_),
    .ZN(_24118_));
 NAND3_X2 _55326_ (.A1(_23775_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [455]),
    .A3(_23512_),
    .ZN(_24119_));
 NAND2_X4 _55327_ (.A1(_24118_),
    .A2(_24119_),
    .ZN(_24120_));
 AOI221_X2 _55328_ (.A(_24120_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2954]),
    .B2(_10838_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2170]),
    .C2(_23660_),
    .ZN(_24121_));
 AND4_X4 _55329_ (.A1(_24109_),
    .A2(net14),
    .A3(net35),
    .A4(net34),
    .ZN(_24122_));
 AND3_X1 _55330_ (.A1(_23035_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [847]),
    .A3(_22969_),
    .ZN(_24123_));
 AOI21_X4 _55331_ (.A(_24123_),
    .B1(_23267_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [798]),
    .ZN(_24124_));
 OAI221_X2 _55332_ (.A(_24124_),
    .B1(_22843_),
    .B2(_11201_),
    .C1(_22869_),
    .C2(_11207_),
    .ZN(_24125_));
 BUF_X32 _55333_ (.A(_23390_),
    .Z(_24126_));
 NAND3_X1 _55334_ (.A1(_24126_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1925]),
    .A3(_22935_),
    .ZN(_24127_));
 NAND3_X2 _55335_ (.A1(_23125_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1729]),
    .A3(_22935_),
    .ZN(_24128_));
 NAND3_X2 _55336_ (.A1(_23059_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1778]),
    .A3(_22935_),
    .ZN(_24129_));
 NAND3_X2 _55337_ (.A1(_23127_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1876]),
    .A3(_23009_),
    .ZN(_24130_));
 NAND4_X4 _55338_ (.A1(_24127_),
    .A2(_24128_),
    .A3(_24129_),
    .A4(_24130_),
    .ZN(_24131_));
 NAND3_X4 _55339_ (.A1(_24045_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [161]),
    .A3(_22951_),
    .ZN(_24132_));
 NAND3_X4 _55340_ (.A1(_23076_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2709]),
    .A3(_23134_),
    .ZN(_24133_));
 NAND3_X2 _55341_ (.A1(_23189_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1631]),
    .A3(_23141_),
    .ZN(_24134_));
 NAND3_X4 _55342_ (.A1(_23025_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1680]),
    .A3(_23830_),
    .ZN(_24135_));
 NAND4_X4 _55343_ (.A1(_24132_),
    .A2(_24133_),
    .A3(_24134_),
    .A4(_24135_),
    .ZN(_24136_));
 NAND3_X4 _55344_ (.A1(_23020_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [553]),
    .A3(_23063_),
    .ZN(_24137_));
 NAND3_X2 _55345_ (.A1(_22972_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2660]),
    .A3(_23023_),
    .ZN(_24138_));
 NAND3_X2 _55346_ (.A1(_23276_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2562]),
    .A3(_23143_),
    .ZN(_24139_));
 NAND3_X2 _55347_ (.A1(_22978_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2611]),
    .A3(_23029_),
    .ZN(_24140_));
 NAND4_X4 _55348_ (.A1(_24137_),
    .A2(_24138_),
    .A3(_24139_),
    .A4(_24140_),
    .ZN(_24141_));
 NOR4_X1 _55349_ (.A1(_24125_),
    .A2(_24131_),
    .A3(_24136_),
    .A4(_24141_),
    .ZN(_24142_));
 NAND3_X4 _55350_ (.A1(_22985_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2121]),
    .A3(_10942_),
    .ZN(_24143_));
 NAND3_X4 _55351_ (.A1(_24126_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3101]),
    .A3(_22991_),
    .ZN(_24144_));
 NAND3_X4 _55352_ (.A1(_22994_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1974]),
    .A3(_23554_),
    .ZN(_24145_));
 NAND3_X4 _55353_ (.A1(_22998_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3003]),
    .A3(_23000_),
    .ZN(_24146_));
 NAND4_X4 _55354_ (.A1(_24143_),
    .A2(_24144_),
    .A3(_24145_),
    .A4(_24146_),
    .ZN(_24147_));
 NAND3_X2 _55355_ (.A1(_24126_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2317]),
    .A3(_23006_),
    .ZN(_24148_));
 NAND3_X4 _55356_ (.A1(_22944_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [308]),
    .A3(_22951_),
    .ZN(_24149_));
 NAND3_X2 _55357_ (.A1(_23536_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2219]),
    .A3(_24046_),
    .ZN(_24150_));
 NAND3_X2 _55358_ (.A1(_24050_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2268]),
    .A3(_24052_),
    .ZN(_24151_));
 NAND4_X4 _55359_ (.A1(_24148_),
    .A2(_24149_),
    .A3(_24150_),
    .A4(_24151_),
    .ZN(_24152_));
 NAND3_X2 _55360_ (.A1(_22968_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2758]),
    .A3(_23128_),
    .ZN(_24153_));
 NAND3_X2 _55361_ (.A1(_22972_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3052]),
    .A3(_10790_),
    .ZN(_24154_));
 NAND3_X4 _55362_ (.A1(_22961_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1484]),
    .A3(_23277_),
    .ZN(_24155_));
 NAND3_X4 _55363_ (.A1(_23071_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1435]),
    .A3(_22981_),
    .ZN(_24156_));
 NAND4_X2 _55364_ (.A1(_24153_),
    .A2(_24154_),
    .A3(_24155_),
    .A4(_24156_),
    .ZN(_24157_));
 NAND3_X1 _55365_ (.A1(_23140_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2464]),
    .A3(_23134_),
    .ZN(_24158_));
 NAND3_X4 _55366_ (.A1(_23036_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [63]),
    .A3(_22959_),
    .ZN(_24159_));
 NAND3_X4 _55367_ (.A1(_23145_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1239]),
    .A3(_23205_),
    .ZN(_24160_));
 NAND3_X2 _55368_ (.A1(_23426_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2415]),
    .A3(_23043_),
    .ZN(_24161_));
 NAND4_X4 _55369_ (.A1(_24158_),
    .A2(_24159_),
    .A3(_24160_),
    .A4(_24161_),
    .ZN(_24162_));
 NOR4_X4 _55370_ (.A1(_24147_),
    .A2(_24152_),
    .A3(_24157_),
    .A4(_24162_),
    .ZN(_24163_));
 NAND3_X2 _55371_ (.A1(_22524_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2856]),
    .A3(_23000_),
    .ZN(_24164_));
 AOI22_X4 _55372_ (.A1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2807]),
    .A2(_21536_),
    .B1(_22911_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2023]),
    .ZN(_24165_));
 OAI211_X4 _55373_ (.A(_24164_),
    .B(_24165_),
    .C1(_10774_),
    .C2(_21475_),
    .ZN(_24166_));
 NAND3_X4 _55374_ (.A1(_23054_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [357]),
    .A3(_22940_),
    .ZN(_24167_));
 NAND3_X4 _55375_ (.A1(_24045_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1337]),
    .A3(_24026_),
    .ZN(_24168_));
 NAND3_X2 _55376_ (.A1(_23020_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2513]),
    .A3(_23014_),
    .ZN(_24169_));
 NAND3_X4 _55377_ (.A1(_23133_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1582]),
    .A3(_22956_),
    .ZN(_24170_));
 NAND4_X4 _55378_ (.A1(_24167_),
    .A2(_24168_),
    .A3(_24169_),
    .A4(_24170_),
    .ZN(_24171_));
 NAND3_X1 _55379_ (.A1(_23192_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [210]),
    .A3(_23187_),
    .ZN(_24172_));
 NAND3_X4 _55380_ (.A1(_23194_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1190]),
    .A3(_23274_),
    .ZN(_24173_));
 NAND3_X2 _55381_ (.A1(_23837_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2366]),
    .A3(_23143_),
    .ZN(_24174_));
 NAND3_X1 _55382_ (.A1(_22978_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [259]),
    .A3(_23086_),
    .ZN(_24175_));
 NAND4_X1 _55383_ (.A1(_24172_),
    .A2(_24173_),
    .A3(_24174_),
    .A4(_24175_),
    .ZN(_24176_));
 NAND3_X2 _55384_ (.A1(_23200_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [945]),
    .A3(_22973_),
    .ZN(_24177_));
 NAND3_X2 _55385_ (.A1(_23071_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [651]),
    .A3(_23072_),
    .ZN(_24178_));
 NAND3_X2 _55386_ (.A1(_23280_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [700]),
    .A3(_23208_),
    .ZN(_24179_));
 NAND3_X2 _55387_ (.A1(_23207_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [406]),
    .A3(_23208_),
    .ZN(_24180_));
 NAND4_X4 _55388_ (.A1(_24177_),
    .A2(_24178_),
    .A3(_24179_),
    .A4(_24180_),
    .ZN(_24181_));
 NOR4_X1 _55389_ (.A1(_24166_),
    .A2(_24171_),
    .A3(_24176_),
    .A4(_24181_),
    .ZN(_24182_));
 NAND4_X1 _55390_ (.A1(_24122_),
    .A2(_24142_),
    .A3(_24163_),
    .A4(_24182_),
    .ZN(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [14]));
 NAND3_X1 _55391_ (.A1(_23236_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [358]),
    .A3(_23709_),
    .ZN(_24183_));
 AOI22_X2 _55392_ (.A1(_23248_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [211]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [64]),
    .B2(_23714_),
    .ZN(_24184_));
 NAND3_X1 _55393_ (.A1(_23434_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [260]),
    .A3(_23709_),
    .ZN(_24185_));
 BUF_X32 _55394_ (.A(_10817_),
    .Z(_24186_));
 NAND3_X1 _55395_ (.A1(_24186_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [309]),
    .A3(_23709_),
    .ZN(_24187_));
 AND4_X1 _55396_ (.A1(_24183_),
    .A2(_24184_),
    .A3(_24185_),
    .A4(_24187_),
    .ZN(_24188_));
 NAND3_X1 _55397_ (.A1(_23806_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [456]),
    .A3(_23161_),
    .ZN(_24189_));
 OAI21_X1 _55398_ (.A(_24189_),
    .B1(_11165_),
    .B2(_22740_),
    .ZN(_24190_));
 AOI221_X2 _55399_ (.A(_24190_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [554]),
    .B2(_11147_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [505]),
    .C2(_11153_),
    .ZN(_24191_));
 NAND3_X1 _55400_ (.A1(_23492_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [750]),
    .A3(_23151_),
    .ZN(_24192_));
 NAND3_X1 _55401_ (.A1(_22942_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [701]),
    .A3(_23510_),
    .ZN(_24193_));
 NAND2_X1 _55402_ (.A1(_24192_),
    .A2(_24193_),
    .ZN(_24194_));
 AOI221_X2 _55403_ (.A(_24194_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [652]),
    .B2(_22642_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [603]),
    .C2(_23515_),
    .ZN(_24195_));
 AND3_X2 _55404_ (.A1(_23158_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [162]),
    .A3(_23159_),
    .ZN(_24196_));
 AOI221_X4 _55405_ (.A(_24196_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [113]),
    .B2(_23453_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [15]),
    .C2(_23164_),
    .ZN(_24197_));
 AND4_X4 _55406_ (.A1(_24188_),
    .A2(_24191_),
    .A3(net33),
    .A4(_24197_),
    .ZN(_24198_));
 AND3_X1 _55407_ (.A1(_23217_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1142]),
    .A3(_23938_),
    .ZN(_24199_));
 AOI221_X2 _55408_ (.A(_24199_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1093]),
    .B2(_23332_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1044]),
    .C2(_22435_),
    .ZN(_24200_));
 AOI22_X2 _55409_ (.A1(_22459_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [995]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [848]),
    .B2(_23268_),
    .ZN(_24201_));
 AND3_X1 _55410_ (.A1(_10877_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [799]),
    .A3(_23938_),
    .ZN(_24202_));
 AOI221_X4 _55411_ (.A(_24202_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [897]),
    .B2(_11106_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [946]),
    .C2(_11100_),
    .ZN(_24203_));
 AND3_X1 _55412_ (.A1(_10866_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1240]),
    .A3(_22979_),
    .ZN(_24204_));
 AOI221_X2 _55413_ (.A(_24204_),
    .B1(_11059_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1289]),
    .C1(_23748_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1338]),
    .ZN(_24205_));
 NAND4_X4 _55414_ (.A1(_24200_),
    .A2(_24201_),
    .A3(_24203_),
    .A4(_24205_),
    .ZN(_24206_));
 AND3_X4 _55415_ (.A1(_10877_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2367]),
    .A3(_10890_),
    .ZN(_24207_));
 AOI221_X2 _55416_ (.A(_24207_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2465]),
    .B2(_10916_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2514]),
    .C2(_10912_),
    .ZN(_24208_));
 AND3_X1 _55417_ (.A1(_10824_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2612]),
    .A3(_10890_),
    .ZN(_24209_));
 AOI221_X4 _55418_ (.A(_24209_),
    .B1(_21600_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2661]),
    .C1(_21573_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2710]),
    .ZN(_24210_));
 AND3_X1 _55419_ (.A1(_10866_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2808]),
    .A3(_10787_),
    .ZN(_24211_));
 AOI221_X2 _55420_ (.A(_24211_),
    .B1(_10851_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2857]),
    .C1(_21466_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2906]),
    .ZN(_24212_));
 AOI22_X4 _55421_ (.A1(_21654_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2563]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2416]),
    .B2(_10922_),
    .ZN(_24213_));
 NAND4_X4 _55422_ (.A1(_24208_),
    .A2(_24210_),
    .A3(_24212_),
    .A4(_24213_),
    .ZN(_24214_));
 AOI22_X4 _55423_ (.A1(_10800_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3102]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3053]),
    .B2(_10813_),
    .ZN(_24215_));
 NAND3_X2 _55424_ (.A1(_22958_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3004]),
    .A3(_23033_),
    .ZN(_24216_));
 NAND3_X2 _55425_ (.A1(_23022_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2759]),
    .A3(_10790_),
    .ZN(_24217_));
 NAND3_X1 _55426_ (.A1(_23276_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2955]),
    .A3(_10790_),
    .ZN(_24218_));
 NAND4_X4 _55427_ (.A1(_24215_),
    .A2(_24216_),
    .A3(_24217_),
    .A4(_24218_),
    .ZN(_24219_));
 AOI22_X4 _55428_ (.A1(_23315_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1534]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1485]),
    .B2(_23095_),
    .ZN(_24220_));
 NAND3_X1 _55429_ (.A1(_23022_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1191]),
    .A3(_23274_),
    .ZN(_24221_));
 NAND3_X2 _55430_ (.A1(_22975_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1436]),
    .A3(_23277_),
    .ZN(_24222_));
 NAND3_X2 _55431_ (.A1(_23839_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1387]),
    .A3(_22981_),
    .ZN(_24223_));
 NAND4_X4 _55432_ (.A1(_24220_),
    .A2(_24221_),
    .A3(_24222_),
    .A4(_24223_),
    .ZN(_24224_));
 NOR4_X1 _55433_ (.A1(_24206_),
    .A2(_24214_),
    .A3(_24219_),
    .A4(_24224_),
    .ZN(_24225_));
 AND3_X1 _55434_ (.A1(_23487_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1926]),
    .A3(_23519_),
    .ZN(_24226_));
 AND3_X1 _55435_ (.A1(_23215_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1828]),
    .A3(_23402_),
    .ZN(_24227_));
 AND3_X1 _55436_ (.A1(_10816_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1877]),
    .A3(_10987_),
    .ZN(_24228_));
 OR3_X2 _55437_ (.A1(_24226_),
    .A2(_24227_),
    .A3(_24228_),
    .ZN(_24229_));
 AOI221_X2 _55438_ (.A(_24229_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1779]),
    .B2(_11003_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1632]),
    .C2(_23604_),
    .ZN(_24230_));
 NAND3_X2 _55439_ (.A1(_22985_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2122]),
    .A3(_10942_),
    .ZN(_24231_));
 OAI21_X4 _55440_ (.A(_24231_),
    .B1(_10969_),
    .B2(_21912_),
    .ZN(_24232_));
 NAND3_X1 _55441_ (.A1(_23054_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2318]),
    .A3(_23006_),
    .ZN(_24233_));
 NAND3_X2 _55442_ (.A1(_23127_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2269]),
    .A3(_23561_),
    .ZN(_24234_));
 NAND3_X2 _55443_ (.A1(_23011_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2171]),
    .A3(_24046_),
    .ZN(_24235_));
 NAND3_X2 _55444_ (.A1(_24029_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2220]),
    .A3(_24052_),
    .ZN(_24236_));
 NAND4_X4 _55445_ (.A1(_24233_),
    .A2(_24234_),
    .A3(_24235_),
    .A4(_24236_),
    .ZN(_24237_));
 NAND3_X2 _55446_ (.A1(_23125_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1730]),
    .A3(_22935_),
    .ZN(_24238_));
 NAND3_X2 _55447_ (.A1(_23008_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1583]),
    .A3(_23009_),
    .ZN(_24239_));
 NAND3_X2 _55448_ (.A1(_23016_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1681]),
    .A3(_22956_),
    .ZN(_24240_));
 NAND3_X4 _55449_ (.A1(_24238_),
    .A2(_24239_),
    .A3(_24240_),
    .ZN(_24241_));
 NAND3_X1 _55450_ (.A1(_23133_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1975]),
    .A3(_24052_),
    .ZN(_24242_));
 OAI21_X2 _55451_ (.A(_24242_),
    .B1(_10973_),
    .B2(_21947_),
    .ZN(_24243_));
 NOR4_X4 _55452_ (.A1(_24232_),
    .A2(_24237_),
    .A3(_24241_),
    .A4(_24243_),
    .ZN(_24244_));
 NAND4_X1 _55453_ (.A1(_24198_),
    .A2(_24225_),
    .A3(net32),
    .A4(_24244_),
    .ZN(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [15]));
 NAND3_X1 _55454_ (.A1(_23438_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [653]),
    .A3(_23237_),
    .ZN(_24245_));
 AND3_X1 _55455_ (.A1(_22896_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [751]),
    .A3(_11145_),
    .ZN(_24246_));
 AOI221_X2 _55456_ (.A(_24246_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [702]),
    .B2(_11131_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [604]),
    .C2(_11141_),
    .ZN(_24247_));
 AND3_X1 _55457_ (.A1(_10873_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [16]),
    .A3(_11173_),
    .ZN(_24248_));
 AOI221_X2 _55458_ (.A(_24248_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [114]),
    .B2(_11200_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [163]),
    .C2(_11195_),
    .ZN(_24249_));
 NAND3_X1 _55459_ (.A1(_10779_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [555]),
    .A3(_23055_),
    .ZN(_24250_));
 NAND3_X1 _55460_ (.A1(_23288_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [506]),
    .A3(_23055_),
    .ZN(_24251_));
 NAND3_X1 _55461_ (.A1(_10878_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [408]),
    .A3(_23055_),
    .ZN(_24252_));
 NAND3_X2 _55462_ (.A1(_10867_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [457]),
    .A3(_23055_),
    .ZN(_24253_));
 AND4_X1 _55463_ (.A1(_24250_),
    .A2(_24251_),
    .A3(_24252_),
    .A4(_24253_),
    .ZN(_24254_));
 AND4_X4 _55464_ (.A1(_24245_),
    .A2(_24247_),
    .A3(net59),
    .A4(_24254_),
    .ZN(_24255_));
 NAND3_X2 _55465_ (.A1(_22967_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [800]),
    .A3(_23879_),
    .ZN(_24256_));
 OAI221_X2 _55466_ (.A(_24256_),
    .B1(_11107_),
    .B2(_22531_),
    .C1(_11101_),
    .C2(_22507_),
    .ZN(_24257_));
 AND3_X1 _55467_ (.A1(_23019_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1339]),
    .A3(_23608_),
    .ZN(_24258_));
 AND3_X1 _55468_ (.A1(_10857_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1290]),
    .A3(_11036_),
    .ZN(_24259_));
 OAI22_X2 _55469_ (.A1(_11070_),
    .A2(_22373_),
    .B1(_22342_),
    .B2(_11066_),
    .ZN(_24260_));
 NOR4_X1 _55470_ (.A1(_24257_),
    .A2(_24258_),
    .A3(_24259_),
    .A4(_24260_),
    .ZN(_24261_));
 BUF_X32 _55471_ (.A(_10803_),
    .Z(_24262_));
 NAND3_X1 _55472_ (.A1(_24262_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1535]),
    .A3(_23412_),
    .ZN(_24263_));
 NAND3_X1 _55473_ (.A1(_23242_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1388]),
    .A3(_23693_),
    .ZN(_24264_));
 NAND3_X1 _55474_ (.A1(_22997_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1437]),
    .A3(_23050_),
    .ZN(_24265_));
 NAND3_X1 _55475_ (.A1(_23935_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1486]),
    .A3(_23050_),
    .ZN(_24266_));
 AND4_X2 _55476_ (.A1(_24263_),
    .A2(_24264_),
    .A3(_24265_),
    .A4(_24266_),
    .ZN(_24267_));
 NAND3_X4 _55477_ (.A1(_22949_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1143]),
    .A3(_22969_),
    .ZN(_24268_));
 OAI221_X2 _55478_ (.A(_24268_),
    .B1(_22447_),
    .B2(_11091_),
    .C1(_11086_),
    .C2(_22424_),
    .ZN(_24269_));
 NAND3_X1 _55479_ (.A1(_10803_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [359]),
    .A3(_22938_),
    .ZN(_24270_));
 OAI221_X2 _55480_ (.A(_24270_),
    .B1(_22783_),
    .B2(_11187_),
    .C1(_11182_),
    .C2(_22767_),
    .ZN(_24271_));
 OAI22_X2 _55481_ (.A1(_11096_),
    .A2(_22469_),
    .B1(_22559_),
    .B2(_11111_),
    .ZN(_24272_));
 NAND3_X1 _55482_ (.A1(_10843_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [212]),
    .A3(_11175_),
    .ZN(_24273_));
 NAND3_X2 _55483_ (.A1(_23035_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [65]),
    .A3(_11175_),
    .ZN(_24274_));
 NAND2_X4 _55484_ (.A1(_24273_),
    .A2(_24274_),
    .ZN(_24275_));
 NOR4_X4 _55485_ (.A1(_24269_),
    .A2(net31),
    .A3(_24272_),
    .A4(_24275_),
    .ZN(_24276_));
 AND4_X4 _55486_ (.A1(_24255_),
    .A2(_24261_),
    .A3(_24267_),
    .A4(_24276_),
    .ZN(_24277_));
 NAND3_X2 _55487_ (.A1(_22953_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2907]),
    .A3(_10788_),
    .ZN(_24278_));
 OAI21_X1 _55488_ (.A(_24278_),
    .B1(_10852_),
    .B2(_21515_),
    .ZN(_24279_));
 AOI221_X4 _55489_ (.A(_24279_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2760]),
    .B2(_21289_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2809]),
    .C2(_21536_),
    .ZN(_24280_));
 NAND3_X1 _55490_ (.A1(_10845_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2956]),
    .A3(_10791_),
    .ZN(_24281_));
 AND3_X1 _55491_ (.A1(_10829_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3005]),
    .A3(_10788_),
    .ZN(_24282_));
 AOI221_X2 _55492_ (.A(_24282_),
    .B1(_23225_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3054]),
    .C1(_23224_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3103]),
    .ZN(_24283_));
 AND3_X4 _55493_ (.A1(_24280_),
    .A2(_24281_),
    .A3(_24283_),
    .ZN(_24284_));
 NAND3_X1 _55494_ (.A1(_23340_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2564]),
    .A3(_10893_),
    .ZN(_24285_));
 AND3_X1 _55495_ (.A1(_23168_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2613]),
    .A3(_23669_),
    .ZN(_24286_));
 AOI221_X4 _55496_ (.A(_24286_),
    .B1(_23374_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2662]),
    .C1(_23373_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2711]),
    .ZN(_24287_));
 AOI22_X2 _55497_ (.A1(_23587_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2515]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2466]),
    .B2(_21705_),
    .ZN(_24288_));
 AOI22_X2 _55498_ (.A1(_10929_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2368]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2417]),
    .B2(_10922_),
    .ZN(_24289_));
 AND4_X4 _55499_ (.A1(_24285_),
    .A2(_24287_),
    .A3(_24288_),
    .A4(_24289_),
    .ZN(_24290_));
 AND3_X1 _55500_ (.A1(_22521_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1682]),
    .A3(_10987_),
    .ZN(_24291_));
 AOI221_X2 _55501_ (.A(_24291_),
    .B1(_11025_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1584]),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1731]),
    .C2(_22078_),
    .ZN(_24292_));
 NAND3_X1 _55502_ (.A1(_22994_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1976]),
    .A3(_23554_),
    .ZN(_24293_));
 NAND3_X2 _55503_ (.A1(_10858_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2074]),
    .A3(_23554_),
    .ZN(_24294_));
 NAND3_X2 _55504_ (.A1(_23004_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2123]),
    .A3(_23006_),
    .ZN(_24295_));
 NAND4_X4 _55505_ (.A1(net50),
    .A2(_24293_),
    .A3(_24294_),
    .A4(_24295_),
    .ZN(_24296_));
 AOI22_X2 _55506_ (.A1(_10956_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2172]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2025]),
    .B2(_22911_),
    .ZN(_24297_));
 NAND3_X1 _55507_ (.A1(_23127_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2270]),
    .A3(_23561_),
    .ZN(_24298_));
 NAND3_X1 _55508_ (.A1(_23067_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2319]),
    .A3(_24046_),
    .ZN(_24299_));
 NAND3_X2 _55509_ (.A1(_24029_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2221]),
    .A3(_24052_),
    .ZN(_24300_));
 NAND4_X2 _55510_ (.A1(_24297_),
    .A2(_24298_),
    .A3(_24299_),
    .A4(_24300_),
    .ZN(_24301_));
 NAND3_X1 _55511_ (.A1(_23236_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1927]),
    .A3(_23830_),
    .ZN(_24302_));
 NAND3_X1 _55512_ (.A1(_22975_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1829]),
    .A3(_23830_),
    .ZN(_24303_));
 OAI211_X2 _55513_ (.A(_24302_),
    .B(_24303_),
    .C1(_10994_),
    .C2(_22018_),
    .ZN(_24304_));
 OAI22_X4 _55514_ (.A1(_11004_),
    .A2(_22069_),
    .B1(_22144_),
    .B2(_11020_),
    .ZN(_24305_));
 NOR4_X4 _55515_ (.A1(_24296_),
    .A2(_24301_),
    .A3(_24304_),
    .A4(_24305_),
    .ZN(_24306_));
 NAND4_X1 _55516_ (.A1(_24277_),
    .A2(_24284_),
    .A3(_24290_),
    .A4(_24306_),
    .ZN(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [16]));
 AOI22_X4 _55517_ (.A1(_23373_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2712]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2663]),
    .B2(_23374_),
    .ZN(_24307_));
 OAI221_X2 _55518_ (.A(_24307_),
    .B1(_21643_),
    .B2(_10903_),
    .C1(_21664_),
    .C2(_10908_),
    .ZN(_24308_));
 AOI22_X4 _55519_ (.A1(_23587_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2516]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2467]),
    .B2(_21705_),
    .ZN(_24309_));
 OAI221_X2 _55520_ (.A(_24309_),
    .B1(_21754_),
    .B2(_10923_),
    .C1(_21776_),
    .C2(_10930_),
    .ZN(_24310_));
 AOI22_X2 _55521_ (.A1(_23485_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1977]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2026]),
    .B2(_22911_),
    .ZN(_24311_));
 OAI221_X2 _55522_ (.A(_24311_),
    .B1(_21914_),
    .B2(_10969_),
    .C1(_10963_),
    .C2(_21889_),
    .ZN(_24312_));
 NAND3_X2 _55523_ (.A1(_22950_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2320]),
    .A3(_23561_),
    .ZN(_24313_));
 NAND3_X2 _55524_ (.A1(_24050_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2271]),
    .A3(_24046_),
    .ZN(_24314_));
 NAND3_X2 _55525_ (.A1(_23192_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2173]),
    .A3(_23894_),
    .ZN(_24315_));
 NAND3_X2 _55526_ (.A1(_22958_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2222]),
    .A3(_23894_),
    .ZN(_24316_));
 NAND4_X4 _55527_ (.A1(_24313_),
    .A2(_24314_),
    .A3(_24315_),
    .A4(_24316_),
    .ZN(_24317_));
 NOR4_X4 _55528_ (.A1(_24308_),
    .A2(_24310_),
    .A3(_24312_),
    .A4(_24317_),
    .ZN(_24318_));
 AND3_X1 _55529_ (.A1(_23492_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [752]),
    .A3(_23151_),
    .ZN(_24319_));
 AOI221_X2 _55530_ (.A(_24319_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [703]),
    .B2(_11131_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [605]),
    .C2(_23106_),
    .ZN(_24320_));
 NAND3_X1 _55531_ (.A1(_23982_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [507]),
    .A3(_11126_),
    .ZN(_24321_));
 AOI22_X4 _55532_ (.A1(_23610_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [409]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [458]),
    .B2(_11158_),
    .ZN(_24322_));
 NAND3_X1 _55533_ (.A1(_23003_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [556]),
    .A3(_23346_),
    .ZN(_24323_));
 NAND3_X1 _55534_ (.A1(_23252_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [654]),
    .A3(_23346_),
    .ZN(_24324_));
 AND4_X2 _55535_ (.A1(_24321_),
    .A2(_24322_),
    .A3(_24323_),
    .A4(_24324_),
    .ZN(_24325_));
 NAND3_X1 _55536_ (.A1(_23982_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [899]),
    .A3(_23321_),
    .ZN(_24326_));
 AOI22_X1 _55537_ (.A1(_23267_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [801]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [850]),
    .B2(_22544_),
    .ZN(_24327_));
 NAND3_X1 _55538_ (.A1(_23003_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [948]),
    .A3(_11081_),
    .ZN(_24328_));
 NAND3_X1 _55539_ (.A1(_23757_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1046]),
    .A3(_23879_),
    .ZN(_24329_));
 AND4_X1 _55540_ (.A1(_24326_),
    .A2(_24327_),
    .A3(_24328_),
    .A4(_24329_),
    .ZN(_24330_));
 AND3_X1 _55541_ (.A1(_23459_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1144]),
    .A3(_23460_),
    .ZN(_24331_));
 AOI221_X2 _55542_ (.A(_24331_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1095]),
    .B2(_23332_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [997]),
    .C2(_23104_),
    .ZN(_24332_));
 AND4_X4 _55543_ (.A1(_24320_),
    .A2(_24325_),
    .A3(_24330_),
    .A4(_24332_),
    .ZN(_24333_));
 AOI22_X4 _55544_ (.A1(_23290_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1732]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1683]),
    .B2(_23591_),
    .ZN(_24334_));
 AOI22_X4 _55545_ (.A1(_23595_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1585]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1634]),
    .B2(_23604_),
    .ZN(_24335_));
 OAI211_X4 _55546_ (.A(_24334_),
    .B(_24335_),
    .C1(_22071_),
    .C2(_11004_),
    .ZN(_24336_));
 AOI22_X2 _55547_ (.A1(_23213_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2908]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2859]),
    .B2(_21502_),
    .ZN(_24337_));
 AOI22_X2 _55548_ (.A1(_23625_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2761]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2810]),
    .B2(_21536_),
    .ZN(_24338_));
 OAI211_X4 _55549_ (.A(_24337_),
    .B(_24338_),
    .C1(_21454_),
    .C2(_10840_),
    .ZN(_24339_));
 NAND4_X2 _55550_ (.A1(_10751_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3104]),
    .A3(_23033_),
    .A4(_10795_),
    .ZN(_24340_));
 NAND3_X2 _55551_ (.A1(_23536_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3006]),
    .A3(_23128_),
    .ZN(_24341_));
 NAND4_X2 _55552_ (.A1(_10809_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3055]),
    .A3(_10790_),
    .A4(_10795_),
    .ZN(_24342_));
 NAND3_X4 _55553_ (.A1(_24340_),
    .A2(_24341_),
    .A3(_24342_),
    .ZN(_24343_));
 NAND3_X2 _55554_ (.A1(_23560_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1928]),
    .A3(_23009_),
    .ZN(_24344_));
 NAND3_X2 _55555_ (.A1(_23888_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1879]),
    .A3(_22956_),
    .ZN(_24345_));
 NAND3_X2 _55556_ (.A1(_22958_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1830]),
    .A3(_23141_),
    .ZN(_24346_));
 NAND3_X4 _55557_ (.A1(_24344_),
    .A2(_24345_),
    .A3(_24346_),
    .ZN(_24347_));
 NOR4_X1 _55558_ (.A1(_24336_),
    .A2(_24339_),
    .A3(_24343_),
    .A4(_24347_),
    .ZN(_24348_));
 AOI22_X4 _55559_ (.A1(_11206_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [17]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [66]),
    .B2(_23490_),
    .ZN(_24349_));
 OAI221_X2 _55560_ (.A(_24349_),
    .B1(_22847_),
    .B2(_11201_),
    .C1(_11197_),
    .C2(_22819_),
    .ZN(_24350_));
 NAND3_X2 _55561_ (.A1(_23054_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1536]),
    .A3(_22945_),
    .ZN(_24351_));
 NAND3_X2 _55562_ (.A1(_23059_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1389]),
    .A3(_24026_),
    .ZN(_24352_));
 NAND3_X2 _55563_ (.A1(_24050_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1487]),
    .A3(_11037_),
    .ZN(_24353_));
 NAND3_X2 _55564_ (.A1(_24029_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1438]),
    .A3(_23566_),
    .ZN(_24354_));
 NAND4_X4 _55565_ (.A1(_24351_),
    .A2(_24352_),
    .A3(_24353_),
    .A4(_24354_),
    .ZN(_24355_));
 NAND3_X2 _55566_ (.A1(_22955_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1340]),
    .A3(_23566_),
    .ZN(_24356_));
 NAND3_X2 _55567_ (.A1(_23025_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1291]),
    .A3(_23277_),
    .ZN(_24357_));
 NAND3_X1 _55568_ (.A1(_23837_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1193]),
    .A3(_22981_),
    .ZN(_24358_));
 NAND3_X2 _55569_ (.A1(_23145_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1242]),
    .A3(_22981_),
    .ZN(_24359_));
 NAND4_X4 _55570_ (.A1(_24356_),
    .A2(_24357_),
    .A3(_24358_),
    .A4(_24359_),
    .ZN(_24360_));
 NAND3_X1 _55571_ (.A1(_23076_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [360]),
    .A3(_23835_),
    .ZN(_24361_));
 NAND3_X1 _55572_ (.A1(_22978_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [262]),
    .A3(_23196_),
    .ZN(_24362_));
 NAND3_X1 _55573_ (.A1(_23839_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [213]),
    .A3(_23086_),
    .ZN(_24363_));
 NAND3_X1 _55574_ (.A1(_23280_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [311]),
    .A3(_23086_),
    .ZN(_24364_));
 NAND4_X2 _55575_ (.A1(_24361_),
    .A2(_24362_),
    .A3(_24363_),
    .A4(_24364_),
    .ZN(_24365_));
 NOR4_X4 _55576_ (.A1(_24350_),
    .A2(_24355_),
    .A3(_24360_),
    .A4(_24365_),
    .ZN(_24366_));
 NAND4_X1 _55577_ (.A1(_24318_),
    .A2(_24333_),
    .A3(_24348_),
    .A4(_24366_),
    .ZN(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [17]));
 NAND3_X1 _55578_ (.A1(_22897_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3105]),
    .A3(_22989_),
    .ZN(_24367_));
 NAND3_X2 _55579_ (.A1(_10867_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2811]),
    .A3(_22989_),
    .ZN(_24368_));
 NAND2_X1 _55580_ (.A1(_24367_),
    .A2(_24368_),
    .ZN(_24369_));
 AOI221_X2 _55581_ (.A(_24369_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2762]),
    .B2(_21289_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3056]),
    .C2(_10813_),
    .ZN(_24370_));
 NAND3_X2 _55582_ (.A1(_23166_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2909]),
    .A3(_23794_),
    .ZN(_24371_));
 OAI21_X4 _55583_ (.A(_24371_),
    .B1(_10852_),
    .B2(_21518_),
    .ZN(_24372_));
 AOI221_X4 _55584_ (.A(_24372_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2713]),
    .B2(_21573_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2615]),
    .C2(_23627_),
    .ZN(_24373_));
 NAND3_X1 _55585_ (.A1(_23492_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1145]),
    .A3(_22905_),
    .ZN(_24374_));
 NAND3_X2 _55586_ (.A1(_23153_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [998]),
    .A3(_23494_),
    .ZN(_24375_));
 NAND2_X4 _55587_ (.A1(_24374_),
    .A2(_24375_),
    .ZN(_24376_));
 AOI221_X2 _55588_ (.A(_24376_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2076]),
    .B2(_22910_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2027]),
    .C2(_23156_),
    .ZN(_24377_));
 NAND3_X1 _55589_ (.A1(_24186_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1488]),
    .A3(_23412_),
    .ZN(_24378_));
 NAND3_X4 _55590_ (.A1(_22987_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2517]),
    .A3(_10892_),
    .ZN(_24379_));
 NAND3_X1 _55591_ (.A1(_10804_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1537]),
    .A3(_23050_),
    .ZN(_24380_));
 NAND3_X1 _55592_ (.A1(_22523_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1292]),
    .A3(_23050_),
    .ZN(_24381_));
 AND4_X4 _55593_ (.A1(_24378_),
    .A2(_24379_),
    .A3(_24380_),
    .A4(_24381_),
    .ZN(_24382_));
 AND4_X1 _55594_ (.A1(net30),
    .A2(_24373_),
    .A3(_24377_),
    .A4(_24382_),
    .ZN(_24383_));
 AOI22_X4 _55595_ (.A1(_23325_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1194]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1243]),
    .B2(_23048_),
    .ZN(_24384_));
 NAND3_X2 _55596_ (.A1(_22524_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [116]),
    .A3(_23341_),
    .ZN(_24385_));
 OAI211_X4 _55597_ (.A(_24384_),
    .B(_24385_),
    .C1(_22821_),
    .C2(_11197_),
    .ZN(_24386_));
 NAND3_X4 _55598_ (.A1(_23008_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [410]),
    .A3(_23057_),
    .ZN(_24387_));
 NAND3_X2 _55599_ (.A1(_23059_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2174]),
    .A3(_23006_),
    .ZN(_24388_));
 NAND3_X1 _55600_ (.A1(_22944_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2272]),
    .A3(_23561_),
    .ZN(_24389_));
 NAND3_X2 _55601_ (.A1(_23536_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2223]),
    .A3(_23561_),
    .ZN(_24390_));
 NAND4_X4 _55602_ (.A1(_24387_),
    .A2(_24388_),
    .A3(_24389_),
    .A4(_24390_),
    .ZN(_24391_));
 NAND3_X4 _55603_ (.A1(_24045_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1341]),
    .A3(_24026_),
    .ZN(_24392_));
 NAND3_X1 _55604_ (.A1(_23140_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2468]),
    .A3(_23134_),
    .ZN(_24393_));
 NAND3_X4 _55605_ (.A1(_23888_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [704]),
    .A3(_23201_),
    .ZN(_24394_));
 NAND3_X1 _55606_ (.A1(_23036_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2419]),
    .A3(_23026_),
    .ZN(_24395_));
 NAND4_X1 _55607_ (.A1(_24392_),
    .A2(_24393_),
    .A3(_24394_),
    .A4(_24395_),
    .ZN(_24396_));
 NAND3_X2 _55608_ (.A1(_23020_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2125]),
    .A3(_24052_),
    .ZN(_24397_));
 NAND3_X4 _55609_ (.A1(_23236_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [361]),
    .A3(_22959_),
    .ZN(_24398_));
 NAND3_X2 _55610_ (.A1(_23236_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2321]),
    .A3(_23832_),
    .ZN(_24399_));
 NAND3_X2 _55611_ (.A1(_23837_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1978]),
    .A3(_23832_),
    .ZN(_24400_));
 NAND4_X4 _55612_ (.A1(_24397_),
    .A2(_24398_),
    .A3(_24399_),
    .A4(_24400_),
    .ZN(_24401_));
 NOR4_X1 _55613_ (.A1(_24386_),
    .A2(_24391_),
    .A3(_24396_),
    .A4(_24401_),
    .ZN(_24402_));
 NAND3_X4 _55614_ (.A1(_22985_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [557]),
    .A3(_11127_),
    .ZN(_24403_));
 NAND3_X4 _55615_ (.A1(_22242_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1439]),
    .A3(_23051_),
    .ZN(_24404_));
 NAND3_X2 _55616_ (.A1(_22524_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [900]),
    .A3(_23880_),
    .ZN(_24405_));
 NAND3_X4 _55617_ (.A1(_23368_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1390]),
    .A3(_22945_),
    .ZN(_24406_));
 NAND4_X4 _55618_ (.A1(_24403_),
    .A2(_24404_),
    .A3(_24405_),
    .A4(_24406_),
    .ZN(_24407_));
 NAND3_X1 _55619_ (.A1(_24126_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [753]),
    .A3(_23057_),
    .ZN(_24408_));
 NAND3_X2 _55620_ (.A1(_23059_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [606]),
    .A3(_23060_),
    .ZN(_24409_));
 NAND3_X4 _55621_ (.A1(_23011_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2958]),
    .A3(_23128_),
    .ZN(_24410_));
 NAND3_X4 _55622_ (.A1(_24029_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [655]),
    .A3(_23063_),
    .ZN(_24411_));
 NAND4_X4 _55623_ (.A1(_24408_),
    .A2(_24409_),
    .A3(_24410_),
    .A4(_24411_),
    .ZN(_24412_));
 NAND3_X4 _55624_ (.A1(_23560_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1929]),
    .A3(_23009_),
    .ZN(_24413_));
 NAND3_X1 _55625_ (.A1(_22972_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [312]),
    .A3(_22959_),
    .ZN(_24414_));
 NAND3_X1 _55626_ (.A1(_23194_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [18]),
    .A3(_22959_),
    .ZN(_24415_));
 NAND3_X1 _55627_ (.A1(_23271_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [214]),
    .A3(_23196_),
    .ZN(_24416_));
 NAND4_X2 _55628_ (.A1(_24413_),
    .A2(_24414_),
    .A3(_24415_),
    .A4(_24416_),
    .ZN(_24417_));
 NAND3_X4 _55629_ (.A1(_10844_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1782]),
    .A3(_23141_),
    .ZN(_24418_));
 NAND3_X1 _55630_ (.A1(_22975_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [263]),
    .A3(_22959_),
    .ZN(_24419_));
 NAND3_X4 _55631_ (.A1(_23028_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1096]),
    .A3(_23547_),
    .ZN(_24420_));
 NAND3_X2 _55632_ (.A1(_23426_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [67]),
    .A3(_23086_),
    .ZN(_24421_));
 NAND4_X2 _55633_ (.A1(_24418_),
    .A2(_24419_),
    .A3(_24420_),
    .A4(_24421_),
    .ZN(_24422_));
 NOR4_X4 _55634_ (.A1(_24407_),
    .A2(_24412_),
    .A3(_24417_),
    .A4(_24422_),
    .ZN(_24423_));
 NAND3_X1 _55635_ (.A1(_22988_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1733]),
    .A3(_10990_),
    .ZN(_24424_));
 NAND3_X2 _55636_ (.A1(_22994_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1586]),
    .A3(_23116_),
    .ZN(_24425_));
 NAND3_X2 _55637_ (.A1(_22944_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1880]),
    .A3(_23116_),
    .ZN(_24426_));
 NAND3_X2 _55638_ (.A1(_23377_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1635]),
    .A3(_23116_),
    .ZN(_24427_));
 NAND4_X4 _55639_ (.A1(_24424_),
    .A2(_24425_),
    .A3(_24426_),
    .A4(_24427_),
    .ZN(_24428_));
 NAND3_X2 _55640_ (.A1(_23125_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [949]),
    .A3(_23882_),
    .ZN(_24429_));
 NAND3_X1 _55641_ (.A1(_23062_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [851]),
    .A3(_23882_),
    .ZN(_24430_));
 NAND3_X4 _55642_ (.A1(_23062_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [459]),
    .A3(_23063_),
    .ZN(_24431_));
 NAND3_X2 _55643_ (.A1(_23016_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [508]),
    .A3(_23063_),
    .ZN(_24432_));
 NAND4_X4 _55644_ (.A1(_24429_),
    .A2(_24430_),
    .A3(_24431_),
    .A4(_24432_),
    .ZN(_24433_));
 NAND3_X2 _55645_ (.A1(_23192_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2566]),
    .A3(_23068_),
    .ZN(_24434_));
 NAND3_X1 _55646_ (.A1(_23194_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2370]),
    .A3(_23026_),
    .ZN(_24435_));
 NAND3_X2 _55647_ (.A1(_22961_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2664]),
    .A3(_23143_),
    .ZN(_24436_));
 NAND3_X4 _55648_ (.A1(_22978_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3007]),
    .A3(_23037_),
    .ZN(_24437_));
 NAND4_X4 _55649_ (.A1(_24434_),
    .A2(_24435_),
    .A3(_24436_),
    .A4(_24437_),
    .ZN(_24438_));
 NAND3_X2 _55650_ (.A1(_23032_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [802]),
    .A3(_22973_),
    .ZN(_24439_));
 NAND3_X4 _55651_ (.A1(_23039_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1684]),
    .A3(_23146_),
    .ZN(_24440_));
 NAND3_X4 _55652_ (.A1(_23575_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1831]),
    .A3(_23146_),
    .ZN(_24441_));
 NAND3_X4 _55653_ (.A1(_23575_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1047]),
    .A3(_23317_),
    .ZN(_24442_));
 NAND4_X4 _55654_ (.A1(_24439_),
    .A2(_24440_),
    .A3(_24441_),
    .A4(_24442_),
    .ZN(_24443_));
 NOR4_X4 _55655_ (.A1(_24428_),
    .A2(_24433_),
    .A3(_24438_),
    .A4(_24443_),
    .ZN(_24444_));
 NAND4_X1 _55656_ (.A1(_24383_),
    .A2(_24402_),
    .A3(_24423_),
    .A4(_24444_),
    .ZN(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [18]));
 NAND3_X4 _55657_ (.A1(_10779_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2126]),
    .A3(_10940_),
    .ZN(_24445_));
 NAND3_X1 _55658_ (.A1(_10867_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2028]),
    .A3(_22913_),
    .ZN(_24446_));
 NAND2_X4 _55659_ (.A1(_24445_),
    .A2(_24446_),
    .ZN(_24447_));
 AOI221_X4 _55660_ (.A(_24447_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1440]),
    .B2(_22232_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1097]),
    .C2(_23333_),
    .ZN(_24448_));
 NAND3_X1 _55661_ (.A1(_22907_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [803]),
    .A3(_22905_),
    .ZN(_24449_));
 NAND3_X4 _55662_ (.A1(_23721_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2469]),
    .A3(_23481_),
    .ZN(_24450_));
 NAND2_X1 _55663_ (.A1(_24449_),
    .A2(_24450_),
    .ZN(_24451_));
 AOI221_X4 _55664_ (.A(_24451_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1244]),
    .B2(_11065_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [950]),
    .C2(_23047_),
    .ZN(_24452_));
 NAND3_X1 _55665_ (.A1(_23153_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2959]),
    .A3(_23498_),
    .ZN(_24453_));
 NAND3_X2 _55666_ (.A1(_10829_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3008]),
    .A3(_23498_),
    .ZN(_24454_));
 NAND2_X4 _55667_ (.A1(_24453_),
    .A2(_24454_),
    .ZN(_24455_));
 AOI221_X4 _55668_ (.A(_24455_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [656]),
    .B2(_22642_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [754]),
    .C2(_22597_),
    .ZN(_24456_));
 NAND3_X1 _55669_ (.A1(_23721_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1685]),
    .A3(_22921_),
    .ZN(_24457_));
 NAND3_X1 _55670_ (.A1(_23775_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1636]),
    .A3(_22923_),
    .ZN(_24458_));
 NAND2_X1 _55671_ (.A1(_24457_),
    .A2(_24458_),
    .ZN(_24459_));
 AOI221_X4 _55672_ (.A(_24459_),
    .B1(_11003_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1783]),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1587]),
    .C2(_23395_),
    .ZN(_24460_));
 AND4_X2 _55673_ (.A1(_24448_),
    .A2(_24452_),
    .A3(_24456_),
    .A4(_24460_),
    .ZN(_24461_));
 NAND3_X1 _55674_ (.A1(_23150_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [362]),
    .A3(_23643_),
    .ZN(_24462_));
 NAND3_X4 _55675_ (.A1(_22920_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [705]),
    .A3(_23151_),
    .ZN(_24463_));
 NAND2_X4 _55676_ (.A1(_24462_),
    .A2(_24463_),
    .ZN(_24464_));
 AOI221_X2 _55677_ (.A(_24464_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2518]),
    .B2(_10912_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2420]),
    .C2(_10922_),
    .ZN(_24465_));
 NAND3_X2 _55678_ (.A1(_22915_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [852]),
    .A3(_23494_),
    .ZN(_24466_));
 BUF_X32 _55679_ (.A(_10901_),
    .Z(_24467_));
 NAND3_X2 _55680_ (.A1(_24467_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1048]),
    .A3(_23494_),
    .ZN(_24468_));
 NAND2_X4 _55681_ (.A1(_24466_),
    .A2(_24468_),
    .ZN(_24469_));
 AOI221_X4 _55682_ (.A(_24469_),
    .B1(_22910_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2077]),
    .C1(_23467_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1734]),
    .ZN(_24470_));
 NAND3_X2 _55683_ (.A1(_23518_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2567]),
    .A3(_23481_),
    .ZN(_24471_));
 NAND3_X2 _55684_ (.A1(_24467_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2616]),
    .A3(_23012_),
    .ZN(_24472_));
 NAND2_X4 _55685_ (.A1(_24471_),
    .A2(_24472_),
    .ZN(_24473_));
 AOI221_X4 _55686_ (.A(_24473_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [999]),
    .B2(_11094_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1146]),
    .C2(_23331_),
    .ZN(_24474_));
 NAND3_X4 _55687_ (.A1(_23524_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [313]),
    .A3(_23258_),
    .ZN(_24475_));
 NAND3_X2 _55688_ (.A1(_23733_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [460]),
    .A3(_23255_),
    .ZN(_24476_));
 NAND2_X1 _55689_ (.A1(_24475_),
    .A2(_24476_),
    .ZN(_24477_));
 AOI221_X4 _55690_ (.A(_24477_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [264]),
    .B2(_22777_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [607]),
    .C2(_23515_),
    .ZN(_24478_));
 AND4_X1 _55691_ (.A1(_24465_),
    .A2(_24470_),
    .A3(_24474_),
    .A4(_24478_),
    .ZN(_24479_));
 NAND3_X4 _55692_ (.A1(_22985_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [558]),
    .A3(_22995_),
    .ZN(_24480_));
 NAND3_X4 _55693_ (.A1(_22988_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2910]),
    .A3(_22991_),
    .ZN(_24481_));
 NAND3_X4 _55694_ (.A1(_22994_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [411]),
    .A3(_22995_),
    .ZN(_24482_));
 NAND3_X4 _55695_ (.A1(_22944_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3057]),
    .A3(_23000_),
    .ZN(_24483_));
 NAND4_X4 _55696_ (.A1(_24480_),
    .A2(_24481_),
    .A3(_24482_),
    .A4(_24483_),
    .ZN(_24484_));
 NAND3_X2 _55697_ (.A1(_23054_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2322]),
    .A3(_23006_),
    .ZN(_24485_));
 NAND3_X2 _55698_ (.A1(_22950_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2714]),
    .A3(_23131_),
    .ZN(_24486_));
 NAND3_X2 _55699_ (.A1(_22968_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2371]),
    .A3(_23014_),
    .ZN(_24487_));
 NAND3_X2 _55700_ (.A1(_24050_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2665]),
    .A3(_23068_),
    .ZN(_24488_));
 NAND4_X4 _55701_ (.A1(_24485_),
    .A2(_24486_),
    .A3(_24487_),
    .A4(_24488_),
    .ZN(_24489_));
 NAND3_X4 _55702_ (.A1(_23560_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1930]),
    .A3(_23009_),
    .ZN(_24490_));
 NAND3_X2 _55703_ (.A1(_23189_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2812]),
    .A3(_10790_),
    .ZN(_24491_));
 NAND3_X2 _55704_ (.A1(_23025_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2861]),
    .A3(_10790_),
    .ZN(_24492_));
 NAND3_X2 _55705_ (.A1(_23837_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2763]),
    .A3(_23037_),
    .ZN(_24493_));
 NAND4_X4 _55706_ (.A1(_24490_),
    .A2(_24491_),
    .A3(_24492_),
    .A4(_24493_),
    .ZN(_24494_));
 NAND3_X2 _55707_ (.A1(_23032_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1979]),
    .A3(_23894_),
    .ZN(_24495_));
 NAND3_X2 _55708_ (.A1(_23276_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2175]),
    .A3(_23832_),
    .ZN(_24496_));
 NAND3_X2 _55709_ (.A1(_23280_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1881]),
    .A3(_23146_),
    .ZN(_24497_));
 NAND3_X2 _55710_ (.A1(_23575_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1832]),
    .A3(_23576_),
    .ZN(_24498_));
 NAND4_X4 _55711_ (.A1(_24495_),
    .A2(_24496_),
    .A3(_24497_),
    .A4(_24498_),
    .ZN(_24499_));
 NOR4_X1 _55712_ (.A1(_24484_),
    .A2(_24489_),
    .A3(_24494_),
    .A4(_24499_),
    .ZN(_24500_));
 NAND3_X1 _55713_ (.A1(_22907_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1195]),
    .A3(_11035_),
    .ZN(_24501_));
 NAND3_X4 _55714_ (.A1(_23775_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [68]),
    .A3(_11174_),
    .ZN(_24502_));
 NAND2_X1 _55715_ (.A1(_24501_),
    .A2(_24502_),
    .ZN(_24503_));
 AOI221_X4 _55716_ (.A(_24503_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1391]),
    .B2(_23094_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1538]),
    .C2(_23179_),
    .ZN(_24504_));
 NAND3_X1 _55717_ (.A1(_10856_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [901]),
    .A3(_23804_),
    .ZN(_24505_));
 NAND3_X1 _55718_ (.A1(_23173_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1293]),
    .A3(_23701_),
    .ZN(_24506_));
 NAND2_X1 _55719_ (.A1(_24505_),
    .A2(_24506_),
    .ZN(_24507_));
 AOI221_X4 _55720_ (.A(_24507_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [509]),
    .B2(_11152_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1342]),
    .C2(_23748_),
    .ZN(_24508_));
 NAND3_X1 _55721_ (.A1(_23935_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2273]),
    .A3(_23553_),
    .ZN(_24509_));
 NAND3_X4 _55722_ (.A1(_23390_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3106]),
    .A3(_22999_),
    .ZN(_24510_));
 NAND3_X4 _55723_ (.A1(_10818_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1489]),
    .A3(_23608_),
    .ZN(_24511_));
 NAND3_X1 _55724_ (.A1(_23303_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2224]),
    .A3(_23005_),
    .ZN(_24512_));
 AND4_X4 _55725_ (.A1(_24509_),
    .A2(_24510_),
    .A3(_24511_),
    .A4(_24512_),
    .ZN(_24513_));
 NAND3_X1 _55726_ (.A1(_10879_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [19]),
    .A3(_23250_),
    .ZN(_24514_));
 NAND3_X1 _55727_ (.A1(_23003_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [166]),
    .A3(_22939_),
    .ZN(_24515_));
 NAND3_X1 _55728_ (.A1(_23306_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [117]),
    .A3(_22939_),
    .ZN(_24516_));
 NAND3_X1 _55729_ (.A1(_22932_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [215]),
    .A3(_11175_),
    .ZN(_24517_));
 AND4_X4 _55730_ (.A1(_24514_),
    .A2(_24515_),
    .A3(_24516_),
    .A4(_24517_),
    .ZN(_24518_));
 AND4_X1 _55731_ (.A1(_24504_),
    .A2(_24508_),
    .A3(_24513_),
    .A4(_24518_),
    .ZN(_24519_));
 NAND4_X1 _55732_ (.A1(_24461_),
    .A2(_24479_),
    .A3(_24500_),
    .A4(_24519_),
    .ZN(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [19]));
 AND3_X1 _55733_ (.A1(_23288_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1294]),
    .A3(_22898_),
    .ZN(_24520_));
 AOI221_X4 _55734_ (.A(_24520_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1245]),
    .B2(_23048_),
    .C1(_22282_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1343]),
    .ZN(_24521_));
 NAND3_X1 _55735_ (.A1(_23408_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [706]),
    .A3(_11124_),
    .ZN(_24522_));
 OAI221_X2 _55736_ (.A(_24522_),
    .B1(_11142_),
    .B2(_22676_),
    .C1(_11121_),
    .C2(_22612_),
    .ZN(_24523_));
 AOI221_X2 _55737_ (.A(_24523_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [657]),
    .B2(_22642_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [412]),
    .C2(_23610_),
    .ZN(_24524_));
 NAND3_X1 _55738_ (.A1(_10842_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1392]),
    .A3(_22979_),
    .ZN(_24525_));
 OAI221_X2 _55739_ (.A(_24525_),
    .B1(_11042_),
    .B2(_22223_),
    .C1(_11032_),
    .C2(_22196_),
    .ZN(_24526_));
 AOI221_X2 _55740_ (.A(_24526_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1441]),
    .B2(_22232_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1196]),
    .C2(_23103_),
    .ZN(_24527_));
 AND3_X1 _55741_ (.A1(_10797_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [363]),
    .A3(_11185_),
    .ZN(_24528_));
 AND3_X1 _55742_ (.A1(_10811_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [314]),
    .A3(_11185_),
    .ZN(_24529_));
 AND3_X1 _55743_ (.A1(_10901_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [265]),
    .A3(_11185_),
    .ZN(_24530_));
 OR3_X1 _55744_ (.A1(_24528_),
    .A2(_24529_),
    .A3(_24530_),
    .ZN(_24531_));
 AOI221_X2 _55745_ (.A(_24531_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [216]),
    .B2(_11190_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [69]),
    .C2(_23714_),
    .ZN(_24532_));
 AND4_X4 _55746_ (.A1(_24521_),
    .A2(net29),
    .A3(net28),
    .A4(net49),
    .ZN(_24533_));
 AOI22_X4 _55747_ (.A1(_23587_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2519]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2470]),
    .B2(_21705_),
    .ZN(_24534_));
 AOI22_X4 _55748_ (.A1(_23213_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2911]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2862]),
    .B2(_21502_),
    .ZN(_24535_));
 NAND3_X2 _55749_ (.A1(_10880_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2372]),
    .A3(_10893_),
    .ZN(_24536_));
 NAND3_X2 _55750_ (.A1(_10869_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2813]),
    .A3(_23361_),
    .ZN(_24537_));
 NAND4_X4 _55751_ (.A1(_24534_),
    .A2(_24535_),
    .A3(_24536_),
    .A4(_24537_),
    .ZN(_24538_));
 AOI22_X2 _55752_ (.A1(_10800_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3107]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3058]),
    .B2(_10813_),
    .ZN(_24539_));
 NAND3_X2 _55753_ (.A1(_23340_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2960]),
    .A3(_22991_),
    .ZN(_24540_));
 NAND3_X2 _55754_ (.A1(_22242_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3009]),
    .A3(_22991_),
    .ZN(_24541_));
 NAND3_X2 _55755_ (.A1(_22994_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2764]),
    .A3(_23000_),
    .ZN(_24542_));
 NAND4_X4 _55756_ (.A1(_24539_),
    .A2(_24540_),
    .A3(_24541_),
    .A4(_24542_),
    .ZN(_24543_));
 AOI22_X4 _55757_ (.A1(_23373_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2715]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2666]),
    .B2(_23374_),
    .ZN(_24544_));
 NAND3_X1 _55758_ (.A1(_23114_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2421]),
    .A3(_23120_),
    .ZN(_24545_));
 NAND3_X1 _55759_ (.A1(_22998_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2617]),
    .A3(_23120_),
    .ZN(_24546_));
 NAND3_X1 _55760_ (.A1(_23368_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2568]),
    .A3(_23120_),
    .ZN(_24547_));
 NAND4_X1 _55761_ (.A1(_24544_),
    .A2(_24545_),
    .A3(_24546_),
    .A4(_24547_),
    .ZN(_24548_));
 NOR3_X1 _55762_ (.A1(_24538_),
    .A2(_24543_),
    .A3(_24548_),
    .ZN(_24549_));
 AND3_X1 _55763_ (.A1(_23509_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [167]),
    .A3(_11174_),
    .ZN(_24550_));
 AOI221_X4 _55764_ (.A(_24550_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [118]),
    .B2(_23453_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [20]),
    .C2(_23164_),
    .ZN(_24551_));
 NAND3_X1 _55765_ (.A1(_10868_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [853]),
    .A3(_23329_),
    .ZN(_24552_));
 AOI22_X1 _55766_ (.A1(_23047_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [951]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [902]),
    .B2(_23265_),
    .ZN(_24553_));
 NAND3_X1 _55767_ (.A1(_10879_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [804]),
    .A3(_11081_),
    .ZN(_24554_));
 NAND3_X1 _55768_ (.A1(_23252_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1049]),
    .A3(_11081_),
    .ZN(_24555_));
 AND4_X1 _55769_ (.A1(_24552_),
    .A2(_24553_),
    .A3(_24554_),
    .A4(_24555_),
    .ZN(_24556_));
 AND3_X1 _55770_ (.A1(_23176_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [461]),
    .A3(_23255_),
    .ZN(_24557_));
 AOI221_X4 _55771_ (.A(_24557_),
    .B1(_11152_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [510]),
    .C1(_11147_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [559]),
    .ZN(_24558_));
 AND3_X1 _55772_ (.A1(_23459_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1147]),
    .A3(_23460_),
    .ZN(_24559_));
 AOI221_X2 _55773_ (.A(_24559_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1098]),
    .B2(_23332_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1000]),
    .C2(_23104_),
    .ZN(_24560_));
 AND4_X4 _55774_ (.A1(_24551_),
    .A2(_24556_),
    .A3(_24558_),
    .A4(_24560_),
    .ZN(_24561_));
 AOI22_X4 _55775_ (.A1(_23097_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2323]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2274]),
    .B2(_21816_),
    .ZN(_24562_));
 OAI221_X2 _55776_ (.A(_24562_),
    .B1(_21855_),
    .B2(_10951_),
    .C1(_21872_),
    .C2(_10957_),
    .ZN(_24563_));
 AND3_X1 _55777_ (.A1(_23041_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2029]),
    .A3(_10940_),
    .ZN(_24564_));
 AOI21_X2 _55778_ (.A(_24564_),
    .B1(_23485_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1980]),
    .ZN(_24565_));
 NAND3_X2 _55779_ (.A1(_23016_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2078]),
    .A3(_24046_),
    .ZN(_24566_));
 OAI211_X4 _55780_ (.A(_24565_),
    .B(_24566_),
    .C1(_10963_),
    .C2(_21892_),
    .ZN(_24567_));
 NAND3_X4 _55781_ (.A1(_23236_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1931]),
    .A3(_23146_),
    .ZN(_24568_));
 OAI221_X2 _55782_ (.A(_24568_),
    .B1(_22055_),
    .B2(_10998_),
    .C1(_10994_),
    .C2(_22021_),
    .ZN(_24569_));
 AOI22_X4 _55783_ (.A1(_23595_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1588]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1637]),
    .B2(_23604_),
    .ZN(_24570_));
 NAND3_X1 _55784_ (.A1(_23039_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1686]),
    .A3(_23146_),
    .ZN(_24571_));
 NAND3_X2 _55785_ (.A1(_23421_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1735]),
    .A3(_23576_),
    .ZN(_24572_));
 NAND3_X1 _55786_ (.A1(_23839_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1784]),
    .A3(_23576_),
    .ZN(_24573_));
 NAND4_X4 _55787_ (.A1(_24570_),
    .A2(_24571_),
    .A3(_24572_),
    .A4(_24573_),
    .ZN(_24574_));
 NOR4_X4 _55788_ (.A1(_24563_),
    .A2(_24567_),
    .A3(_24569_),
    .A4(_24574_),
    .ZN(_24575_));
 NAND4_X1 _55789_ (.A1(_24533_),
    .A2(_24549_),
    .A3(_24561_),
    .A4(_24575_),
    .ZN(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [20]));
 AND3_X1 _55790_ (.A1(_22897_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [756]),
    .A3(_23504_),
    .ZN(_24576_));
 AOI221_X2 _55791_ (.A(_24576_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [707]),
    .B2(_11131_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [609]),
    .C2(_23106_),
    .ZN(_24577_));
 NAND3_X1 _55792_ (.A1(_23084_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1197]),
    .A3(_11036_),
    .ZN(_24578_));
 OAI21_X1 _55793_ (.A(_24578_),
    .B1(_11066_),
    .B2(_22344_),
    .ZN(_24579_));
 OAI22_X2 _55794_ (.A1(_11055_),
    .A2(_22296_),
    .B1(_22321_),
    .B2(_11061_),
    .ZN(_24580_));
 AOI211_X2 _55795_ (.A(_24579_),
    .B(_24580_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1442]),
    .C2(_23326_),
    .ZN(_24581_));
 NAND3_X1 _55796_ (.A1(_23207_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [413]),
    .A3(_23237_),
    .ZN(_24582_));
 AOI22_X2 _55797_ (.A1(_23622_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [560]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [511]),
    .B2(_23689_),
    .ZN(_24583_));
 NAND3_X1 _55798_ (.A1(_23113_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [462]),
    .A3(_23346_),
    .ZN(_24584_));
 NAND3_X1 _55799_ (.A1(_22997_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [658]),
    .A3(_23346_),
    .ZN(_24585_));
 AND4_X4 _55800_ (.A1(_24582_),
    .A2(_24583_),
    .A3(_24584_),
    .A4(_24585_),
    .ZN(_24586_));
 AND3_X1 _55801_ (.A1(_23518_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1393]),
    .A3(_23848_),
    .ZN(_24587_));
 AOI221_X4 _55802_ (.A(_24587_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1491]),
    .B2(_22210_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1540]),
    .C2(_23179_),
    .ZN(_24588_));
 AND4_X4 _55803_ (.A1(net48),
    .A2(_24581_),
    .A3(_24586_),
    .A4(_24588_),
    .ZN(_24589_));
 NAND3_X1 _55804_ (.A1(_24262_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2324]),
    .A3(_23600_),
    .ZN(_24590_));
 AOI22_X2 _55805_ (.A1(_10956_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2177]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2030]),
    .B2(_23156_),
    .ZN(_24591_));
 NAND3_X1 _55806_ (.A1(_23385_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2226]),
    .A3(_10941_),
    .ZN(_24592_));
 NAND3_X1 _55807_ (.A1(_23935_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2275]),
    .A3(_10941_),
    .ZN(_24593_));
 AND4_X4 _55808_ (.A1(_24590_),
    .A2(_24591_),
    .A3(_24592_),
    .A4(_24593_),
    .ZN(_24594_));
 NAND3_X1 _55809_ (.A1(_23245_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1932]),
    .A3(_23576_),
    .ZN(_24595_));
 AOI22_X2 _55810_ (.A1(_11003_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1785]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1638]),
    .B2(_23396_),
    .ZN(_24596_));
 NAND3_X1 _55811_ (.A1(_10818_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1883]),
    .A3(_10989_),
    .ZN(_24597_));
 NAND3_X1 _55812_ (.A1(_23252_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1834]),
    .A3(_10989_),
    .ZN(_24598_));
 AND4_X1 _55813_ (.A1(_24595_),
    .A2(_24596_),
    .A3(_24597_),
    .A4(_24598_),
    .ZN(_24599_));
 AND3_X1 _55814_ (.A1(_23173_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1687]),
    .A3(_23662_),
    .ZN(_24600_));
 AOI221_X4 _55815_ (.A(_24600_),
    .B1(_11025_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1589]),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1736]),
    .C2(_22078_),
    .ZN(_24601_));
 AND3_X1 _55816_ (.A1(_23083_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1981]),
    .A3(_23169_),
    .ZN(_24602_));
 AOI221_X2 _55817_ (.A(_24602_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2079]),
    .B2(_23233_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2128]),
    .C2(_23736_),
    .ZN(_24603_));
 AND4_X4 _55818_ (.A1(_24594_),
    .A2(_24599_),
    .A3(_24601_),
    .A4(net27),
    .ZN(_24604_));
 NAND3_X1 _55819_ (.A1(_23221_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2569]),
    .A3(_23422_),
    .ZN(_24605_));
 AND3_X1 _55820_ (.A1(_10824_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2618]),
    .A3(_10886_),
    .ZN(_24606_));
 AOI221_X1 _55821_ (.A(_24606_),
    .B1(_21600_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2667]),
    .C1(_21573_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2716]),
    .ZN(_24607_));
 AOI22_X1 _55822_ (.A1(_23587_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2520]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2471]),
    .B2(_21705_),
    .ZN(_24608_));
 AOI22_X2 _55823_ (.A1(_10929_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2373]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2422]),
    .B2(_23301_),
    .ZN(_24609_));
 AND4_X1 _55824_ (.A1(_24605_),
    .A2(_24607_),
    .A3(_24608_),
    .A4(_24609_),
    .ZN(_24610_));
 AND3_X1 _55825_ (.A1(_23721_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2863]),
    .A3(_10788_),
    .ZN(_24611_));
 AOI221_X4 _55826_ (.A(_24611_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2814]),
    .B2(_21536_),
    .C1(_23213_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2912]),
    .ZN(_24612_));
 NAND4_X1 _55827_ (.A1(_10751_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3108]),
    .A3(_10825_),
    .A4(_10795_),
    .ZN(_24613_));
 NAND3_X2 _55828_ (.A1(_24467_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3010]),
    .A3(_23794_),
    .ZN(_24614_));
 NAND4_X1 _55829_ (.A1(_10809_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3059]),
    .A3(_10825_),
    .A4(_10795_),
    .ZN(_24615_));
 NAND3_X1 _55830_ (.A1(_24613_),
    .A2(_24614_),
    .A3(_24615_),
    .ZN(_24616_));
 AOI221_X4 _55831_ (.A(_24616_),
    .B1(_22918_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2961]),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2765]),
    .C2(_21289_),
    .ZN(_24617_));
 AND3_X4 _55832_ (.A1(_24610_),
    .A2(_24612_),
    .A3(_24617_),
    .ZN(_24618_));
 AND3_X1 _55833_ (.A1(_23382_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [805]),
    .A3(_23804_),
    .ZN(_24619_));
 AOI221_X4 _55834_ (.A(_24619_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [903]),
    .B2(_11106_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [952]),
    .C2(_11100_),
    .ZN(_24620_));
 NAND3_X1 _55835_ (.A1(_22993_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [21]),
    .A3(_23246_),
    .ZN(_24621_));
 AND3_X1 _55836_ (.A1(_10901_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [266]),
    .A3(_11185_),
    .ZN(_24622_));
 AOI221_X2 _55837_ (.A(_24622_),
    .B1(_11181_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [315]),
    .C1(_11170_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [364]),
    .ZN(_24623_));
 AOI22_X2 _55838_ (.A1(_22806_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [168]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [119]),
    .B2(_23453_),
    .ZN(_24624_));
 AOI22_X2 _55839_ (.A1(_11190_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [217]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [70]),
    .B2(_11211_),
    .ZN(_24625_));
 AND4_X4 _55840_ (.A1(_24621_),
    .A2(_24623_),
    .A3(_24624_),
    .A4(_24625_),
    .ZN(_24626_));
 AND3_X1 _55841_ (.A1(_23459_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1148]),
    .A3(_23460_),
    .ZN(_24627_));
 AOI221_X2 _55842_ (.A(_24627_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1099]),
    .B2(_23332_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1050]),
    .C2(_22435_),
    .ZN(_24628_));
 AOI22_X2 _55843_ (.A1(_22459_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1001]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [854]),
    .B2(_23268_),
    .ZN(_24629_));
 AND4_X4 _55844_ (.A1(_24620_),
    .A2(_24626_),
    .A3(_24628_),
    .A4(_24629_),
    .ZN(_24630_));
 NAND4_X1 _55845_ (.A1(_24589_),
    .A2(_24604_),
    .A3(_24618_),
    .A4(_24630_),
    .ZN(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [21]));
 AND3_X1 _55846_ (.A1(_23019_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [169]),
    .A3(_11175_),
    .ZN(_24631_));
 AOI21_X4 _55847_ (.A(_24631_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [120]),
    .B2(_22827_),
    .ZN(_24632_));
 OAI221_X2 _55848_ (.A(_24632_),
    .B1(_22653_),
    .B2(_11137_),
    .C1(_22786_),
    .C2(_11187_),
    .ZN(_24633_));
 AND4_X2 _55849_ (.A1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3060]),
    .A2(_10809_),
    .A3(_22989_),
    .A4(_10795_),
    .ZN(_24634_));
 AOI21_X4 _55850_ (.A(_24634_),
    .B1(_10800_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3109]),
    .ZN(_24635_));
 OAI221_X2 _55851_ (.A(_24635_),
    .B1(_22712_),
    .B2(_11154_),
    .C1(_22872_),
    .C2(_11207_),
    .ZN(_24636_));
 AOI22_X4 _55852_ (.A1(_23485_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1982]),
    .B1(_23591_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1688]),
    .ZN(_24637_));
 NAND3_X2 _55853_ (.A1(_23127_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1492]),
    .A3(_24026_),
    .ZN(_24638_));
 OAI211_X4 _55854_ (.A(_24637_),
    .B(_24638_),
    .C1(_22199_),
    .C2(_11032_),
    .ZN(_24639_));
 NAND3_X4 _55855_ (.A1(_23008_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2374]),
    .A3(_23131_),
    .ZN(_24640_));
 NAND3_X4 _55856_ (.A1(_23011_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [610]),
    .A3(_23060_),
    .ZN(_24641_));
 NAND3_X4 _55857_ (.A1(_22958_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1835]),
    .A3(_23141_),
    .ZN(_24642_));
 NAND3_X1 _55858_ (.A1(_23888_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [316]),
    .A3(_23835_),
    .ZN(_24643_));
 NAND4_X1 _55859_ (.A1(_24640_),
    .A2(_24641_),
    .A3(_24642_),
    .A4(_24643_),
    .ZN(_24644_));
 NOR4_X1 _55860_ (.A1(_24633_),
    .A2(_24636_),
    .A3(_24639_),
    .A4(_24644_),
    .ZN(_24645_));
 NAND3_X4 _55861_ (.A1(_23150_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [757]),
    .A3(_23504_),
    .ZN(_24646_));
 NAND3_X4 _55862_ (.A1(_22920_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2668]),
    .A3(_23481_),
    .ZN(_24647_));
 NAND2_X4 _55863_ (.A1(_24646_),
    .A2(_24647_),
    .ZN(_24648_));
 AOI221_X4 _55864_ (.A(_24648_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1933]),
    .B2(_21978_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1786]),
    .C2(_11003_),
    .ZN(_24649_));
 NAND3_X1 _55865_ (.A1(_23509_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1737]),
    .A3(_22921_),
    .ZN(_24650_));
 NAND3_X1 _55866_ (.A1(_23751_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2276]),
    .A3(_23657_),
    .ZN(_24651_));
 NAND2_X1 _55867_ (.A1(_24650_),
    .A2(_24651_),
    .ZN(_24652_));
 AOI221_X2 _55868_ (.A(_24652_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2129]),
    .B2(_23736_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1590]),
    .C2(_23395_),
    .ZN(_24653_));
 NAND3_X4 _55869_ (.A1(_23487_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [365]),
    .A3(_23159_),
    .ZN(_24654_));
 NAND3_X1 _55870_ (.A1(_23733_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1247]),
    .A3(_23848_),
    .ZN(_24655_));
 NAND2_X2 _55871_ (.A1(_24654_),
    .A2(_24655_),
    .ZN(_24656_));
 AOI221_X2 _55872_ (.A(_24656_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1884]),
    .B2(_10993_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1198]),
    .C2(_23103_),
    .ZN(_24657_));
 NAND3_X4 _55873_ (.A1(_23166_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2521]),
    .A3(_23012_),
    .ZN(_24658_));
 NAND3_X1 _55874_ (.A1(_23733_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1639]),
    .A3(_23662_),
    .ZN(_24659_));
 NAND2_X1 _55875_ (.A1(_24658_),
    .A2(_24659_),
    .ZN(_24660_));
 AOI221_X4 _55876_ (.A(_24660_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2080]),
    .B2(_10968_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2031]),
    .C2(_23156_),
    .ZN(_24661_));
 AND4_X4 _55877_ (.A1(_24649_),
    .A2(_24653_),
    .A3(_24657_),
    .A4(_24661_),
    .ZN(_24662_));
 NAND3_X2 _55878_ (.A1(_22985_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [561]),
    .A3(_22995_),
    .ZN(_24663_));
 NAND3_X2 _55879_ (.A1(_23114_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [463]),
    .A3(_22995_),
    .ZN(_24664_));
 NAND3_X4 _55880_ (.A1(_22994_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2766]),
    .A3(_23000_),
    .ZN(_24665_));
 NAND3_X4 _55881_ (.A1(_10858_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2864]),
    .A3(_23123_),
    .ZN(_24666_));
 NAND4_X4 _55882_ (.A1(_24663_),
    .A2(_24664_),
    .A3(_24665_),
    .A4(_24666_),
    .ZN(_24667_));
 NAND3_X2 _55883_ (.A1(_23004_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [953]),
    .A3(_23880_),
    .ZN(_24668_));
 NAND3_X4 _55884_ (.A1(_23125_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2913]),
    .A3(_23123_),
    .ZN(_24669_));
 NAND3_X2 _55885_ (.A1(_23011_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1002]),
    .A3(_23882_),
    .ZN(_24670_));
 NAND3_X2 _55886_ (.A1(_23133_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [806]),
    .A3(_22970_),
    .ZN(_24671_));
 NAND4_X4 _55887_ (.A1(_24668_),
    .A2(_24669_),
    .A3(_24670_),
    .A4(_24671_),
    .ZN(_24672_));
 NAND3_X2 _55888_ (.A1(_23560_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1149]),
    .A3(_23882_),
    .ZN(_24673_));
 NAND3_X4 _55889_ (.A1(_23022_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [414]),
    .A3(_23201_),
    .ZN(_24674_));
 NAND3_X2 _55890_ (.A1(_22975_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1051]),
    .A3(_22976_),
    .ZN(_24675_));
 NAND3_X2 _55891_ (.A1(_23028_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1100]),
    .A3(_23891_),
    .ZN(_24676_));
 NAND4_X4 _55892_ (.A1(_24673_),
    .A2(_24674_),
    .A3(_24675_),
    .A4(_24676_),
    .ZN(_24677_));
 NAND3_X4 _55893_ (.A1(_10844_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2178]),
    .A3(_23894_),
    .ZN(_24678_));
 NAND3_X4 _55894_ (.A1(_22975_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3011]),
    .A3(_23037_),
    .ZN(_24679_));
 NAND3_X4 _55895_ (.A1(_23039_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [904]),
    .A3(_23547_),
    .ZN(_24680_));
 NAND3_X4 _55896_ (.A1(_23575_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2227]),
    .A3(_23600_),
    .ZN(_24681_));
 NAND4_X4 _55897_ (.A1(_24678_),
    .A2(_24679_),
    .A3(_24680_),
    .A4(_24681_),
    .ZN(_24682_));
 NOR4_X4 _55898_ (.A1(_24667_),
    .A2(_24672_),
    .A3(_24677_),
    .A4(_24682_),
    .ZN(_24683_));
 NAND3_X4 _55899_ (.A1(_10805_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2325]),
    .A3(_23554_),
    .ZN(_24684_));
 NAND3_X4 _55900_ (.A1(_23114_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [855]),
    .A3(_23880_),
    .ZN(_24685_));
 NAND3_X2 _55901_ (.A1(_23114_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2815]),
    .A3(_23000_),
    .ZN(_24686_));
 NAND3_X4 _55902_ (.A1(_22933_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2962]),
    .A3(_23123_),
    .ZN(_24687_));
 NAND4_X4 _55903_ (.A1(_24684_),
    .A2(_24685_),
    .A3(_24686_),
    .A4(_24687_),
    .ZN(_24688_));
 NAND3_X1 _55904_ (.A1(_23125_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1345]),
    .A3(_22945_),
    .ZN(_24689_));
 NAND3_X2 _55905_ (.A1(_10858_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1296]),
    .A3(_24026_),
    .ZN(_24690_));
 NAND3_X4 _55906_ (.A1(_24029_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1443]),
    .A3(_11037_),
    .ZN(_24691_));
 NAND3_X4 _55907_ (.A1(_23189_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [71]),
    .A3(_23187_),
    .ZN(_24692_));
 NAND4_X4 _55908_ (.A1(_24689_),
    .A2(_24690_),
    .A3(_24691_),
    .A4(_24692_),
    .ZN(_24693_));
 NAND3_X1 _55909_ (.A1(_23067_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2717]),
    .A3(_23068_),
    .ZN(_24694_));
 NAND3_X1 _55910_ (.A1(_10844_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [218]),
    .A3(_22959_),
    .ZN(_24695_));
 NAND3_X1 _55911_ (.A1(_23071_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2619]),
    .A3(_23143_),
    .ZN(_24696_));
 NAND3_X4 _55912_ (.A1(_23028_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [708]),
    .A3(_23072_),
    .ZN(_24697_));
 NAND4_X1 _55913_ (.A1(_24694_),
    .A2(_24695_),
    .A3(_24696_),
    .A4(_24697_),
    .ZN(_24698_));
 NAND3_X2 _55914_ (.A1(_10844_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2570]),
    .A3(_23134_),
    .ZN(_24699_));
 NAND3_X4 _55915_ (.A1(_23271_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1394]),
    .A3(_22981_),
    .ZN(_24700_));
 NAND3_X2 _55916_ (.A1(_23042_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2423]),
    .A3(_23043_),
    .ZN(_24701_));
 NAND3_X1 _55917_ (.A1(_23204_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2472]),
    .A3(_23422_),
    .ZN(_24702_));
 NAND4_X4 _55918_ (.A1(_24699_),
    .A2(_24700_),
    .A3(_24701_),
    .A4(_24702_),
    .ZN(_24703_));
 NOR4_X2 _55919_ (.A1(_24688_),
    .A2(_24693_),
    .A3(_24698_),
    .A4(_24703_),
    .ZN(_24704_));
 NAND4_X1 _55920_ (.A1(_24645_),
    .A2(_24662_),
    .A3(_24683_),
    .A4(_24704_),
    .ZN(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [22]));
 AOI22_X4 _55921_ (.A1(_10800_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3110]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3061]),
    .B2(_10813_),
    .ZN(_24705_));
 NAND3_X1 _55922_ (.A1(_23839_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2963]),
    .A3(_23431_),
    .ZN(_24706_));
 NAND3_X1 _55923_ (.A1(_23575_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3012]),
    .A3(_23431_),
    .ZN(_24707_));
 AND3_X4 _55924_ (.A1(_24705_),
    .A2(_24706_),
    .A3(_24707_),
    .ZN(_24708_));
 NAND3_X2 _55925_ (.A1(_23215_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2228]),
    .A3(_10939_),
    .ZN(_24709_));
 OAI221_X2 _55926_ (.A(_24709_),
    .B1(_10946_),
    .B2(_21836_),
    .C1(_10937_),
    .C2(_21809_),
    .ZN(_24710_));
 AOI221_X2 _55927_ (.A(_24710_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2179]),
    .B2(_10955_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1983]),
    .C2(_23485_),
    .ZN(_24711_));
 NAND3_X2 _55928_ (.A1(_23230_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2767]),
    .A3(_23174_),
    .ZN(_24712_));
 OAI21_X1 _55929_ (.A(_24712_),
    .B1(_10864_),
    .B2(_21551_),
    .ZN(_24713_));
 AOI221_X2 _55930_ (.A(_24713_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2914]),
    .B2(_21466_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2865]),
    .C2(_21502_),
    .ZN(_24714_));
 AND3_X1 _55931_ (.A1(_23806_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2032]),
    .A3(_22962_),
    .ZN(_24715_));
 AOI221_X4 _55932_ (.A(_24715_),
    .B1(_22910_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2081]),
    .C1(_10962_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2130]),
    .ZN(_24716_));
 AND4_X1 _55933_ (.A1(_24708_),
    .A2(net26),
    .A3(_24714_),
    .A4(_24716_),
    .ZN(_24717_));
 NAND3_X2 _55934_ (.A1(_23408_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1493]),
    .A3(_22979_),
    .ZN(_24718_));
 NAND3_X4 _55935_ (.A1(_10842_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1395]),
    .A3(_22979_),
    .ZN(_24719_));
 OAI211_X4 _55936_ (.A(_24718_),
    .B(_24719_),
    .C1(_11032_),
    .C2(_22202_),
    .ZN(_24720_));
 AOI221_X4 _55937_ (.A(_24720_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1444]),
    .B2(_22232_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1199]),
    .C2(_23103_),
    .ZN(_24721_));
 AND3_X1 _55938_ (.A1(_23487_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1150]),
    .A3(_23804_),
    .ZN(_24722_));
 AOI221_X2 _55939_ (.A(_24722_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1101]),
    .B2(_22410_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1003]),
    .C2(_23104_),
    .ZN(_24723_));
 AOI22_X2 _55940_ (.A1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1052]),
    .A2(_23632_),
    .B1(_23268_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [856]),
    .ZN(_24724_));
 NAND3_X1 _55941_ (.A1(_22987_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [954]),
    .A3(_23321_),
    .ZN(_24725_));
 AND3_X1 _55942_ (.A1(_10920_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1248]),
    .A3(_11034_),
    .ZN(_24726_));
 AOI221_X2 _55943_ (.A(_24726_),
    .B1(_11059_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1297]),
    .C1(_11054_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1346]),
    .ZN(_24727_));
 NAND3_X1 _55944_ (.A1(_23455_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [807]),
    .A3(_23879_),
    .ZN(_24728_));
 NAND3_X1 _55945_ (.A1(_23306_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [905]),
    .A3(_23879_),
    .ZN(_24729_));
 AND4_X1 _55946_ (.A1(_24725_),
    .A2(_24727_),
    .A3(_24728_),
    .A4(_24729_),
    .ZN(_24730_));
 AND4_X4 _55947_ (.A1(_24721_),
    .A2(_24723_),
    .A3(_24724_),
    .A4(_24730_),
    .ZN(_24731_));
 NAND3_X1 _55948_ (.A1(_23150_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [366]),
    .A3(_23643_),
    .ZN(_24732_));
 NAND3_X1 _55949_ (.A1(_22942_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [317]),
    .A3(_11174_),
    .ZN(_24733_));
 NAND2_X1 _55950_ (.A1(_24732_),
    .A2(_24733_),
    .ZN(_24734_));
 AOI221_X2 _55951_ (.A(_24734_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [268]),
    .B2(_22777_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [219]),
    .C2(_23248_),
    .ZN(_24735_));
 NAND3_X1 _55952_ (.A1(_23158_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [170]),
    .A3(_23159_),
    .ZN(_24736_));
 NAND3_X1 _55953_ (.A1(_23173_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [121]),
    .A3(_23258_),
    .ZN(_24737_));
 NAND2_X1 _55954_ (.A1(_24736_),
    .A2(_24737_),
    .ZN(_24738_));
 AOI221_X2 _55955_ (.A(_24738_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [23]),
    .B2(_11205_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [72]),
    .C2(_23714_),
    .ZN(_24739_));
 NAND3_X1 _55956_ (.A1(_23242_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [611]),
    .A3(_11126_),
    .ZN(_24740_));
 AOI22_X2 _55957_ (.A1(_11147_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [562]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [513]),
    .B2(_23689_),
    .ZN(_24741_));
 NAND3_X1 _55958_ (.A1(_23293_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [464]),
    .A3(_23056_),
    .ZN(_24742_));
 NAND3_X1 _55959_ (.A1(_23455_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [415]),
    .A3(_23056_),
    .ZN(_24743_));
 AND4_X4 _55960_ (.A1(_24740_),
    .A2(_24741_),
    .A3(_24742_),
    .A4(_24743_),
    .ZN(_24744_));
 AND3_X1 _55961_ (.A1(_23408_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [709]),
    .A3(_23255_),
    .ZN(_24745_));
 AOI221_X4 _55962_ (.A(_24745_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [660]),
    .B2(_22642_),
    .C1(_22597_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [758]),
    .ZN(_24746_));
 AND4_X4 _55963_ (.A1(_24735_),
    .A2(_24739_),
    .A3(_24744_),
    .A4(_24746_),
    .ZN(_24747_));
 AND3_X1 _55964_ (.A1(_23751_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1885]),
    .A3(_22923_),
    .ZN(_24748_));
 AOI221_X4 _55965_ (.A(_24748_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1836]),
    .B2(_23286_),
    .C1(_23584_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1934]),
    .ZN(_24749_));
 NAND3_X1 _55966_ (.A1(_23113_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1640]),
    .A3(_23393_),
    .ZN(_24750_));
 AOI22_X4 _55967_ (.A1(_23467_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1738]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1689]),
    .B2(_22105_),
    .ZN(_24751_));
 NAND3_X1 _55968_ (.A1(_23296_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1787]),
    .A3(_23294_),
    .ZN(_24752_));
 NAND3_X1 _55969_ (.A1(_23455_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1591]),
    .A3(_23398_),
    .ZN(_24753_));
 AND4_X4 _55970_ (.A1(_24750_),
    .A2(_24751_),
    .A3(_24752_),
    .A4(_24753_),
    .ZN(_24754_));
 AND3_X1 _55971_ (.A1(_23168_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2620]),
    .A3(_23669_),
    .ZN(_24755_));
 AOI221_X4 _55972_ (.A(_24755_),
    .B1(_23374_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2669]),
    .C1(_23373_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2718]),
    .ZN(_24756_));
 NAND3_X1 _55973_ (.A1(_22967_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2375]),
    .A3(_23013_),
    .ZN(_24757_));
 OAI21_X1 _55974_ (.A(_24757_),
    .B1(_10923_),
    .B2(_21756_),
    .ZN(_24758_));
 AND3_X1 _55975_ (.A1(_22954_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2522]),
    .A3(_23013_),
    .ZN(_24759_));
 AND3_X1 _55976_ (.A1(_10843_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2571]),
    .A3(_10891_),
    .ZN(_24760_));
 AND3_X1 _55977_ (.A1(_22522_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2473]),
    .A3(_10891_),
    .ZN(_24761_));
 NOR4_X2 _55978_ (.A1(_24758_),
    .A2(_24759_),
    .A3(_24760_),
    .A4(_24761_),
    .ZN(_24762_));
 AND4_X4 _55979_ (.A1(_24749_),
    .A2(_24754_),
    .A3(_24756_),
    .A4(_24762_),
    .ZN(_24763_));
 NAND4_X1 _55980_ (.A1(_24717_),
    .A2(_24731_),
    .A3(_24747_),
    .A4(_24763_),
    .ZN(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [23]));
 AND3_X1 _55981_ (.A1(_22953_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2915]),
    .A3(_10788_),
    .ZN(_24764_));
 AOI221_X4 _55982_ (.A(_24764_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2866]),
    .B2(_21502_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2817]),
    .C2(_21536_),
    .ZN(_24765_));
 NAND3_X1 _55983_ (.A1(_23217_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1935]),
    .A3(_23402_),
    .ZN(_24766_));
 OAI221_X2 _55984_ (.A(_24766_),
    .B1(_22057_),
    .B2(_10998_),
    .C1(_10994_),
    .C2(_22027_),
    .ZN(_24767_));
 AOI221_X2 _55985_ (.A(_24767_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1788]),
    .B2(_11002_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1641]),
    .C2(_23604_),
    .ZN(_24768_));
 NAND3_X1 _55986_ (.A1(_23245_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3111]),
    .A3(_23360_),
    .ZN(_24769_));
 NAND3_X1 _55987_ (.A1(_23240_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3062]),
    .A3(_22990_),
    .ZN(_24770_));
 NAND2_X2 _55988_ (.A1(_24769_),
    .A2(_24770_),
    .ZN(_24771_));
 AND3_X1 _55989_ (.A1(_22932_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2964]),
    .A3(_10789_),
    .ZN(_24772_));
 AND3_X1 _55990_ (.A1(_23084_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2768]),
    .A3(_10789_),
    .ZN(_24773_));
 AND3_X1 _55991_ (.A1(_10830_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3013]),
    .A3(_10789_),
    .ZN(_24774_));
 NOR4_X4 _55992_ (.A1(_24771_),
    .A2(_24772_),
    .A3(_24773_),
    .A4(_24774_),
    .ZN(_24775_));
 NAND3_X1 _55993_ (.A1(_10868_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2033]),
    .A3(_23600_),
    .ZN(_24776_));
 AOI22_X2 _55994_ (.A1(_23097_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2327]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2278]),
    .B2(_21816_),
    .ZN(_24777_));
 NAND3_X1 _55995_ (.A1(_23367_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2180]),
    .A3(_23553_),
    .ZN(_24778_));
 NAND3_X1 _55996_ (.A1(_23252_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2229]),
    .A3(_23553_),
    .ZN(_24779_));
 AND4_X4 _55997_ (.A1(_24776_),
    .A2(_24777_),
    .A3(_24778_),
    .A4(_24779_),
    .ZN(_24780_));
 AND4_X1 _55998_ (.A1(_24765_),
    .A2(net25),
    .A3(net10),
    .A4(_24780_),
    .ZN(_24781_));
 AND3_X1 _55999_ (.A1(_10816_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [710]),
    .A3(_11124_),
    .ZN(_24782_));
 AOI221_X2 _56000_ (.A(_24782_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [661]),
    .B2(_22642_),
    .C1(_22597_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [759]),
    .ZN(_24783_));
 OAI221_X2 _56001_ (.A(_24783_),
    .B1(_22679_),
    .B2(_11142_),
    .C1(_22743_),
    .C2(_11165_),
    .ZN(_24784_));
 NAND3_X1 _56002_ (.A1(_23560_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [367]),
    .A3(_22951_),
    .ZN(_24785_));
 OAI221_X2 _56003_ (.A(_24785_),
    .B1(_22789_),
    .B2(_11187_),
    .C1(_11182_),
    .C2(_22770_),
    .ZN(_24786_));
 NAND3_X1 _56004_ (.A1(_22933_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [220]),
    .A3(_23341_),
    .ZN(_24787_));
 NAND3_X1 _56005_ (.A1(_23377_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [73]),
    .A3(_22940_),
    .ZN(_24788_));
 NAND2_X2 _56006_ (.A1(_24787_),
    .A2(_24788_),
    .ZN(_24789_));
 AND3_X1 _56007_ (.A1(_10779_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [563]),
    .A3(_11125_),
    .ZN(_24790_));
 AOI21_X4 _56008_ (.A(_24790_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [514]),
    .B2(_11153_),
    .ZN(_24791_));
 NAND3_X4 _56009_ (.A1(_23189_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [465]),
    .A3(_23201_),
    .ZN(_24792_));
 NAND3_X4 _56010_ (.A1(_23837_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [24]),
    .A3(_22959_),
    .ZN(_24793_));
 AOI22_X4 _56011_ (.A1(_11196_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [171]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [122]),
    .B2(_22827_),
    .ZN(_24794_));
 NAND4_X2 _56012_ (.A1(_24791_),
    .A2(_24792_),
    .A3(_24793_),
    .A4(_24794_),
    .ZN(_24795_));
 NOR4_X4 _56013_ (.A1(net47),
    .A2(_24786_),
    .A3(_24789_),
    .A4(_24795_),
    .ZN(_24796_));
 AOI22_X2 _56014_ (.A1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1396]),
    .A2(_23094_),
    .B1(_23325_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1200]),
    .ZN(_24797_));
 AOI22_X4 _56015_ (.A1(_23315_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1543]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1494]),
    .B2(_23095_),
    .ZN(_24798_));
 OAI211_X4 _56016_ (.A(_24797_),
    .B(_24798_),
    .C1(_22245_),
    .C2(_11046_),
    .ZN(_24799_));
 NAND3_X4 _56017_ (.A1(_24050_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1102]),
    .A3(_23882_),
    .ZN(_24800_));
 OAI221_X2 _56018_ (.A(_24800_),
    .B1(_11096_),
    .B2(_22474_),
    .C1(_11076_),
    .C2(_22401_),
    .ZN(_24801_));
 NAND3_X2 _56019_ (.A1(_23145_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1249]),
    .A3(_23277_),
    .ZN(_24802_));
 OAI221_X2 _56020_ (.A(_24802_),
    .B1(_11061_),
    .B2(_22324_),
    .C1(_11055_),
    .C2(_22300_),
    .ZN(_24803_));
 AOI22_X4 _56021_ (.A1(_23267_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [808]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [857]),
    .B2(_23268_),
    .ZN(_24804_));
 NAND3_X2 _56022_ (.A1(_23078_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [906]),
    .A3(_22976_),
    .ZN(_24805_));
 NAND3_X2 _56023_ (.A1(_23080_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1053]),
    .A3(_23547_),
    .ZN(_24806_));
 NAND3_X2 _56024_ (.A1(_23421_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [955]),
    .A3(_23317_),
    .ZN(_24807_));
 NAND4_X4 _56025_ (.A1(_24804_),
    .A2(_24805_),
    .A3(_24806_),
    .A4(_24807_),
    .ZN(_24808_));
 NOR4_X4 _56026_ (.A1(_24799_),
    .A2(_24801_),
    .A3(_24803_),
    .A4(_24808_),
    .ZN(_24809_));
 AND3_X1 _56027_ (.A1(_10856_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1690]),
    .A3(_22923_),
    .ZN(_24810_));
 AOI221_X4 _56028_ (.A(_24810_),
    .B1(_11025_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1592]),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1739]),
    .C2(_22078_),
    .ZN(_24811_));
 NAND3_X1 _56029_ (.A1(_23113_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2425]),
    .A3(_10892_),
    .ZN(_24812_));
 AOI22_X4 _56030_ (.A1(_23587_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2523]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2474]),
    .B2(_21705_),
    .ZN(_24813_));
 NAND3_X1 _56031_ (.A1(_23455_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2376]),
    .A3(_23119_),
    .ZN(_24814_));
 NAND3_X1 _56032_ (.A1(_23757_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2621]),
    .A3(_23119_),
    .ZN(_24815_));
 AND4_X1 _56033_ (.A1(_24812_),
    .A2(_24813_),
    .A3(_24814_),
    .A4(_24815_),
    .ZN(_24816_));
 AND3_X1 _56034_ (.A1(_22521_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2082]),
    .A3(_23169_),
    .ZN(_24817_));
 AOI221_X4 _56035_ (.A(_24817_),
    .B1(_10976_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1984]),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2131]),
    .C2(_23736_),
    .ZN(_24818_));
 AND3_X1 _56036_ (.A1(_23309_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2572]),
    .A3(_23310_),
    .ZN(_24819_));
 AOI221_X4 _56037_ (.A(_24819_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2670]),
    .B2(_21600_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2719]),
    .C2(_21573_),
    .ZN(_24820_));
 AND4_X4 _56038_ (.A1(_24811_),
    .A2(_24816_),
    .A3(_24818_),
    .A4(_24820_),
    .ZN(_24821_));
 NAND4_X4 _56039_ (.A1(_24781_),
    .A2(net9),
    .A3(net3),
    .A4(_24821_),
    .ZN(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [24]));
 NAND3_X1 _56040_ (.A1(_23438_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1054]),
    .A3(_23317_),
    .ZN(_24822_));
 AND3_X1 _56041_ (.A1(_22896_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1152]),
    .A3(_11079_),
    .ZN(_24823_));
 AOI221_X2 _56042_ (.A(_24823_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1103]),
    .B2(_11085_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1005]),
    .C2(_11094_),
    .ZN(_24824_));
 AND3_X2 _56043_ (.A1(_10855_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [907]),
    .A3(_11089_),
    .ZN(_24825_));
 AOI221_X2 _56044_ (.A(_24825_),
    .B1(_11114_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [809]),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [956]),
    .C2(_11099_),
    .ZN(_24826_));
 NAND3_X1 _56045_ (.A1(_10868_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [858]),
    .A3(_23329_),
    .ZN(_24827_));
 AND4_X4 _56046_ (.A1(_24822_),
    .A2(_24824_),
    .A3(_24826_),
    .A4(_24827_),
    .ZN(_24828_));
 AND3_X1 _56047_ (.A1(_22907_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [417]),
    .A3(_23151_),
    .ZN(_24829_));
 AOI221_X4 _56048_ (.A(_24829_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [515]),
    .B2(_23689_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [564]),
    .C2(_11147_),
    .ZN(_24830_));
 AND3_X1 _56049_ (.A1(_10829_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [662]),
    .A3(_23512_),
    .ZN(_24831_));
 AOI221_X4 _56050_ (.A(_24831_),
    .B1(_11131_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [711]),
    .C1(_23638_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [760]),
    .ZN(_24832_));
 AOI22_X2 _56051_ (.A1(_23106_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [613]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [466]),
    .B2(_11159_),
    .ZN(_24833_));
 AND4_X4 _56052_ (.A1(_24828_),
    .A2(_24830_),
    .A3(_24832_),
    .A4(_24833_),
    .ZN(_24834_));
 AOI22_X2 _56053_ (.A1(_23224_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3112]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3063]),
    .B2(_10813_),
    .ZN(_24835_));
 NAND3_X1 _56054_ (.A1(_23221_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2965]),
    .A3(_23431_),
    .ZN(_24836_));
 NAND3_X1 _56055_ (.A1(_23434_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3014]),
    .A3(_23673_),
    .ZN(_24837_));
 AND3_X2 _56056_ (.A1(_24835_),
    .A2(_24836_),
    .A3(_24837_),
    .ZN(_24838_));
 OAI22_X2 _56057_ (.A1(_10875_),
    .A2(_21321_),
    .B1(_21553_),
    .B2(_10864_),
    .ZN(_24839_));
 AOI221_X2 _56058_ (.A(_24839_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2916]),
    .B2(_21466_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2867]),
    .C2(_21502_),
    .ZN(_24840_));
 OAI22_X1 _56059_ (.A1(_10977_),
    .A2(_21975_),
    .B1(_21950_),
    .B2(_10973_),
    .ZN(_24841_));
 AOI221_X4 _56060_ (.A(_24841_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2132]),
    .B2(_10961_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2083]),
    .C2(_21900_),
    .ZN(_24842_));
 NAND3_X1 _56061_ (.A1(_22241_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2230]),
    .A3(_10941_),
    .ZN(_24843_));
 NAND3_X1 _56062_ (.A1(_23390_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2328]),
    .A3(_23388_),
    .ZN(_24844_));
 NAND3_X1 _56063_ (.A1(_23296_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2181]),
    .A3(_23388_),
    .ZN(_24845_));
 NAND3_X1 _56064_ (.A1(_10818_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2279]),
    .A3(_23005_),
    .ZN(_24846_));
 AND4_X4 _56065_ (.A1(_24843_),
    .A2(_24844_),
    .A3(_24845_),
    .A4(_24846_),
    .ZN(_24847_));
 AND4_X4 _56066_ (.A1(_24838_),
    .A2(_24840_),
    .A3(_24842_),
    .A4(_24847_),
    .ZN(_24848_));
 AND3_X1 _56067_ (.A1(_23284_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [368]),
    .A3(_11174_),
    .ZN(_24849_));
 AOI221_X2 _56068_ (.A(_24849_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [319]),
    .B2(_11181_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [270]),
    .C2(_23446_),
    .ZN(_24850_));
 NAND3_X1 _56069_ (.A1(_22993_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [25]),
    .A3(_23246_),
    .ZN(_24851_));
 AOI22_X4 _56070_ (.A1(_22806_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [172]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [123]),
    .B2(_23453_),
    .ZN(_24852_));
 NAND3_X1 _56071_ (.A1(_23367_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [221]),
    .A3(_22939_),
    .ZN(_24853_));
 NAND3_X1 _56072_ (.A1(_23293_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [74]),
    .A3(_22939_),
    .ZN(_24854_));
 AND4_X4 _56073_ (.A1(_24851_),
    .A2(_24852_),
    .A3(_24853_),
    .A4(_24854_),
    .ZN(_24855_));
 NAND3_X1 _56074_ (.A1(_23113_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1250]),
    .A3(_23050_),
    .ZN(_24856_));
 AOI22_X2 _56075_ (.A1(_22282_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1348]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1299]),
    .B2(_11060_),
    .ZN(_24857_));
 NAND3_X1 _56076_ (.A1(_23455_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1201]),
    .A3(_23608_),
    .ZN(_24858_));
 NAND3_X1 _56077_ (.A1(_23303_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1446]),
    .A3(_23608_),
    .ZN(_24859_));
 AND4_X4 _56078_ (.A1(_24856_),
    .A2(_24857_),
    .A3(_24858_),
    .A4(_24859_),
    .ZN(_24860_));
 AND3_X1 _56079_ (.A1(_23309_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1397]),
    .A3(_22979_),
    .ZN(_24861_));
 AOI221_X4 _56080_ (.A(_24861_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1495]),
    .B2(_22210_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1544]),
    .C2(_23179_),
    .ZN(_24862_));
 AND4_X4 _56081_ (.A1(_24850_),
    .A2(_24855_),
    .A3(_24860_),
    .A4(_24862_),
    .ZN(_24863_));
 AND3_X1 _56082_ (.A1(_23751_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1887]),
    .A3(_23519_),
    .ZN(_24864_));
 AOI221_X4 _56083_ (.A(_24864_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1838]),
    .B2(_22044_),
    .C1(_23584_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1936]),
    .ZN(_24865_));
 AOI22_X1 _56084_ (.A1(_23290_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1740]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1691]),
    .B2(_23591_),
    .ZN(_24866_));
 NAND3_X1 _56085_ (.A1(_23328_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1789]),
    .A3(_23576_),
    .ZN(_24867_));
 AOI22_X2 _56086_ (.A1(_23595_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1593]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1642]),
    .B2(_23396_),
    .ZN(_24868_));
 AND3_X4 _56087_ (.A1(_24866_),
    .A2(_24867_),
    .A3(_24868_),
    .ZN(_24869_));
 NAND3_X1 _56088_ (.A1(_22987_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2524]),
    .A3(_10892_),
    .ZN(_24870_));
 AOI22_X1 _56089_ (.A1(_23300_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2377]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2426]),
    .B2(_23301_),
    .ZN(_24871_));
 NAND3_X1 _56090_ (.A1(_23306_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2475]),
    .A3(_23304_),
    .ZN(_24872_));
 NAND3_X1 _56091_ (.A1(_23303_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2622]),
    .A3(_23304_),
    .ZN(_24873_));
 AND4_X2 _56092_ (.A1(_24870_),
    .A2(_24871_),
    .A3(_24872_),
    .A4(_24873_),
    .ZN(_24874_));
 AND3_X1 _56093_ (.A1(_23217_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2720]),
    .A3(_23310_),
    .ZN(_24875_));
 AOI221_X2 _56094_ (.A(_24875_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2671]),
    .B2(_21600_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2573]),
    .C2(_21654_),
    .ZN(_24876_));
 AND4_X4 _56095_ (.A1(_24865_),
    .A2(_24869_),
    .A3(_24874_),
    .A4(_24876_),
    .ZN(_24877_));
 NAND4_X2 _56096_ (.A1(_24834_),
    .A2(_24848_),
    .A3(_24863_),
    .A4(_24877_),
    .ZN(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [25]));
 NAND3_X1 _56097_ (.A1(_23438_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3015]),
    .A3(_23431_),
    .ZN(_24878_));
 AOI22_X2 _56098_ (.A1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2770]),
    .A2(_23625_),
    .B1(_10839_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2966]),
    .ZN(_24879_));
 NAND3_X1 _56099_ (.A1(_24186_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3064]),
    .A3(_23222_),
    .ZN(_24880_));
 NAND3_X1 _56100_ (.A1(_23245_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3113]),
    .A3(_23222_),
    .ZN(_24881_));
 AND4_X4 _56101_ (.A1(_24878_),
    .A2(_24879_),
    .A3(_24880_),
    .A4(_24881_),
    .ZN(_24882_));
 NAND3_X1 _56102_ (.A1(_23408_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1496]),
    .A3(_22979_),
    .ZN(_24883_));
 OAI221_X2 _56103_ (.A(_24883_),
    .B1(_22247_),
    .B2(_11046_),
    .C1(_11032_),
    .C2(_22204_),
    .ZN(_24884_));
 AOI221_X2 _56104_ (.A(_24884_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1398]),
    .B2(_23094_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1202]),
    .C2(_23103_),
    .ZN(_24885_));
 AND3_X1 _56105_ (.A1(_10842_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2574]),
    .A3(_10886_),
    .ZN(_24886_));
 AOI221_X4 _56106_ (.A(_24886_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2672]),
    .B2(_21600_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2721]),
    .C2(_10887_),
    .ZN(_24887_));
 AND3_X1 _56107_ (.A1(_10855_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2476]),
    .A3(_10886_),
    .ZN(_24888_));
 AOI221_X2 _56108_ (.A(_24888_),
    .B1(_10928_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2378]),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2525]),
    .C2(_10911_),
    .ZN(_24889_));
 AOI22_X2 _56109_ (.A1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2623]),
    .A2(_23627_),
    .B1(_23301_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2427]),
    .ZN(_24890_));
 AND3_X1 _56110_ (.A1(_10854_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2868]),
    .A3(net106),
    .ZN(_24891_));
 AOI221_X2 _56111_ (.A(_24891_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2819]),
    .B2(_10863_),
    .C1(_10773_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2917]),
    .ZN(_24892_));
 AND4_X4 _56112_ (.A1(_24887_),
    .A2(_24889_),
    .A3(_24890_),
    .A4(_24892_),
    .ZN(_24893_));
 AND3_X1 _56113_ (.A1(_10797_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1153]),
    .A3(_11089_),
    .ZN(_24894_));
 AOI221_X2 _56114_ (.A(_24894_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1104]),
    .B2(_11085_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1006]),
    .C2(_11094_),
    .ZN(_24895_));
 AOI22_X2 _56115_ (.A1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1055]),
    .A2(_23632_),
    .B1(_22544_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [859]),
    .ZN(_24896_));
 AND3_X1 _56116_ (.A1(_10873_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [810]),
    .A3(_11089_),
    .ZN(_24897_));
 AOI221_X4 _56117_ (.A(_24897_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [908]),
    .B2(_11105_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [957]),
    .C2(_11099_),
    .ZN(_24898_));
 AND3_X1 _56118_ (.A1(_10920_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1251]),
    .A3(_11034_),
    .ZN(_24899_));
 AOI221_X2 _56119_ (.A(_24899_),
    .B1(_11059_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1300]),
    .C1(_11054_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1349]),
    .ZN(_24900_));
 AND4_X4 _56120_ (.A1(_24895_),
    .A2(_24896_),
    .A3(_24898_),
    .A4(_24900_),
    .ZN(_24901_));
 AND4_X4 _56121_ (.A1(_24882_),
    .A2(net24),
    .A3(_24893_),
    .A4(_24901_),
    .ZN(_24902_));
 NAND3_X1 _56122_ (.A1(_10880_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [26]),
    .A3(_23341_),
    .ZN(_24903_));
 AND3_X1 _56123_ (.A1(_23751_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [320]),
    .A3(_23159_),
    .ZN(_24904_));
 AOI221_X4 _56124_ (.A(_24904_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [271]),
    .B2(_22777_),
    .C1(_23615_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [369]),
    .ZN(_24905_));
 AOI22_X1 _56125_ (.A1(_11196_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [173]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [124]),
    .B2(_22827_),
    .ZN(_24906_));
 AOI22_X1 _56126_ (.A1(_23248_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [222]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [75]),
    .B2(_23490_),
    .ZN(_24907_));
 AND4_X2 _56127_ (.A1(_24903_),
    .A2(_24905_),
    .A3(_24906_),
    .A4(_24907_),
    .ZN(_24908_));
 NAND3_X2 _56128_ (.A1(_22242_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [663]),
    .A3(_11127_),
    .ZN(_24909_));
 AND3_X1 _56129_ (.A1(_23524_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [712]),
    .A3(_23255_),
    .ZN(_24910_));
 AOI221_X4 _56130_ (.A(_24910_),
    .B1(_23515_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [614]),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [761]),
    .C2(_22597_),
    .ZN(_24911_));
 AOI22_X2 _56131_ (.A1(_23622_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [565]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [516]),
    .B2(_11153_),
    .ZN(_24912_));
 AOI22_X2 _56132_ (.A1(_23610_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [418]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [467]),
    .B2(_11159_),
    .ZN(_24913_));
 AND4_X4 _56133_ (.A1(_24909_),
    .A2(_24911_),
    .A3(_24912_),
    .A4(_24913_),
    .ZN(_24914_));
 AND3_X1 _56134_ (.A1(_23382_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1986]),
    .A3(_23231_),
    .ZN(_24915_));
 AOI221_X4 _56135_ (.A(_24915_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2084]),
    .B2(_23233_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2133]),
    .C2(_10962_),
    .ZN(_24916_));
 OAI22_X2 _56136_ (.A1(_11026_),
    .A2(_22172_),
    .B1(_22148_),
    .B2(_11020_),
    .ZN(_24917_));
 OAI22_X2 _56137_ (.A1(_11009_),
    .A2(_22094_),
    .B1(_22124_),
    .B2(_11013_),
    .ZN(_24918_));
 AOI211_X2 _56138_ (.A(_24917_),
    .B(_24918_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1790]),
    .C2(_11003_),
    .ZN(_24919_));
 NAND3_X1 _56139_ (.A1(_22997_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2231]),
    .A3(_23553_),
    .ZN(_24920_));
 AOI22_X2 _56140_ (.A1(_23660_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2182]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2035]),
    .B2(_21937_),
    .ZN(_24921_));
 NAND3_X1 _56141_ (.A1(_10818_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2280]),
    .A3(_23005_),
    .ZN(_24922_));
 NAND3_X1 _56142_ (.A1(_22949_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2329]),
    .A3(_23005_),
    .ZN(_24923_));
 AND4_X4 _56143_ (.A1(_24920_),
    .A2(_24921_),
    .A3(_24922_),
    .A4(_24923_),
    .ZN(_24924_));
 AND3_X1 _56144_ (.A1(_23215_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1839]),
    .A3(_23402_),
    .ZN(_24925_));
 AOI221_X4 _56145_ (.A(_24925_),
    .B1(_10993_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1888]),
    .C1(_21978_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1937]),
    .ZN(_24926_));
 AND4_X4 _56146_ (.A1(_24916_),
    .A2(_24919_),
    .A3(_24924_),
    .A4(_24926_),
    .ZN(_24927_));
 NAND4_X4 _56147_ (.A1(_24902_),
    .A2(_24908_),
    .A3(_24914_),
    .A4(_24927_),
    .ZN(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [26]));
 OAI22_X2 _56148_ (.A1(_10774_),
    .A2(_21488_),
    .B1(_21523_),
    .B2(_10852_),
    .ZN(_24928_));
 AOI221_X2 _56149_ (.A(_24928_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2771]),
    .B2(_10874_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2820]),
    .C2(_21536_),
    .ZN(_24929_));
 NAND3_X2 _56150_ (.A1(_23340_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2967]),
    .A3(_23361_),
    .ZN(_24930_));
 AND3_X1 _56151_ (.A1(_10816_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3065]),
    .A3(_10825_),
    .ZN(_24931_));
 AOI221_X2 _56152_ (.A(_24931_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3016]),
    .B2(_10826_),
    .C1(_10799_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3114]),
    .ZN(_24932_));
 AND3_X1 _56153_ (.A1(_22521_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2477]),
    .A3(_23310_),
    .ZN(_24933_));
 AOI221_X4 _56154_ (.A(_24933_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2428]),
    .B2(_10921_),
    .C1(_10912_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2526]),
    .ZN(_24934_));
 NAND4_X4 _56155_ (.A1(_24929_),
    .A2(_24930_),
    .A3(_24932_),
    .A4(_24934_),
    .ZN(_24935_));
 AND3_X1 _56156_ (.A1(_10824_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1840]),
    .A3(_10987_),
    .ZN(_24936_));
 AOI221_X4 _56157_ (.A(_24936_),
    .B1(_10993_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1889]),
    .C1(_21978_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1938]),
    .ZN(_24937_));
 NAND3_X4 _56158_ (.A1(_22933_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1791]),
    .A3(_23116_),
    .ZN(_24938_));
 AOI22_X4 _56159_ (.A1(_23290_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1742]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1693]),
    .B2(_23591_),
    .ZN(_24939_));
 AOI22_X2 _56160_ (.A1(_23595_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1595]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1644]),
    .B2(_23604_),
    .ZN(_24940_));
 NAND4_X4 _56161_ (.A1(_24937_),
    .A2(_24938_),
    .A3(_24939_),
    .A4(_24940_),
    .ZN(_24941_));
 AND3_X1 _56162_ (.A1(_10866_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [468]),
    .A3(_11124_),
    .ZN(_24942_));
 AOI221_X4 _56163_ (.A(_24942_),
    .B1(_11152_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [517]),
    .C1(_11146_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [566]),
    .ZN(_24943_));
 AND3_X1 _56164_ (.A1(_23084_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [419]),
    .A3(_11125_),
    .ZN(_24944_));
 AOI21_X2 _56165_ (.A(_24944_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [615]),
    .B2(_23106_),
    .ZN(_24945_));
 NAND3_X4 _56166_ (.A1(_23536_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [664]),
    .A3(_23060_),
    .ZN(_24946_));
 AOI22_X4 _56167_ (.A1(_23638_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [762]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [713]),
    .B2(_23092_),
    .ZN(_24947_));
 NAND4_X4 _56168_ (.A1(_24943_),
    .A2(_24945_),
    .A3(_24946_),
    .A4(_24947_),
    .ZN(_24948_));
 AND3_X1 _56169_ (.A1(_10798_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1154]),
    .A3(_11079_),
    .ZN(_24949_));
 AOI221_X2 _56170_ (.A(_24949_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1105]),
    .B2(_11085_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1056]),
    .C2(_11090_),
    .ZN(_24950_));
 OAI221_X2 _56171_ (.A(net46),
    .B1(_22476_),
    .B2(_11096_),
    .C1(_22587_),
    .C2(_11115_),
    .ZN(_24951_));
 NOR4_X2 _56172_ (.A1(_24935_),
    .A2(_24941_),
    .A3(_24948_),
    .A4(net23),
    .ZN(_24952_));
 AND3_X1 _56173_ (.A1(_10824_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2624]),
    .A3(_23310_),
    .ZN(_24953_));
 AOI221_X2 _56174_ (.A(_24953_),
    .B1(_21601_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2673]),
    .C1(_21573_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2722]),
    .ZN(_24954_));
 NAND3_X2 _56175_ (.A1(_23368_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2575]),
    .A3(_10893_),
    .ZN(_24955_));
 OAI211_X4 _56176_ (.A(net45),
    .B(_24955_),
    .C1(_21785_),
    .C2(_10930_),
    .ZN(_24956_));
 NAND3_X2 _56177_ (.A1(_23377_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2036]),
    .A3(_23561_),
    .ZN(_24957_));
 OAI221_X2 _56178_ (.A(_24957_),
    .B1(_10969_),
    .B2(_21921_),
    .C1(_10963_),
    .C2(_21894_),
    .ZN(_24958_));
 NAND3_X1 _56179_ (.A1(_23076_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2330]),
    .A3(_24052_),
    .ZN(_24959_));
 NAND3_X1 _56180_ (.A1(_23888_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2281]),
    .A3(_23894_),
    .ZN(_24960_));
 OAI211_X2 _56181_ (.A(_24959_),
    .B(_24960_),
    .C1(_21859_),
    .C2(_10951_),
    .ZN(_24961_));
 NAND3_X2 _56182_ (.A1(_23008_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1987]),
    .A3(_24046_),
    .ZN(_24962_));
 OAI21_X4 _56183_ (.A(_24962_),
    .B1(_10957_),
    .B2(_21874_),
    .ZN(_24963_));
 NOR4_X4 _56184_ (.A1(_24956_),
    .A2(_24958_),
    .A3(_24961_),
    .A4(_24963_),
    .ZN(_24964_));
 NAND3_X2 _56185_ (.A1(_23340_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [223]),
    .A3(_23341_),
    .ZN(_24965_));
 AND3_X1 _56186_ (.A1(_23524_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [321]),
    .A3(_23258_),
    .ZN(_24966_));
 AOI221_X4 _56187_ (.A(_24966_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [272]),
    .B2(_22777_),
    .C1(_23615_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [370]),
    .ZN(_24967_));
 AOI22_X2 _56188_ (.A1(_11196_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [174]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [125]),
    .B2(_22827_),
    .ZN(_24968_));
 AOI22_X2 _56189_ (.A1(_11206_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [27]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [76]),
    .B2(_23490_),
    .ZN(_24969_));
 AND4_X4 _56190_ (.A1(_24965_),
    .A2(_24967_),
    .A3(_24968_),
    .A4(_24969_),
    .ZN(_24970_));
 NAND3_X1 _56191_ (.A1(_23340_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1399]),
    .A3(_23051_),
    .ZN(_24971_));
 NAND3_X1 _56192_ (.A1(_23083_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1203]),
    .A3(_22979_),
    .ZN(_24972_));
 OAI21_X1 _56193_ (.A(_24972_),
    .B1(_11066_),
    .B2(_22347_),
    .ZN(_24973_));
 AOI221_X4 _56194_ (.A(_24973_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1350]),
    .B2(_23748_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1301]),
    .C2(_23262_),
    .ZN(_24974_));
 AND3_X1 _56195_ (.A1(_23459_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1546]),
    .A3(_23701_),
    .ZN(_24975_));
 AOI221_X4 _56196_ (.A(_24975_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1497]),
    .B2(_22210_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1448]),
    .C2(_22232_),
    .ZN(_24976_));
 AND3_X1 _56197_ (.A1(_10778_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [958]),
    .A3(_23938_),
    .ZN(_24977_));
 AOI221_X4 _56198_ (.A(_24977_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [909]),
    .B2(_11106_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [860]),
    .C2(_22544_),
    .ZN(_24978_));
 AND4_X4 _56199_ (.A1(_24971_),
    .A2(_24974_),
    .A3(_24976_),
    .A4(_24978_),
    .ZN(_24979_));
 NAND4_X4 _56200_ (.A1(_24952_),
    .A2(net8),
    .A3(_24970_),
    .A4(_24979_),
    .ZN(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [27]));
 AND3_X1 _56201_ (.A1(_23721_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [518]),
    .A3(_23504_),
    .ZN(_24980_));
 AOI221_X4 _56202_ (.A(_24980_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [469]),
    .B2(_11158_),
    .C1(_23622_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [567]),
    .ZN(_24981_));
 NAND3_X2 _56203_ (.A1(_23217_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [763]),
    .A3(_11124_),
    .ZN(_24982_));
 OAI221_X2 _56204_ (.A(_24982_),
    .B1(_22656_),
    .B2(_11137_),
    .C1(_11132_),
    .C2(_22636_),
    .ZN(_24983_));
 AOI221_X2 _56205_ (.A(_24983_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [616]),
    .B2(_23515_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [420]),
    .C2(_23610_),
    .ZN(_24984_));
 AND3_X1 _56206_ (.A1(_23284_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [371]),
    .A3(_11174_),
    .ZN(_24985_));
 AOI221_X2 _56207_ (.A(_24985_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [322]),
    .B2(_11181_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [273]),
    .C2(_23446_),
    .ZN(_24986_));
 NAND3_X1 _56208_ (.A1(_23982_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [126]),
    .A3(_23246_),
    .ZN(_24987_));
 AOI22_X1 _56209_ (.A1(_23164_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [28]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [77]),
    .B2(_23714_),
    .ZN(_24988_));
 NAND3_X1 _56210_ (.A1(_23367_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [224]),
    .A3(_23451_),
    .ZN(_24989_));
 NAND3_X1 _56211_ (.A1(_23003_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [175]),
    .A3(_23250_),
    .ZN(_24990_));
 AND4_X1 _56212_ (.A1(_24987_),
    .A2(_24988_),
    .A3(_24989_),
    .A4(_24990_),
    .ZN(_24991_));
 AND4_X4 _56213_ (.A1(_24981_),
    .A2(net22),
    .A3(_24986_),
    .A4(_24991_),
    .ZN(_24992_));
 NAND3_X2 _56214_ (.A1(_22988_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2135]),
    .A3(_23554_),
    .ZN(_24993_));
 OAI221_X2 _56215_ (.A(_24993_),
    .B1(_21954_),
    .B2(_10973_),
    .C1(_10969_),
    .C2(_21923_),
    .ZN(_24994_));
 NAND3_X1 _56216_ (.A1(_23367_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2184]),
    .A3(_23388_),
    .ZN(_24995_));
 NAND3_X1 _56217_ (.A1(_23455_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1988]),
    .A3(_23388_),
    .ZN(_24996_));
 AND2_X2 _56218_ (.A1(_24995_),
    .A2(_24996_),
    .ZN(_24997_));
 NAND3_X2 _56219_ (.A1(_10831_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2233]),
    .A3(_23006_),
    .ZN(_24998_));
 NAND3_X1 _56220_ (.A1(_22944_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2282]),
    .A3(_23561_),
    .ZN(_24999_));
 NAND3_X2 _56221_ (.A1(_23560_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2331]),
    .A3(_23561_),
    .ZN(_25000_));
 NAND4_X4 _56222_ (.A1(_24997_),
    .A2(_24998_),
    .A3(_24999_),
    .A4(_25000_),
    .ZN(_25001_));
 OAI22_X4 _56223_ (.A1(_21667_),
    .A2(_10908_),
    .B1(_10930_),
    .B2(_21788_),
    .ZN(_25002_));
 NAND3_X1 _56224_ (.A1(_23236_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2723]),
    .A3(_23026_),
    .ZN(_25003_));
 NAND3_X1 _56225_ (.A1(_22961_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2674]),
    .A3(_23026_),
    .ZN(_25004_));
 OAI211_X2 _56226_ (.A(_25003_),
    .B(_25004_),
    .C1(_21646_),
    .C2(_10903_),
    .ZN(_25005_));
 NOR4_X4 _56227_ (.A1(_24994_),
    .A2(_25001_),
    .A3(_25002_),
    .A4(_25005_),
    .ZN(_25006_));
 AND3_X1 _56228_ (.A1(_10824_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1057]),
    .A3(_23938_),
    .ZN(_25007_));
 AOI221_X2 _56229_ (.A(_25007_),
    .B1(_23332_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1106]),
    .C1(_23331_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1155]),
    .ZN(_25008_));
 NAND3_X2 _56230_ (.A1(_22994_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [812]),
    .A3(_23880_),
    .ZN(_25009_));
 OAI211_X4 _56231_ (.A(_25008_),
    .B(_25009_),
    .C1(_22478_),
    .C2(_11096_),
    .ZN(_25010_));
 AOI22_X4 _56232_ (.A1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1400]),
    .A2(_23094_),
    .B1(_23325_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1204]),
    .ZN(_25011_));
 NAND3_X2 _56233_ (.A1(_22944_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1498]),
    .A3(_24026_),
    .ZN(_25012_));
 NAND3_X1 _56234_ (.A1(_23536_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1449]),
    .A3(_11037_),
    .ZN(_25013_));
 NAND3_X2 _56235_ (.A1(_23067_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1547]),
    .A3(_11037_),
    .ZN(_25014_));
 NAND4_X4 _56236_ (.A1(_25011_),
    .A2(_25012_),
    .A3(_25013_),
    .A4(_25014_),
    .ZN(_25015_));
 NAND3_X4 _56237_ (.A1(_23421_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [959]),
    .A3(_23891_),
    .ZN(_25016_));
 OAI221_X2 _56238_ (.A(_25016_),
    .B1(_22565_),
    .B2(_11111_),
    .C1(_11107_),
    .C2(_22537_),
    .ZN(_25017_));
 NAND3_X1 _56239_ (.A1(_23204_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1302]),
    .A3(_23205_),
    .ZN(_25018_));
 OAI221_X2 _56240_ (.A(_25018_),
    .B1(_22349_),
    .B2(_11066_),
    .C1(_11055_),
    .C2(_22304_),
    .ZN(_25019_));
 NOR4_X4 _56241_ (.A1(_25010_),
    .A2(_25015_),
    .A3(_25017_),
    .A4(_25019_),
    .ZN(_25020_));
 AND3_X1 _56242_ (.A1(_10816_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1890]),
    .A3(_10987_),
    .ZN(_25021_));
 AOI221_X4 _56243_ (.A(_25021_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1841]),
    .B2(_10997_),
    .C1(_21978_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1939]),
    .ZN(_25022_));
 NAND3_X2 _56244_ (.A1(_23368_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1792]),
    .A3(_23116_),
    .ZN(_25023_));
 AOI22_X2 _56245_ (.A1(_23290_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1743]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1694]),
    .B2(_23591_),
    .ZN(_25024_));
 AOI22_X4 _56246_ (.A1(_23595_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1596]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1645]),
    .B2(_23604_),
    .ZN(_25025_));
 NAND4_X4 _56247_ (.A1(_25022_),
    .A2(_25023_),
    .A3(_25024_),
    .A4(_25025_),
    .ZN(_25026_));
 AND3_X1 _56248_ (.A1(_10824_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3017]),
    .A3(_10825_),
    .ZN(_25027_));
 AOI221_X2 _56249_ (.A(_25027_),
    .B1(_10812_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3066]),
    .C1(_10799_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3115]),
    .ZN(_25028_));
 OAI21_X4 _56250_ (.A(_25028_),
    .B1(_21458_),
    .B2(_10840_),
    .ZN(_25029_));
 AOI22_X4 _56251_ (.A1(_23213_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2919]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2870]),
    .B2(_21502_),
    .ZN(_25030_));
 NAND3_X4 _56252_ (.A1(_23036_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2821]),
    .A3(_23037_),
    .ZN(_25031_));
 OAI211_X4 _56253_ (.A(_25030_),
    .B(_25031_),
    .C1(_21325_),
    .C2(_10875_),
    .ZN(_25032_));
 NAND3_X1 _56254_ (.A1(_23426_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2429]),
    .A3(_23422_),
    .ZN(_25033_));
 OAI221_X2 _56255_ (.A(_25033_),
    .B1(_10917_),
    .B2(_21727_),
    .C1(_10913_),
    .C2(_21698_),
    .ZN(_25034_));
 NOR4_X1 _56256_ (.A1(_25026_),
    .A2(_25029_),
    .A3(_25032_),
    .A4(_25034_),
    .ZN(_25035_));
 NAND4_X1 _56257_ (.A1(_24992_),
    .A2(_25006_),
    .A3(net7),
    .A4(_25035_),
    .ZN(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [28]));
 NAND3_X1 _56258_ (.A1(_23221_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1401]),
    .A3(_23931_),
    .ZN(_25036_));
 NAND3_X1 _56259_ (.A1(_24262_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1548]),
    .A3(_23931_),
    .ZN(_25037_));
 NAND3_X1 _56260_ (.A1(_24186_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1499]),
    .A3(_23931_),
    .ZN(_25038_));
 NAND3_X1 _56261_ (.A1(_23385_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1450]),
    .A3(_23412_),
    .ZN(_25039_));
 AND4_X4 _56262_ (.A1(_25036_),
    .A2(_25037_),
    .A3(_25038_),
    .A4(_25039_),
    .ZN(_25040_));
 OAI22_X2 _56263_ (.A1(_11070_),
    .A2(_22377_),
    .B1(_22351_),
    .B2(_11066_),
    .ZN(_25041_));
 AOI221_X4 _56264_ (.A(_25041_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1352]),
    .B2(_23748_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1303]),
    .C2(_23262_),
    .ZN(_25042_));
 AND3_X1 _56265_ (.A1(_10856_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [519]),
    .A3(_23512_),
    .ZN(_25043_));
 AOI221_X4 _56266_ (.A(_25043_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [470]),
    .B2(_11158_),
    .C1(_23622_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [568]),
    .ZN(_25044_));
 NAND3_X1 _56267_ (.A1(_10798_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [764]),
    .A3(_11124_),
    .ZN(_25045_));
 NAND3_X1 _56268_ (.A1(_10816_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [715]),
    .A3(_11124_),
    .ZN(_25046_));
 OAI211_X2 _56269_ (.A(_25045_),
    .B(_25046_),
    .C1(_22658_),
    .C2(_11137_),
    .ZN(_25047_));
 AOI221_X2 _56270_ (.A(_25047_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [617]),
    .B2(_23515_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [421]),
    .C2(_22733_),
    .ZN(_25048_));
 AND4_X4 _56271_ (.A1(_25040_),
    .A2(_25042_),
    .A3(_25044_),
    .A4(_25048_),
    .ZN(_25049_));
 NAND3_X1 _56272_ (.A1(_23236_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3116]),
    .A3(_23431_),
    .ZN(_25050_));
 NAND3_X1 _56273_ (.A1(_23280_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3067]),
    .A3(_23673_),
    .ZN(_25051_));
 NAND3_X1 _56274_ (.A1(_23434_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3018]),
    .A3(_23673_),
    .ZN(_25052_));
 AND3_X2 _56275_ (.A1(_25050_),
    .A2(_25051_),
    .A3(_25052_),
    .ZN(_25053_));
 NAND3_X1 _56276_ (.A1(_22954_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2920]),
    .A3(_22928_),
    .ZN(_25054_));
 OAI21_X2 _56277_ (.A(_25054_),
    .B1(_10852_),
    .B2(_21525_),
    .ZN(_25055_));
 OAI22_X2 _56278_ (.A1(_10875_),
    .A2(_21327_),
    .B1(_21557_),
    .B2(_10864_),
    .ZN(_25056_));
 AOI211_X2 _56279_ (.A(_25055_),
    .B(_25056_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2969]),
    .C2(_10839_),
    .ZN(_25057_));
 AND3_X1 _56280_ (.A1(_23524_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1891]),
    .A3(_23662_),
    .ZN(_25058_));
 AOI221_X4 _56281_ (.A(_25058_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1842]),
    .B2(_22044_),
    .C1(_21978_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1940]),
    .ZN(_25059_));
 NAND3_X1 _56282_ (.A1(_22993_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1597]),
    .A3(_23393_),
    .ZN(_25060_));
 AOI22_X4 _56283_ (.A1(_23467_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1744]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1695]),
    .B2(_22105_),
    .ZN(_25061_));
 NAND3_X1 _56284_ (.A1(_23296_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1793]),
    .A3(_23294_),
    .ZN(_25062_));
 NAND3_X1 _56285_ (.A1(_23035_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1646]),
    .A3(_23398_),
    .ZN(_25063_));
 AND4_X4 _56286_ (.A1(_25060_),
    .A2(_25061_),
    .A3(_25062_),
    .A4(_25063_),
    .ZN(_25064_));
 AND4_X1 _56287_ (.A1(_25053_),
    .A2(_25057_),
    .A3(_25059_),
    .A4(_25064_),
    .ZN(_25065_));
 AOI22_X4 _56288_ (.A1(_23485_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1989]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2038]),
    .B2(_22911_),
    .ZN(_25066_));
 OAI221_X2 _56289_ (.A(_25066_),
    .B1(_21925_),
    .B2(_10969_),
    .C1(_10963_),
    .C2(_21896_),
    .ZN(_25067_));
 AOI22_X2 _56290_ (.A1(_23097_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2332]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2283]),
    .B2(_21816_),
    .ZN(_25068_));
 NAND3_X2 _56291_ (.A1(_23536_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2234]),
    .A3(_24046_),
    .ZN(_25069_));
 OAI211_X4 _56292_ (.A(_25068_),
    .B(_25069_),
    .C1(_21878_),
    .C2(_10957_),
    .ZN(_25070_));
 NAND3_X2 _56293_ (.A1(_23067_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2724]),
    .A3(_23014_),
    .ZN(_25071_));
 NAND3_X2 _56294_ (.A1(_10844_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2577]),
    .A3(_23023_),
    .ZN(_25072_));
 NAND3_X1 _56295_ (.A1(_22975_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2626]),
    .A3(_23026_),
    .ZN(_25073_));
 NAND3_X2 _56296_ (.A1(_23028_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2675]),
    .A3(_23029_),
    .ZN(_25074_));
 NAND4_X4 _56297_ (.A1(_25071_),
    .A2(_25072_),
    .A3(_25073_),
    .A4(_25074_),
    .ZN(_25075_));
 NAND3_X1 _56298_ (.A1(_22955_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2528]),
    .A3(_23134_),
    .ZN(_25076_));
 NAND3_X1 _56299_ (.A1(_23145_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2430]),
    .A3(_23143_),
    .ZN(_25077_));
 NAND3_X1 _56300_ (.A1(_23039_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2479]),
    .A3(_23043_),
    .ZN(_25078_));
 NAND3_X1 _56301_ (.A1(_23085_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2381]),
    .A3(_23422_),
    .ZN(_25079_));
 NAND4_X2 _56302_ (.A1(_25076_),
    .A2(_25077_),
    .A3(_25078_),
    .A4(_25079_),
    .ZN(_25080_));
 NOR4_X4 _56303_ (.A1(_25067_),
    .A2(_25070_),
    .A3(_25075_),
    .A4(_25080_),
    .ZN(_25081_));
 AND3_X1 _56304_ (.A1(_24467_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [274]),
    .A3(_23159_),
    .ZN(_25082_));
 AOI221_X4 _56305_ (.A(_25082_),
    .B1(_22903_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [323]),
    .C1(_23615_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [372]),
    .ZN(_25083_));
 NAND3_X1 _56306_ (.A1(_22523_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [911]),
    .A3(_23321_),
    .ZN(_25084_));
 AOI22_X2 _56307_ (.A1(_23267_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [813]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [862]),
    .B2(_22544_),
    .ZN(_25085_));
 NAND3_X1 _56308_ (.A1(_23003_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [960]),
    .A3(_11081_),
    .ZN(_25086_));
 NAND3_X1 _56309_ (.A1(_23296_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1009]),
    .A3(_23879_),
    .ZN(_25087_));
 AND4_X4 _56310_ (.A1(_25084_),
    .A2(_25085_),
    .A3(_25086_),
    .A4(_25087_),
    .ZN(_25088_));
 NAND3_X1 _56311_ (.A1(_23242_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [225]),
    .A3(_23451_),
    .ZN(_25089_));
 AOI22_X2 _56312_ (.A1(_23164_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [29]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [78]),
    .B2(_11211_),
    .ZN(_25090_));
 NAND3_X1 _56313_ (.A1(_23306_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [127]),
    .A3(_22939_),
    .ZN(_25091_));
 NAND3_X1 _56314_ (.A1(_23019_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [176]),
    .A3(_22939_),
    .ZN(_25092_));
 AND4_X4 _56315_ (.A1(_25089_),
    .A2(_25090_),
    .A3(_25091_),
    .A4(_25092_),
    .ZN(_25093_));
 AND3_X1 _56316_ (.A1(_23217_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1156]),
    .A3(_23938_),
    .ZN(_25094_));
 AOI221_X2 _56317_ (.A(_25094_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1107]),
    .B2(_23332_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1058]),
    .C2(_22435_),
    .ZN(_25095_));
 AND4_X4 _56318_ (.A1(_25083_),
    .A2(_25088_),
    .A3(_25093_),
    .A4(net44),
    .ZN(_25096_));
 NAND4_X4 _56319_ (.A1(_25049_),
    .A2(_25065_),
    .A3(_25081_),
    .A4(_25096_),
    .ZN(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [29]));
 NAND3_X1 _56320_ (.A1(_23438_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3019]),
    .A3(_23431_),
    .ZN(_25097_));
 AOI22_X2 _56321_ (.A1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2774]),
    .A2(_23625_),
    .B1(_22918_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2970]),
    .ZN(_25098_));
 NAND3_X1 _56322_ (.A1(_24262_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3117]),
    .A3(_23222_),
    .ZN(_25099_));
 NAND3_X2 _56323_ (.A1(_24186_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3068]),
    .A3(_23360_),
    .ZN(_25100_));
 AND4_X4 _56324_ (.A1(_25097_),
    .A2(_25098_),
    .A3(_25099_),
    .A4(_25100_),
    .ZN(_25101_));
 NAND3_X1 _56325_ (.A1(_23221_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [618]),
    .A3(_23237_),
    .ZN(_25102_));
 AND3_X1 _56326_ (.A1(_10797_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [765]),
    .A3(_11145_),
    .ZN(_25103_));
 AOI221_X2 _56327_ (.A(_25103_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [716]),
    .B2(_11131_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [667]),
    .C2(_22642_),
    .ZN(_25104_));
 AOI22_X2 _56328_ (.A1(_23622_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [569]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [520]),
    .B2(_23689_),
    .ZN(_25105_));
 AOI22_X2 _56329_ (.A1(_23610_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [422]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [471]),
    .B2(_11158_),
    .ZN(_25106_));
 AND4_X4 _56330_ (.A1(_25102_),
    .A2(_25104_),
    .A3(_25105_),
    .A4(_25106_),
    .ZN(_25107_));
 AND3_X1 _56331_ (.A1(_22896_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2725]),
    .A3(_10886_),
    .ZN(_25108_));
 AOI221_X2 _56332_ (.A(_25108_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2676]),
    .B2(_10896_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2578]),
    .C2(_21654_),
    .ZN(_25109_));
 AOI22_X1 _56333_ (.A1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2627]),
    .A2(_23627_),
    .B1(_23301_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2431]),
    .ZN(_25110_));
 AND3_X1 _56334_ (.A1(_10854_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2480]),
    .A3(_10886_),
    .ZN(_25111_));
 AOI221_X4 _56335_ (.A(_25111_),
    .B1(_10928_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2382]),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2529]),
    .C2(_10911_),
    .ZN(_25112_));
 AND3_X1 _56336_ (.A1(_10920_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2823]),
    .A3(net107),
    .ZN(_25113_));
 AOI221_X2 _56337_ (.A(_25113_),
    .B1(_10851_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2872]),
    .C1(_10773_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2921]),
    .ZN(_25114_));
 AND4_X4 _56338_ (.A1(_25109_),
    .A2(_25110_),
    .A3(_25112_),
    .A4(_25114_),
    .ZN(_25115_));
 NAND3_X1 _56339_ (.A1(_23385_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1451]),
    .A3(_23412_),
    .ZN(_25116_));
 AND3_X1 _56340_ (.A1(_10811_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1500]),
    .A3(_11034_),
    .ZN(_25117_));
 AOI221_X2 _56341_ (.A(_25117_),
    .B1(_11050_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1402]),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1549]),
    .C2(_11031_),
    .ZN(_25118_));
 AOI22_X2 _56342_ (.A1(_22282_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1353]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1304]),
    .B2(_11060_),
    .ZN(_25119_));
 AOI22_X2 _56343_ (.A1(_23103_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1206]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1255]),
    .B2(_23048_),
    .ZN(_25120_));
 AND4_X4 _56344_ (.A1(_25116_),
    .A2(_25118_),
    .A3(_25119_),
    .A4(_25120_),
    .ZN(_25121_));
 AND4_X1 _56345_ (.A1(_25101_),
    .A2(_25107_),
    .A3(_25115_),
    .A4(_25121_),
    .ZN(_25122_));
 NAND3_X1 _56346_ (.A1(_22524_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2088]),
    .A3(_10942_),
    .ZN(_25123_));
 NAND3_X1 _56347_ (.A1(_23459_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2333]),
    .A3(_23169_),
    .ZN(_25124_));
 OAI21_X1 _56348_ (.A(_25124_),
    .B1(_10946_),
    .B2(_21840_),
    .ZN(_25125_));
 AOI221_X2 _56349_ (.A(_25125_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2235]),
    .B2(_10950_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2186]),
    .C2(_23660_),
    .ZN(_25126_));
 NAND3_X1 _56350_ (.A1(_10781_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2137]),
    .A3(_10942_),
    .ZN(_25127_));
 AOI22_X4 _56351_ (.A1(_23485_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1990]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2039]),
    .B2(_22911_),
    .ZN(_25128_));
 AND4_X4 _56352_ (.A1(_25123_),
    .A2(_25126_),
    .A3(_25127_),
    .A4(_25128_),
    .ZN(_25129_));
 NAND3_X1 _56353_ (.A1(_23340_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1794]),
    .A3(_10990_),
    .ZN(_25130_));
 AND3_X1 _56354_ (.A1(_23524_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1892]),
    .A3(_23662_),
    .ZN(_25131_));
 AOI221_X4 _56355_ (.A(_25131_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1843]),
    .B2(_22044_),
    .C1(_21978_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1941]),
    .ZN(_25132_));
 AOI22_X2 _56356_ (.A1(_23290_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1745]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1696]),
    .B2(_23591_),
    .ZN(_25133_));
 AOI22_X4 _56357_ (.A1(_23595_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1598]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1647]),
    .B2(_23604_),
    .ZN(_25134_));
 AND4_X4 _56358_ (.A1(_25130_),
    .A2(_25132_),
    .A3(_25133_),
    .A4(_25134_),
    .ZN(_25135_));
 AOI22_X4 _56359_ (.A1(_23331_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1157]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1108]),
    .B2(_23333_),
    .ZN(_25136_));
 NAND3_X2 _56360_ (.A1(_22998_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1059]),
    .A3(_23880_),
    .ZN(_25137_));
 OAI211_X4 _56361_ (.A(_25136_),
    .B(_25137_),
    .C1(_22482_),
    .C2(_11096_),
    .ZN(_25138_));
 AOI22_X4 _56362_ (.A1(_23615_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [373]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [324]),
    .B2(_22903_),
    .ZN(_25139_));
 NAND3_X2 _56363_ (.A1(_23062_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [79]),
    .A3(_22951_),
    .ZN(_25140_));
 NAND3_X2 _56364_ (.A1(_23011_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [226]),
    .A3(_23187_),
    .ZN(_25141_));
 NAND3_X2 _56365_ (.A1(_24029_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [275]),
    .A3(_23835_),
    .ZN(_25142_));
 NAND4_X4 _56366_ (.A1(_25139_),
    .A2(_25140_),
    .A3(_25141_),
    .A4(_25142_),
    .ZN(_25143_));
 NAND3_X2 _56367_ (.A1(_22955_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [961]),
    .A3(_22970_),
    .ZN(_25144_));
 NAND3_X2 _56368_ (.A1(_23036_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [863]),
    .A3(_22973_),
    .ZN(_25145_));
 NAND3_X2 _56369_ (.A1(_23078_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [912]),
    .A3(_23891_),
    .ZN(_25146_));
 NAND3_X2 _56370_ (.A1(_23085_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [814]),
    .A3(_23891_),
    .ZN(_25147_));
 NAND4_X4 _56371_ (.A1(_25144_),
    .A2(_25145_),
    .A3(_25146_),
    .A4(_25147_),
    .ZN(_25148_));
 NAND3_X1 _56372_ (.A1(_24045_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [177]),
    .A3(_11176_),
    .ZN(_25149_));
 NAND3_X1 _56373_ (.A1(_23140_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [128]),
    .A3(_23835_),
    .ZN(_25150_));
 NAND3_X1 _56374_ (.A1(_23032_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [30]),
    .A3(_23835_),
    .ZN(_25151_));
 NAND3_X2 _56375_ (.A1(_25149_),
    .A2(_25150_),
    .A3(_25151_),
    .ZN(_25152_));
 NOR4_X4 _56376_ (.A1(_25138_),
    .A2(_25143_),
    .A3(_25148_),
    .A4(_25152_),
    .ZN(_25153_));
 NAND4_X2 _56377_ (.A1(_25122_),
    .A2(_25129_),
    .A3(_25135_),
    .A4(_25153_),
    .ZN(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [30]));
 NAND3_X1 _56378_ (.A1(_23288_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2481]),
    .A3(_23481_),
    .ZN(_25154_));
 NAND3_X4 _56379_ (.A1(_10867_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2824]),
    .A3(_22989_),
    .ZN(_25155_));
 NAND2_X4 _56380_ (.A1(_25154_),
    .A2(_25155_),
    .ZN(_25156_));
 AOI221_X4 _56381_ (.A(_25156_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2089]),
    .B2(_21900_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1746]),
    .C2(_23467_),
    .ZN(_25157_));
 NAND3_X2 _56382_ (.A1(_23166_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2530]),
    .A3(_23012_),
    .ZN(_25158_));
 OAI21_X4 _56383_ (.A(_25158_),
    .B1(_10908_),
    .B2(_21669_),
    .ZN(_25159_));
 AOI221_X4 _56384_ (.A(_25159_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1550]),
    .B2(_23179_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1501]),
    .C2(_23095_),
    .ZN(_25160_));
 NAND3_X2 _56385_ (.A1(_22953_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [962]),
    .A3(_22905_),
    .ZN(_25161_));
 NAND3_X4 _56386_ (.A1(_23284_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2726]),
    .A3(_23481_),
    .ZN(_25162_));
 NAND2_X1 _56387_ (.A1(_25161_),
    .A2(_25162_),
    .ZN(_25163_));
 AOI221_X1 _56388_ (.A(_25163_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2628]),
    .B2(_10902_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [423]),
    .C2(_22733_),
    .ZN(_25164_));
 NAND3_X2 _56389_ (.A1(_23166_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2922]),
    .A3(_10825_),
    .ZN(_25165_));
 OAI21_X4 _56390_ (.A(_25165_),
    .B1(_10852_),
    .B2(_21529_),
    .ZN(_25166_));
 AOI221_X4 _56391_ (.A(_25166_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [374]),
    .B2(_11170_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [227]),
    .C2(_11190_),
    .ZN(_25167_));
 AND4_X2 _56392_ (.A1(_25157_),
    .A2(_25160_),
    .A3(_25164_),
    .A4(_25167_),
    .ZN(_25168_));
 NAND3_X2 _56393_ (.A1(_23150_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1158]),
    .A3(_22905_),
    .ZN(_25169_));
 NAND3_X2 _56394_ (.A1(_22907_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1207]),
    .A3(_11035_),
    .ZN(_25170_));
 NAND2_X4 _56395_ (.A1(_25169_),
    .A2(_25170_),
    .ZN(_25171_));
 AOI221_X2 _56396_ (.A(_25171_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1648]),
    .B2(_11019_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1599]),
    .C2(_23395_),
    .ZN(_25172_));
 NAND3_X1 _56397_ (.A1(_23509_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2138]),
    .A3(_23657_),
    .ZN(_25173_));
 NAND3_X1 _56398_ (.A1(_23382_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1991]),
    .A3(_23657_),
    .ZN(_25174_));
 NAND2_X1 _56399_ (.A1(_25173_),
    .A2(_25174_),
    .ZN(_25175_));
 AOI221_X4 _56400_ (.A(_25175_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1795]),
    .B2(_11002_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1697]),
    .C2(_22105_),
    .ZN(_25176_));
 NAND3_X2 _56401_ (.A1(_23487_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2334]),
    .A3(_23231_),
    .ZN(_25177_));
 NAND3_X2 _56402_ (.A1(_24467_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2236]),
    .A3(_22962_),
    .ZN(_25178_));
 NAND2_X4 _56403_ (.A1(_25177_),
    .A2(_25178_),
    .ZN(_25179_));
 AOI221_X2 _56404_ (.A(_25179_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2040]),
    .B2(_21937_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1060]),
    .C2(_23632_),
    .ZN(_25180_));
 NAND3_X2 _56405_ (.A1(_23810_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1942]),
    .A3(_23519_),
    .ZN(_25181_));
 NAND3_X2 _56406_ (.A1(_23524_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2285]),
    .A3(_23169_),
    .ZN(_25182_));
 NAND2_X4 _56407_ (.A1(_25181_),
    .A2(_25182_),
    .ZN(_25183_));
 AOI221_X2 _56408_ (.A(_25183_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1844]),
    .B2(_22044_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1109]),
    .C2(_23333_),
    .ZN(_25184_));
 AND4_X4 _56409_ (.A1(_25172_),
    .A2(_25176_),
    .A3(_25180_),
    .A4(_25184_),
    .ZN(_25185_));
 NAND3_X1 _56410_ (.A1(_22988_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [570]),
    .A3(_22995_),
    .ZN(_25186_));
 NAND3_X2 _56411_ (.A1(_10880_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [31]),
    .A3(_23341_),
    .ZN(_25187_));
 NAND3_X2 _56412_ (.A1(_23114_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [80]),
    .A3(_23341_),
    .ZN(_25188_));
 NAND3_X2 _56413_ (.A1(_10831_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [668]),
    .A3(_23057_),
    .ZN(_25189_));
 NAND4_X4 _56414_ (.A1(_25186_),
    .A2(_25187_),
    .A3(_25188_),
    .A4(_25189_),
    .ZN(_25190_));
 NAND3_X2 _56415_ (.A1(_23004_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [178]),
    .A3(_22940_),
    .ZN(_25191_));
 NAND3_X4 _56416_ (.A1(_10831_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3020]),
    .A3(_23123_),
    .ZN(_25192_));
 NAND3_X2 _56417_ (.A1(_23127_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3069]),
    .A3(_23128_),
    .ZN(_25193_));
 NAND3_X4 _56418_ (.A1(_23888_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2677]),
    .A3(_23068_),
    .ZN(_25194_));
 NAND4_X4 _56419_ (.A1(_25191_),
    .A2(_25192_),
    .A3(_25193_),
    .A4(_25194_),
    .ZN(_25195_));
 NAND3_X4 _56420_ (.A1(_23020_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1354]),
    .A3(_11037_),
    .ZN(_25196_));
 NAND3_X2 _56421_ (.A1(_23140_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [129]),
    .A3(_22959_),
    .ZN(_25197_));
 NAND3_X1 _56422_ (.A1(_23036_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [472]),
    .A3(_23201_),
    .ZN(_25198_));
 NAND3_X4 _56423_ (.A1(_23145_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1256]),
    .A3(_22981_),
    .ZN(_25199_));
 NAND4_X1 _56424_ (.A1(_25196_),
    .A2(_25197_),
    .A3(_25198_),
    .A4(_25199_),
    .ZN(_25200_));
 NAND3_X1 _56425_ (.A1(_23032_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [815]),
    .A3(_22973_),
    .ZN(_25201_));
 NAND3_X2 _56426_ (.A1(_23276_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1011]),
    .A3(_22976_),
    .ZN(_25202_));
 NAND3_X2 _56427_ (.A1(_23042_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [864]),
    .A3(_23547_),
    .ZN(_25203_));
 NAND3_X2 _56428_ (.A1(_23204_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [913]),
    .A3(_23317_),
    .ZN(_25204_));
 NAND4_X4 _56429_ (.A1(_25201_),
    .A2(_25202_),
    .A3(_25203_),
    .A4(_25204_),
    .ZN(_25205_));
 NOR4_X1 _56430_ (.A1(_25190_),
    .A2(_25195_),
    .A3(_25200_),
    .A4(_25205_),
    .ZN(_25206_));
 AOI22_X4 _56431_ (.A1(_10800_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3118]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1305]),
    .B2(_23262_),
    .ZN(_25207_));
 NAND3_X4 _56432_ (.A1(_23368_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2971]),
    .A3(_23000_),
    .ZN(_25208_));
 OAI211_X4 _56433_ (.A(_25207_),
    .B(_25208_),
    .C1(_21329_),
    .C2(_10875_),
    .ZN(_25209_));
 AOI22_X4 _56434_ (.A1(_22903_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [325]),
    .B1(_23446_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [276]),
    .ZN(_25210_));
 NAND3_X2 _56435_ (.A1(_24050_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [717]),
    .A3(_23060_),
    .ZN(_25211_));
 OAI211_X4 _56436_ (.A(_25210_),
    .B(_25211_),
    .C1(_11121_),
    .C2(_22619_),
    .ZN(_25212_));
 NAND3_X4 _56437_ (.A1(_23192_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2187]),
    .A3(_24052_),
    .ZN(_25213_));
 NAND3_X2 _56438_ (.A1(_10844_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1403]),
    .A3(_23277_),
    .ZN(_25214_));
 NAND3_X1 _56439_ (.A1(_23028_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1893]),
    .A3(_23830_),
    .ZN(_25215_));
 NAND3_X2 _56440_ (.A1(_23080_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1452]),
    .A3(_23205_),
    .ZN(_25216_));
 NAND4_X4 _56441_ (.A1(_25213_),
    .A2(_25214_),
    .A3(_25215_),
    .A4(_25216_),
    .ZN(_25217_));
 NAND3_X4 _56442_ (.A1(_23032_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2383]),
    .A3(_23023_),
    .ZN(_25218_));
 NAND3_X2 _56443_ (.A1(_23271_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [619]),
    .A3(_23072_),
    .ZN(_25219_));
 NAND3_X4 _56444_ (.A1(_23042_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2432]),
    .A3(_23043_),
    .ZN(_25220_));
 NAND3_X2 _56445_ (.A1(_23204_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [521]),
    .A3(_23208_),
    .ZN(_25221_));
 NAND4_X2 _56446_ (.A1(_25218_),
    .A2(_25219_),
    .A3(_25220_),
    .A4(_25221_),
    .ZN(_25222_));
 NOR4_X1 _56447_ (.A1(_25209_),
    .A2(_25212_),
    .A3(_25217_),
    .A4(_25222_),
    .ZN(_25223_));
 NAND4_X1 _56448_ (.A1(_25168_),
    .A2(_25185_),
    .A3(_25206_),
    .A4(_25223_),
    .ZN(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [31]));
 NAND3_X2 _56449_ (.A1(_10817_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [326]),
    .A3(_23643_),
    .ZN(_25224_));
 NAND3_X2 _56450_ (.A1(_10817_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [718]),
    .A3(_23055_),
    .ZN(_25225_));
 NAND2_X4 _56451_ (.A1(_25224_),
    .A2(_25225_),
    .ZN(_25226_));
 AOI221_X4 _56452_ (.A(_25226_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1404]),
    .B2(_23094_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1551]),
    .C2(_23315_),
    .ZN(_25227_));
 NAND3_X1 _56453_ (.A1(_23150_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1943]),
    .A3(_22921_),
    .ZN(_25228_));
 NAND3_X1 _56454_ (.A1(_22915_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1649]),
    .A3(_22921_),
    .ZN(_25229_));
 NAND2_X1 _56455_ (.A1(_25228_),
    .A2(_25229_),
    .ZN(_25230_));
 AOI221_X2 _56456_ (.A(_25230_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1894]),
    .B2(_22003_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1845]),
    .C2(_23286_),
    .ZN(_25231_));
 NAND3_X2 _56457_ (.A1(_23492_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1159]),
    .A3(_22905_),
    .ZN(_25232_));
 NAND3_X2 _56458_ (.A1(_22907_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1208]),
    .A3(_11035_),
    .ZN(_25233_));
 NAND2_X4 _56459_ (.A1(_25232_),
    .A2(_25233_),
    .ZN(_25234_));
 AOI221_X2 _56460_ (.A(_25234_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2090]),
    .B2(_22910_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2041]),
    .C2(_23156_),
    .ZN(_25235_));
 NAND3_X2 _56461_ (.A1(_22953_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [179]),
    .A3(_23643_),
    .ZN(_25236_));
 NAND3_X4 _56462_ (.A1(_23153_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2972]),
    .A3(_23794_),
    .ZN(_25237_));
 NAND2_X4 _56463_ (.A1(_25236_),
    .A2(_25237_),
    .ZN(_25238_));
 AOI221_X4 _56464_ (.A(_25238_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2188]),
    .B2(_10955_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [81]),
    .C2(_23714_),
    .ZN(_25239_));
 AND4_X4 _56465_ (.A1(_25227_),
    .A2(_25231_),
    .A3(_25235_),
    .A4(_25239_),
    .ZN(_25240_));
 NAND3_X4 _56466_ (.A1(_22985_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [571]),
    .A3(_11127_),
    .ZN(_25241_));
 NAND3_X4 _56467_ (.A1(_22988_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2923]),
    .A3(_23361_),
    .ZN(_25242_));
 NAND3_X4 _56468_ (.A1(_10880_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [424]),
    .A3(_22995_),
    .ZN(_25243_));
 NAND3_X4 _56469_ (.A1(_22998_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3021]),
    .A3(_22991_),
    .ZN(_25244_));
 NAND4_X4 _56470_ (.A1(_25241_),
    .A2(_25242_),
    .A3(_25243_),
    .A4(_25244_),
    .ZN(_25245_));
 NAND3_X2 _56471_ (.A1(_23004_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2139]),
    .A3(_23006_),
    .ZN(_25246_));
 NAND3_X2 _56472_ (.A1(_23008_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1600]),
    .A3(_22935_),
    .ZN(_25247_));
 NAND3_X4 _56473_ (.A1(_23059_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2580]),
    .A3(_23131_),
    .ZN(_25248_));
 NAND3_X2 _56474_ (.A1(_10858_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1698]),
    .A3(_23009_),
    .ZN(_25249_));
 NAND4_X4 _56475_ (.A1(_25246_),
    .A2(_25247_),
    .A3(_25248_),
    .A4(_25249_),
    .ZN(_25250_));
 NAND3_X4 _56476_ (.A1(_24045_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2531]),
    .A3(_23131_),
    .ZN(_25251_));
 NAND3_X1 _56477_ (.A1(_23133_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2384]),
    .A3(_23134_),
    .ZN(_25252_));
 NAND3_X1 _56478_ (.A1(_23140_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2482]),
    .A3(_23023_),
    .ZN(_25253_));
 NAND3_X1 _56479_ (.A1(_22961_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2678]),
    .A3(_23026_),
    .ZN(_25254_));
 NAND4_X2 _56480_ (.A1(_25251_),
    .A2(_25252_),
    .A3(_25253_),
    .A4(_25254_),
    .ZN(_25255_));
 NAND3_X1 _56481_ (.A1(_22968_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2776]),
    .A3(_23033_),
    .ZN(_25256_));
 NAND3_X2 _56482_ (.A1(_23189_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2825]),
    .A3(_10790_),
    .ZN(_25257_));
 NAND3_X2 _56483_ (.A1(_23025_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2874]),
    .A3(_23037_),
    .ZN(_25258_));
 NAND3_X2 _56484_ (.A1(_23145_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2433]),
    .A3(_23029_),
    .ZN(_25259_));
 NAND4_X4 _56485_ (.A1(_25256_),
    .A2(_25257_),
    .A3(_25258_),
    .A4(_25259_),
    .ZN(_25260_));
 NOR4_X1 _56486_ (.A1(_25245_),
    .A2(_25250_),
    .A3(_25255_),
    .A4(_25260_),
    .ZN(_25261_));
 AOI22_X2 _56487_ (.A1(_23047_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [963]),
    .B1(_23048_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1257]),
    .ZN(_25262_));
 NAND3_X2 _56488_ (.A1(_22524_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1306]),
    .A3(_23051_),
    .ZN(_25263_));
 OAI211_X4 _56489_ (.A(_25262_),
    .B(_25263_),
    .C1(_22306_),
    .C2(_11055_),
    .ZN(_25264_));
 NAND3_X2 _56490_ (.A1(_23054_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [767]),
    .A3(_23057_),
    .ZN(_25265_));
 NAND3_X1 _56491_ (.A1(_23059_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [620]),
    .A3(_23060_),
    .ZN(_25266_));
 NAND3_X2 _56492_ (.A1(_23062_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [473]),
    .A3(_23060_),
    .ZN(_25267_));
 NAND3_X2 _56493_ (.A1(_23016_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [914]),
    .A3(_22970_),
    .ZN(_25268_));
 NAND4_X4 _56494_ (.A1(_25265_),
    .A2(_25266_),
    .A3(_25267_),
    .A4(_25268_),
    .ZN(_25269_));
 NAND3_X1 _56495_ (.A1(_23067_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2727]),
    .A3(_23014_),
    .ZN(_25270_));
 NAND3_X4 _56496_ (.A1(_23022_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1992]),
    .A3(_22964_),
    .ZN(_25271_));
 NAND3_X4 _56497_ (.A1(_22975_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [669]),
    .A3(_23201_),
    .ZN(_25272_));
 NAND3_X1 _56498_ (.A1(_23071_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2629]),
    .A3(_23029_),
    .ZN(_25273_));
 NAND4_X2 _56499_ (.A1(_25270_),
    .A2(_25271_),
    .A3(_25272_),
    .A4(_25273_),
    .ZN(_25274_));
 NAND3_X4 _56500_ (.A1(_23076_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2335]),
    .A3(_23894_),
    .ZN(_25275_));
 NAND3_X4 _56501_ (.A1(_23078_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [522]),
    .A3(_23201_),
    .ZN(_25276_));
 NAND3_X4 _56502_ (.A1(_23080_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2237]),
    .A3(_23081_),
    .ZN(_25277_));
 NAND3_X4 _56503_ (.A1(_23085_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [32]),
    .A3(_23086_),
    .ZN(_25278_));
 NAND4_X1 _56504_ (.A1(_25275_),
    .A2(_25276_),
    .A3(_25277_),
    .A4(_25278_),
    .ZN(_25279_));
 NOR4_X1 _56505_ (.A1(_25264_),
    .A2(_25269_),
    .A3(_25274_),
    .A4(_25279_),
    .ZN(_25280_));
 AND4_X2 _56506_ (.A1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3070]),
    .A2(_10809_),
    .A3(_22928_),
    .A4(_10795_),
    .ZN(_25281_));
 AOI21_X4 _56507_ (.A(_25281_),
    .B1(_10800_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3119]),
    .ZN(_25282_));
 OAI221_X2 _56508_ (.A(_25282_),
    .B1(_22484_),
    .B2(_11096_),
    .C1(_22569_),
    .C2(_11111_),
    .ZN(_25283_));
 NAND3_X4 _56509_ (.A1(_22933_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1796]),
    .A3(_22935_),
    .ZN(_25284_));
 NAND3_X4 _56510_ (.A1(_23011_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [228]),
    .A3(_22951_),
    .ZN(_25285_));
 NAND3_X4 _56511_ (.A1(_24050_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1502]),
    .A3(_11037_),
    .ZN(_25286_));
 NAND3_X2 _56512_ (.A1(_23140_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [130]),
    .A3(_23835_),
    .ZN(_25287_));
 NAND4_X1 _56513_ (.A1(_25284_),
    .A2(_25285_),
    .A3(_25286_),
    .A4(_25287_),
    .ZN(_25288_));
 NAND3_X2 _56514_ (.A1(_23067_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [375]),
    .A3(_23187_),
    .ZN(_25289_));
 NAND3_X4 _56515_ (.A1(_23200_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1747]),
    .A3(_23830_),
    .ZN(_25290_));
 NAND3_X4 _56516_ (.A1(_23071_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [277]),
    .A3(_23196_),
    .ZN(_25291_));
 NAND3_X4 _56517_ (.A1(_23028_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2286]),
    .A3(_23081_),
    .ZN(_25292_));
 NAND4_X2 _56518_ (.A1(_25289_),
    .A2(_25290_),
    .A3(_25291_),
    .A4(_25292_),
    .ZN(_25293_));
 NAND3_X2 _56519_ (.A1(_23032_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [816]),
    .A3(_22973_),
    .ZN(_25294_));
 NAND3_X1 _56520_ (.A1(_23028_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1110]),
    .A3(_23891_),
    .ZN(_25295_));
 NAND3_X2 _56521_ (.A1(_23575_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1061]),
    .A3(_23547_),
    .ZN(_25296_));
 NAND3_X2 _56522_ (.A1(_23575_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1453]),
    .A3(_23205_),
    .ZN(_25297_));
 NAND4_X4 _56523_ (.A1(_25294_),
    .A2(_25295_),
    .A3(_25296_),
    .A4(_25297_),
    .ZN(_25298_));
 NOR4_X2 _56524_ (.A1(_25283_),
    .A2(_25288_),
    .A3(_25293_),
    .A4(_25298_),
    .ZN(_25299_));
 NAND4_X1 _56525_ (.A1(_25240_),
    .A2(_25261_),
    .A3(_25280_),
    .A4(_25299_),
    .ZN(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [32]));
 AND3_X1 _56526_ (.A1(_23019_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [964]),
    .A3(_22969_),
    .ZN(_25300_));
 AOI21_X2 _56527_ (.A(_25300_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [915]),
    .B2(_23265_),
    .ZN(_25301_));
 OAI221_X2 _56528_ (.A(_25301_),
    .B1(_22451_),
    .B2(_11091_),
    .C1(_22593_),
    .C2(_11115_),
    .ZN(_25302_));
 NAND3_X1 _56529_ (.A1(_24126_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [376]),
    .A3(_23341_),
    .ZN(_25303_));
 NAND3_X1 _56530_ (.A1(_10831_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [278]),
    .A3(_22940_),
    .ZN(_25304_));
 NAND3_X1 _56531_ (.A1(_23377_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [82]),
    .A3(_22940_),
    .ZN(_25305_));
 NAND3_X4 _56532_ (.A1(_23377_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [866]),
    .A3(_23880_),
    .ZN(_25306_));
 NAND4_X2 _56533_ (.A1(_25303_),
    .A2(_25304_),
    .A3(_25305_),
    .A4(_25306_),
    .ZN(_25307_));
 NAND3_X4 _56534_ (.A1(_22933_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2581]),
    .A3(_23131_),
    .ZN(_25308_));
 NAND3_X4 _56535_ (.A1(_23008_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2777]),
    .A3(_23123_),
    .ZN(_25309_));
 NAND3_X2 _56536_ (.A1(_24050_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [327]),
    .A3(_11176_),
    .ZN(_25310_));
 NAND3_X2 _56537_ (.A1(_23189_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2434]),
    .A3(_23068_),
    .ZN(_25311_));
 NAND4_X4 _56538_ (.A1(_25308_),
    .A2(_25309_),
    .A3(_25310_),
    .A4(_25311_),
    .ZN(_25312_));
 NAND3_X2 _56539_ (.A1(_23125_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [572]),
    .A3(_23057_),
    .ZN(_25313_));
 NAND3_X2 _56540_ (.A1(_23062_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [474]),
    .A3(_23063_),
    .ZN(_25314_));
 NAND3_X4 _56541_ (.A1(_23140_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1307]),
    .A3(_23566_),
    .ZN(_25315_));
 NAND3_X2 _56542_ (.A1(_23032_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [425]),
    .A3(_23063_),
    .ZN(_25316_));
 NAND4_X4 _56543_ (.A1(_25313_),
    .A2(_25314_),
    .A3(_25315_),
    .A4(_25316_),
    .ZN(_25317_));
 NOR4_X4 _56544_ (.A1(_25302_),
    .A2(_25307_),
    .A3(_25312_),
    .A4(_25317_),
    .ZN(_25318_));
 AND3_X1 _56545_ (.A1(_10803_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1944]),
    .A3(_10988_),
    .ZN(_25319_));
 AOI21_X4 _56546_ (.A(_25319_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1895]),
    .B2(_22003_),
    .ZN(_25320_));
 AOI22_X4 _56547_ (.A1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [719]),
    .A2(_23092_),
    .B1(_22827_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [131]),
    .ZN(_25321_));
 AOI22_X2 _56548_ (.A1(_23094_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1405]),
    .B1(_23095_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1503]),
    .ZN(_25322_));
 AOI22_X4 _56549_ (.A1(_23097_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2336]),
    .B1(_10976_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1993]),
    .ZN(_25323_));
 AND4_X4 _56550_ (.A1(_25320_),
    .A2(_25321_),
    .A3(_25322_),
    .A4(_25323_),
    .ZN(_25324_));
 NAND3_X2 _56551_ (.A1(_23153_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2973]),
    .A3(_23498_),
    .ZN(_25325_));
 NAND3_X2 _56552_ (.A1(_24467_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3022]),
    .A3(_23794_),
    .ZN(_25326_));
 NAND2_X4 _56553_ (.A1(_25325_),
    .A2(_25326_),
    .ZN(_25327_));
 AOI221_X4 _56554_ (.A(_25327_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [670]),
    .B2(_22642_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [621]),
    .C2(_23515_),
    .ZN(_25328_));
 AND3_X1 _56555_ (.A1(_23390_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1160]),
    .A3(_11081_),
    .ZN(_25329_));
 AOI21_X4 _56556_ (.A(_25329_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1111]),
    .B2(_23333_),
    .ZN(_25330_));
 AOI22_X4 _56557_ (.A1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1209]),
    .A2(_23325_),
    .B1(_22459_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1013]),
    .ZN(_25331_));
 AND4_X4 _56558_ (.A1(_25324_),
    .A2(_25328_),
    .A3(_25330_),
    .A4(_25331_),
    .ZN(_25332_));
 NAND3_X4 _56559_ (.A1(_23221_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [229]),
    .A3(_23709_),
    .ZN(_25333_));
 NAND3_X4 _56560_ (.A1(_10804_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [768]),
    .A3(_11126_),
    .ZN(_25334_));
 NAND3_X4 _56561_ (.A1(_23113_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2042]),
    .A3(_10941_),
    .ZN(_25335_));
 NAND3_X1 _56562_ (.A1(_22523_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2091]),
    .A3(_23553_),
    .ZN(_25336_));
 AND4_X1 _56563_ (.A1(_25333_),
    .A2(_25334_),
    .A3(_25335_),
    .A4(_25336_),
    .ZN(_25337_));
 NAND3_X1 _56564_ (.A1(_23158_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2140]),
    .A3(_23231_),
    .ZN(_25338_));
 NAND3_X1 _56565_ (.A1(_24467_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2238]),
    .A3(_22962_),
    .ZN(_25339_));
 NAND2_X1 _56566_ (.A1(_25338_),
    .A2(_25339_),
    .ZN(_25340_));
 AOI221_X4 _56567_ (.A(_25340_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2287]),
    .B2(_21816_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2189]),
    .C2(_23660_),
    .ZN(_25341_));
 NAND3_X2 _56568_ (.A1(_23173_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2875]),
    .A3(_23174_),
    .ZN(_25342_));
 NAND3_X2 _56569_ (.A1(_23176_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2826]),
    .A3(_10825_),
    .ZN(_25343_));
 NAND2_X4 _56570_ (.A1(_25342_),
    .A2(_25343_),
    .ZN(_25344_));
 AOI221_X4 _56571_ (.A(_25344_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1454]),
    .B2(_22232_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1552]),
    .C2(_23179_),
    .ZN(_25345_));
 NAND3_X1 _56572_ (.A1(_22987_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [180]),
    .A3(_23451_),
    .ZN(_25346_));
 NAND3_X4 _56573_ (.A1(_22523_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [523]),
    .A3(_23056_),
    .ZN(_25347_));
 NAND3_X2 _56574_ (.A1(_23455_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [33]),
    .A3(_22939_),
    .ZN(_25348_));
 NAND3_X4 _56575_ (.A1(_22932_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1797]),
    .A3(_23398_),
    .ZN(_25349_));
 AND4_X4 _56576_ (.A1(_25346_),
    .A2(_25347_),
    .A3(_25348_),
    .A4(_25349_),
    .ZN(_25350_));
 AND4_X4 _56577_ (.A1(_25337_),
    .A2(_25341_),
    .A3(_25345_),
    .A4(_25350_),
    .ZN(_25351_));
 NAND3_X2 _56578_ (.A1(_22988_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1356]),
    .A3(_23051_),
    .ZN(_25352_));
 NAND3_X2 _56579_ (.A1(_23004_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1748]),
    .A3(_23116_),
    .ZN(_25353_));
 NAND3_X2 _56580_ (.A1(_23114_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1258]),
    .A3(_22945_),
    .ZN(_25354_));
 NAND3_X2 _56581_ (.A1(_10831_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1846]),
    .A3(_23116_),
    .ZN(_25355_));
 NAND4_X4 _56582_ (.A1(_25352_),
    .A2(_25353_),
    .A3(_25354_),
    .A4(_25355_),
    .ZN(_25356_));
 NAND3_X2 _56583_ (.A1(_23125_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2532]),
    .A3(_23131_),
    .ZN(_25357_));
 NAND3_X4 _56584_ (.A1(_23560_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3120]),
    .A3(_23128_),
    .ZN(_25358_));
 NAND3_X2 _56585_ (.A1(_23020_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2924]),
    .A3(_23033_),
    .ZN(_25359_));
 NAND3_X4 _56586_ (.A1(_23888_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3071]),
    .A3(_23033_),
    .ZN(_25360_));
 NAND4_X4 _56587_ (.A1(_25357_),
    .A2(_25358_),
    .A3(_25359_),
    .A4(_25360_),
    .ZN(_25361_));
 NAND3_X1 _56588_ (.A1(_23067_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2728]),
    .A3(_23134_),
    .ZN(_25362_));
 NAND3_X1 _56589_ (.A1(_23194_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2385]),
    .A3(_23026_),
    .ZN(_25363_));
 NAND3_X1 _56590_ (.A1(_23071_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2630]),
    .A3(_23029_),
    .ZN(_25364_));
 NAND3_X1 _56591_ (.A1(_23039_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2483]),
    .A3(_23043_),
    .ZN(_25365_));
 NAND4_X2 _56592_ (.A1(_25362_),
    .A2(_25363_),
    .A3(_25364_),
    .A4(_25365_),
    .ZN(_25366_));
 NAND3_X2 _56593_ (.A1(_23022_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1601]),
    .A3(_23141_),
    .ZN(_25367_));
 NAND3_X2 _56594_ (.A1(_23039_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1699]),
    .A3(_23146_),
    .ZN(_25368_));
 NAND3_X4 _56595_ (.A1(_23280_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2679]),
    .A3(_23043_),
    .ZN(_25369_));
 NAND3_X1 _56596_ (.A1(_23426_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1650]),
    .A3(_23576_),
    .ZN(_25370_));
 NAND4_X4 _56597_ (.A1(_25367_),
    .A2(_25368_),
    .A3(_25369_),
    .A4(_25370_),
    .ZN(_25371_));
 NOR4_X2 _56598_ (.A1(_25356_),
    .A2(_25361_),
    .A3(_25366_),
    .A4(_25371_),
    .ZN(_25372_));
 NAND4_X1 _56599_ (.A1(_25318_),
    .A2(_25332_),
    .A3(_25351_),
    .A4(_25372_),
    .ZN(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [33]));
 AND3_X1 _56600_ (.A1(_22920_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [720]),
    .A3(_23504_),
    .ZN(_25373_));
 AOI221_X4 _56601_ (.A(_25373_),
    .B1(_23515_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [622]),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [769]),
    .C2(_23638_),
    .ZN(_25374_));
 NAND3_X1 _56602_ (.A1(_23204_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [132]),
    .A3(_23709_),
    .ZN(_25375_));
 AND3_X1 _56603_ (.A1(_10757_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [573]),
    .A3(_11145_),
    .ZN(_25376_));
 AOI221_X2 _56604_ (.A(_25376_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [524]),
    .B2(_11151_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [426]),
    .C2(_11164_),
    .ZN(_25377_));
 NAND3_X1 _56605_ (.A1(_10780_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [181]),
    .A3(_23246_),
    .ZN(_25378_));
 NAND3_X1 _56606_ (.A1(_22993_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [34]),
    .A3(_23451_),
    .ZN(_25379_));
 AND4_X1 _56607_ (.A1(_25375_),
    .A2(net58),
    .A3(_25378_),
    .A4(_25379_),
    .ZN(_25380_));
 AOI22_X4 _56608_ (.A1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [671]),
    .A2(_23107_),
    .B1(_11159_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [475]),
    .ZN(_25381_));
 NAND3_X1 _56609_ (.A1(_23245_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [377]),
    .A3(_23246_),
    .ZN(_25382_));
 AOI22_X1 _56610_ (.A1(_23248_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [230]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [83]),
    .B2(_11211_),
    .ZN(_25383_));
 NAND3_X1 _56611_ (.A1(_23935_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [328]),
    .A3(_23250_),
    .ZN(_25384_));
 NAND3_X1 _56612_ (.A1(_23252_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [279]),
    .A3(_23250_),
    .ZN(_25385_));
 AND4_X1 _56613_ (.A1(_25382_),
    .A2(_25383_),
    .A3(_25384_),
    .A4(_25385_),
    .ZN(_25386_));
 AND4_X4 _56614_ (.A1(_25374_),
    .A2(_25380_),
    .A3(_25381_),
    .A4(_25386_),
    .ZN(_25387_));
 AND3_X1 _56615_ (.A1(_23721_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2876]),
    .A3(_23498_),
    .ZN(_25388_));
 AOI221_X4 _56616_ (.A(_25388_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2827]),
    .B2(_10863_),
    .C1(_23213_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2925]),
    .ZN(_25389_));
 NAND3_X1 _56617_ (.A1(_23328_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2974]),
    .A3(_23360_),
    .ZN(_25390_));
 AOI22_X2 _56618_ (.A1(_23224_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3121]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3072]),
    .B2(_23225_),
    .ZN(_25391_));
 NAND3_X1 _56619_ (.A1(_10879_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2778]),
    .A3(_22999_),
    .ZN(_25392_));
 NAND3_X1 _56620_ (.A1(_23252_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3023]),
    .A3(_22999_),
    .ZN(_25393_));
 AND4_X4 _56621_ (.A1(_25390_),
    .A2(_25391_),
    .A3(_25392_),
    .A4(_25393_),
    .ZN(_25394_));
 AND3_X1 _56622_ (.A1(_23230_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1994]),
    .A3(_22962_),
    .ZN(_25395_));
 AOI221_X4 _56623_ (.A(_25395_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2092]),
    .B2(_23233_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2141]),
    .C2(_23736_),
    .ZN(_25396_));
 NAND3_X1 _56624_ (.A1(_23935_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2288]),
    .A3(_10941_),
    .ZN(_25397_));
 AOI22_X2 _56625_ (.A1(_10956_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2190]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2043]),
    .B2(_21937_),
    .ZN(_25398_));
 NAND3_X2 _56626_ (.A1(_23757_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2239]),
    .A3(_23388_),
    .ZN(_25399_));
 NAND3_X1 _56627_ (.A1(_23390_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2337]),
    .A3(_23005_),
    .ZN(_25400_));
 AND4_X4 _56628_ (.A1(_25397_),
    .A2(_25398_),
    .A3(_25399_),
    .A4(_25400_),
    .ZN(_25401_));
 AND4_X2 _56629_ (.A1(_25389_),
    .A2(_25394_),
    .A3(_25396_),
    .A4(_25401_),
    .ZN(_25402_));
 NAND3_X1 _56630_ (.A1(_24262_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1553]),
    .A3(_23931_),
    .ZN(_25403_));
 NAND3_X1 _56631_ (.A1(_23339_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1406]),
    .A3(_23412_),
    .ZN(_25404_));
 NAND3_X1 _56632_ (.A1(_22241_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1455]),
    .A3(_23693_),
    .ZN(_25405_));
 NAND3_X1 _56633_ (.A1(_23935_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1504]),
    .A3(_23050_),
    .ZN(_25406_));
 AND4_X4 _56634_ (.A1(_25403_),
    .A2(_25404_),
    .A3(_25405_),
    .A4(_25406_),
    .ZN(_25407_));
 OAI22_X2 _56635_ (.A1(_11115_),
    .A2(_22595_),
    .B1(_22572_),
    .B2(_11111_),
    .ZN(_25408_));
 OAI22_X4 _56636_ (.A1(_11101_),
    .A2(_22515_),
    .B1(_22540_),
    .B2(_11107_),
    .ZN(_25409_));
 AOI211_X2 _56637_ (.A(_25408_),
    .B(_25409_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1063]),
    .C2(_23632_),
    .ZN(_25410_));
 OAI22_X4 _56638_ (.A1(_11070_),
    .A2(_22379_),
    .B1(_22354_),
    .B2(_11066_),
    .ZN(_25411_));
 AOI221_X2 _56639_ (.A(_25411_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1357]),
    .B2(_23748_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1308]),
    .C2(_23262_),
    .ZN(_25412_));
 AND3_X1 _56640_ (.A1(_23459_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1161]),
    .A3(_23460_),
    .ZN(_25413_));
 AOI221_X2 _56641_ (.A(_25413_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1112]),
    .B2(_23332_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1014]),
    .C2(_23104_),
    .ZN(_25414_));
 AND4_X4 _56642_ (.A1(_25407_),
    .A2(_25410_),
    .A3(_25412_),
    .A4(_25414_),
    .ZN(_25415_));
 AND3_X1 _56643_ (.A1(_24467_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1847]),
    .A3(_23519_),
    .ZN(_25416_));
 AOI221_X4 _56644_ (.A(_25416_),
    .B1(_22003_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1896]),
    .C1(_23584_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1945]),
    .ZN(_25417_));
 AND3_X1 _56645_ (.A1(_23288_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1700]),
    .A3(_10988_),
    .ZN(_25418_));
 AOI21_X1 _56646_ (.A(_25418_),
    .B1(_23467_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1749]),
    .ZN(_25419_));
 NAND3_X1 _56647_ (.A1(_10879_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1602]),
    .A3(_10989_),
    .ZN(_25420_));
 NAND3_X1 _56648_ (.A1(_23293_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1651]),
    .A3(_23294_),
    .ZN(_25421_));
 NAND3_X1 _56649_ (.A1(_23296_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1798]),
    .A3(_23398_),
    .ZN(_25422_));
 AND4_X4 _56650_ (.A1(_25419_),
    .A2(_25420_),
    .A3(_25421_),
    .A4(_25422_),
    .ZN(_25423_));
 NAND3_X1 _56651_ (.A1(_22987_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2533]),
    .A3(_10892_),
    .ZN(_25424_));
 AOI22_X2 _56652_ (.A1(_23300_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2386]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2435]),
    .B2(_23301_),
    .ZN(_25425_));
 NAND3_X1 _56653_ (.A1(_23303_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2631]),
    .A3(_23304_),
    .ZN(_25426_));
 NAND3_X1 _56654_ (.A1(_23306_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2484]),
    .A3(_23304_),
    .ZN(_25427_));
 AND4_X4 _56655_ (.A1(_25424_),
    .A2(_25425_),
    .A3(_25426_),
    .A4(_25427_),
    .ZN(_25428_));
 AND3_X1 _56656_ (.A1(_23217_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2729]),
    .A3(_23310_),
    .ZN(_25429_));
 AOI221_X2 _56657_ (.A(_25429_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2680]),
    .B2(_21600_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2582]),
    .C2(_21654_),
    .ZN(_25430_));
 AND4_X2 _56658_ (.A1(_25417_),
    .A2(_25423_),
    .A3(_25428_),
    .A4(_25430_),
    .ZN(_25431_));
 NAND4_X1 _56659_ (.A1(_25387_),
    .A2(_25402_),
    .A3(_25415_),
    .A4(_25431_),
    .ZN(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [34]));
 NAND3_X1 _56660_ (.A1(_23340_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [231]),
    .A3(_23341_),
    .ZN(_25432_));
 NAND3_X2 _56661_ (.A1(_23221_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [623]),
    .A3(_23237_),
    .ZN(_25433_));
 AND3_X1 _56662_ (.A1(_10757_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [574]),
    .A3(_11145_),
    .ZN(_25434_));
 AOI221_X2 _56663_ (.A(_25434_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [525]),
    .B2(_11151_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [427]),
    .C2(_11164_),
    .ZN(_25435_));
 AND3_X1 _56664_ (.A1(_10797_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [770]),
    .A3(_11145_),
    .ZN(_25436_));
 AOI221_X2 _56665_ (.A(_25436_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [721]),
    .B2(_11131_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [672]),
    .C2(_11136_),
    .ZN(_25437_));
 NAND3_X1 _56666_ (.A1(_23113_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [476]),
    .A3(_11126_),
    .ZN(_25438_));
 AND4_X4 _56667_ (.A1(_25433_),
    .A2(_25435_),
    .A3(_25437_),
    .A4(_25438_),
    .ZN(_25439_));
 AND3_X1 _56668_ (.A1(_22942_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [329]),
    .A3(_23159_),
    .ZN(_25440_));
 AOI221_X4 _56669_ (.A(_25440_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [280]),
    .B2(_22777_),
    .C1(_23615_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [378]),
    .ZN(_25441_));
 NAND3_X1 _56670_ (.A1(_22907_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [35]),
    .A3(_23643_),
    .ZN(_25442_));
 NAND3_X1 _56671_ (.A1(_23775_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [84]),
    .A3(_23159_),
    .ZN(_25443_));
 NAND2_X1 _56672_ (.A1(_25442_),
    .A2(_25443_),
    .ZN(_25444_));
 AOI221_X4 _56673_ (.A(_25444_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [133]),
    .B2(_23453_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [182]),
    .C2(_22806_),
    .ZN(_25445_));
 AND4_X4 _56674_ (.A1(_25432_),
    .A2(_25439_),
    .A3(_25441_),
    .A4(_25445_),
    .ZN(_25446_));
 AND3_X1 _56675_ (.A1(_10856_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2485]),
    .A3(_23012_),
    .ZN(_25447_));
 AOI221_X2 _56676_ (.A(_25447_),
    .B1(_23300_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2387]),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2534]),
    .C2(_23587_),
    .ZN(_25448_));
 NAND3_X2 _56677_ (.A1(_10869_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2828]),
    .A3(_23361_),
    .ZN(_25449_));
 NAND3_X1 _56678_ (.A1(_22524_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2877]),
    .A3(_23361_),
    .ZN(_25450_));
 NAND3_X2 _56679_ (.A1(_10781_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2926]),
    .A3(_23361_),
    .ZN(_25451_));
 NAND4_X4 _56680_ (.A1(_25448_),
    .A2(_25449_),
    .A3(_25450_),
    .A4(_25451_),
    .ZN(_25452_));
 AOI22_X4 _56681_ (.A1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2779]),
    .A2(_23625_),
    .B1(_10839_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2975]),
    .ZN(_25453_));
 NAND3_X2 _56682_ (.A1(_10819_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3073]),
    .A3(_22991_),
    .ZN(_25454_));
 NAND3_X2 _56683_ (.A1(_22242_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3024]),
    .A3(_22991_),
    .ZN(_25455_));
 NAND3_X2 _56684_ (.A1(_24126_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3122]),
    .A3(_23000_),
    .ZN(_25456_));
 NAND4_X4 _56685_ (.A1(_25453_),
    .A2(_25454_),
    .A3(_25455_),
    .A4(_25456_),
    .ZN(_25457_));
 AOI22_X4 _56686_ (.A1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2632]),
    .A2(_23627_),
    .B1(_10922_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2436]),
    .ZN(_25458_));
 NAND3_X2 _56687_ (.A1(_22944_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2681]),
    .A3(_23120_),
    .ZN(_25459_));
 NAND3_X2 _56688_ (.A1(_23368_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2583]),
    .A3(_23120_),
    .ZN(_25460_));
 NAND3_X2 _56689_ (.A1(_24126_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2730]),
    .A3(_23120_),
    .ZN(_25461_));
 NAND4_X4 _56690_ (.A1(_25458_),
    .A2(_25459_),
    .A3(_25460_),
    .A4(_25461_),
    .ZN(_25462_));
 NOR3_X2 _56691_ (.A1(_25452_),
    .A2(_25457_),
    .A3(_25462_),
    .ZN(_25463_));
 AND3_X1 _56692_ (.A1(_23153_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1407]),
    .A3(_23848_),
    .ZN(_25464_));
 AOI221_X4 _56693_ (.A(_25464_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1505]),
    .B2(_22210_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1554]),
    .C2(_23179_),
    .ZN(_25465_));
 NAND3_X1 _56694_ (.A1(_23339_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1015]),
    .A3(_23329_),
    .ZN(_25466_));
 AOI22_X1 _56695_ (.A1(_23331_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1162]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1113]),
    .B2(_22410_),
    .ZN(_25467_));
 NAND3_X1 _56696_ (.A1(_23252_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1064]),
    .A3(_11081_),
    .ZN(_25468_));
 NAND3_X1 _56697_ (.A1(_23293_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [868]),
    .A3(_23879_),
    .ZN(_25469_));
 AND4_X2 _56698_ (.A1(_25466_),
    .A2(_25467_),
    .A3(_25468_),
    .A4(_25469_),
    .ZN(_25470_));
 AOI22_X2 _56699_ (.A1(_23325_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1211]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1456]),
    .B2(_23326_),
    .ZN(_25471_));
 NAND3_X2 _56700_ (.A1(_23019_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [966]),
    .A3(_23879_),
    .ZN(_25472_));
 NAND3_X2 _56701_ (.A1(_10857_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [917]),
    .A3(_23879_),
    .ZN(_25473_));
 NAND3_X2 _56702_ (.A1(_22967_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [819]),
    .A3(_22969_),
    .ZN(_25474_));
 NAND3_X4 _56703_ (.A1(_25472_),
    .A2(_25473_),
    .A3(_25474_),
    .ZN(_25475_));
 AND3_X1 _56704_ (.A1(_22954_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1358]),
    .A3(_11036_),
    .ZN(_25476_));
 AND3_X1 _56705_ (.A1(_22522_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1309]),
    .A3(_22980_),
    .ZN(_25477_));
 AND3_X1 _56706_ (.A1(_23041_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1260]),
    .A3(_22980_),
    .ZN(_25478_));
 NOR4_X1 _56707_ (.A1(_25475_),
    .A2(_25476_),
    .A3(_25477_),
    .A4(_25478_),
    .ZN(_25479_));
 AND4_X4 _56708_ (.A1(_25465_),
    .A2(_25470_),
    .A3(_25471_),
    .A4(_25479_),
    .ZN(_25480_));
 AND3_X1 _56709_ (.A1(_23382_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1995]),
    .A3(_23231_),
    .ZN(_25481_));
 AOI221_X4 _56710_ (.A(_25481_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2093]),
    .B2(_23233_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2142]),
    .C2(_10962_),
    .ZN(_25482_));
 NAND3_X1 _56711_ (.A1(_10780_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1750]),
    .A3(_23393_),
    .ZN(_25483_));
 AOI22_X4 _56712_ (.A1(_23395_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1603]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1652]),
    .B2(_23396_),
    .ZN(_25484_));
 NAND3_X1 _56713_ (.A1(_23296_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1799]),
    .A3(_23294_),
    .ZN(_25485_));
 NAND3_X1 _56714_ (.A1(_23306_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1701]),
    .A3(_23398_),
    .ZN(_25486_));
 AND4_X4 _56715_ (.A1(_25483_),
    .A2(_25484_),
    .A3(_25485_),
    .A4(_25486_),
    .ZN(_25487_));
 NAND3_X1 _56716_ (.A1(_22997_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2240]),
    .A3(_23553_),
    .ZN(_25488_));
 AOI22_X1 _56717_ (.A1(_23660_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2191]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2044]),
    .B2(_21937_),
    .ZN(_25489_));
 NAND3_X1 _56718_ (.A1(_22943_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2289]),
    .A3(_23005_),
    .ZN(_25490_));
 NAND3_X1 _56719_ (.A1(_22949_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2338]),
    .A3(_23005_),
    .ZN(_25491_));
 AND4_X1 _56720_ (.A1(_25488_),
    .A2(_25489_),
    .A3(_25490_),
    .A4(_25491_),
    .ZN(_25492_));
 AND3_X1 _56721_ (.A1(_23408_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1897]),
    .A3(_23402_),
    .ZN(_25493_));
 AOI221_X4 _56722_ (.A(_25493_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1848]),
    .B2(_10997_),
    .C1(_21978_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1946]),
    .ZN(_25494_));
 AND4_X4 _56723_ (.A1(_25482_),
    .A2(_25487_),
    .A3(_25492_),
    .A4(_25494_),
    .ZN(_25495_));
 NAND4_X1 _56724_ (.A1(_25446_),
    .A2(_25463_),
    .A3(_25480_),
    .A4(_25495_),
    .ZN(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [35]));
 NAND3_X1 _56725_ (.A1(_23083_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [820]),
    .A3(_23460_),
    .ZN(_25496_));
 NAND3_X1 _56726_ (.A1(_23176_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [869]),
    .A3(_23460_),
    .ZN(_25497_));
 NAND2_X1 _56727_ (.A1(_25496_),
    .A2(_25497_),
    .ZN(_25498_));
 AOI221_X2 _56728_ (.A(_25498_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [967]),
    .B2(_11100_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [918]),
    .C2(_23265_),
    .ZN(_25499_));
 AND3_X1 _56729_ (.A1(_10798_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1163]),
    .A3(_23938_),
    .ZN(_25500_));
 AOI221_X2 _56730_ (.A(_25500_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1114]),
    .B2(_23332_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1065]),
    .C2(_22435_),
    .ZN(_25501_));
 OAI211_X4 _56731_ (.A(net21),
    .B(net43),
    .C1(_22486_),
    .C2(_11096_),
    .ZN(_25502_));
 AND3_X1 _56732_ (.A1(_10798_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2731]),
    .A3(_10890_),
    .ZN(_25503_));
 AOI221_X2 _56733_ (.A(_25503_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2682]),
    .B2(_21600_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2633]),
    .C2(_23627_),
    .ZN(_25504_));
 AOI22_X2 _56734_ (.A1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2584]),
    .A2(_21654_),
    .B1(_10929_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2388]),
    .ZN(_25505_));
 AND3_X1 _56735_ (.A1(_22521_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2486]),
    .A3(_10890_),
    .ZN(_25506_));
 AOI221_X2 _56736_ (.A(_25506_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2437]),
    .B2(_10921_),
    .C1(_10912_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2535]),
    .ZN(_25507_));
 AND3_X1 _56737_ (.A1(_10866_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2829]),
    .A3(_10825_),
    .ZN(_25508_));
 AOI221_X2 _56738_ (.A(_25508_),
    .B1(_10851_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2878]),
    .C1(_21466_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2927]),
    .ZN(_25509_));
 NAND4_X4 _56739_ (.A1(_25504_),
    .A2(_25505_),
    .A3(_25507_),
    .A4(_25509_),
    .ZN(_25510_));
 AOI22_X4 _56740_ (.A1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2780]),
    .A2(_23625_),
    .B1(_10839_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2976]),
    .ZN(_25511_));
 NAND3_X2 _56741_ (.A1(_22950_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3123]),
    .A3(_23123_),
    .ZN(_25512_));
 NAND3_X2 _56742_ (.A1(_23536_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3025]),
    .A3(_23128_),
    .ZN(_25513_));
 NAND3_X2 _56743_ (.A1(_23888_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3074]),
    .A3(_23033_),
    .ZN(_25514_));
 NAND4_X4 _56744_ (.A1(_25511_),
    .A2(_25512_),
    .A3(_25513_),
    .A4(_25514_),
    .ZN(_25515_));
 AND3_X1 _56745_ (.A1(_10824_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [281]),
    .A3(_22937_),
    .ZN(_25516_));
 AOI221_X2 _56746_ (.A(_25516_),
    .B1(_11181_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [330]),
    .C1(_11170_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [379]),
    .ZN(_25517_));
 NAND3_X2 _56747_ (.A1(_23011_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [232]),
    .A3(_23187_),
    .ZN(_25518_));
 AOI22_X2 _56748_ (.A1(_11196_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [183]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [134]),
    .B2(_22827_),
    .ZN(_25519_));
 AOI22_X4 _56749_ (.A1(_11206_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [36]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [85]),
    .B2(_23490_),
    .ZN(_25520_));
 NAND4_X4 _56750_ (.A1(_25517_),
    .A2(_25518_),
    .A3(_25519_),
    .A4(_25520_),
    .ZN(_25521_));
 NOR4_X1 _56751_ (.A1(_25502_),
    .A2(_25510_),
    .A3(_25515_),
    .A4(_25521_),
    .ZN(_25522_));
 AND3_X1 _56752_ (.A1(_22953_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2143]),
    .A3(_22913_),
    .ZN(_25523_));
 AOI221_X4 _56753_ (.A(_25523_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2094]),
    .B2(_22910_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1996]),
    .C2(_23485_),
    .ZN(_25524_));
 NAND3_X1 _56754_ (.A1(_23339_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1800]),
    .A3(_23393_),
    .ZN(_25525_));
 AND3_X1 _56755_ (.A1(_10811_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1898]),
    .A3(_10982_),
    .ZN(_25526_));
 AOI221_X2 _56756_ (.A(_25526_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1849]),
    .B2(_10997_),
    .C1(_10983_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1947]),
    .ZN(_25527_));
 AOI22_X2 _56757_ (.A1(_23467_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1751]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1702]),
    .B2(_22105_),
    .ZN(_25528_));
 AOI22_X2 _56758_ (.A1(_23395_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1604]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1653]),
    .B2(_23396_),
    .ZN(_25529_));
 AND4_X4 _56759_ (.A1(_25525_),
    .A2(_25527_),
    .A3(_25528_),
    .A4(_25529_),
    .ZN(_25530_));
 AND3_X1 _56760_ (.A1(_23168_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2241]),
    .A3(_22962_),
    .ZN(_25531_));
 AOI221_X4 _56761_ (.A(_25531_),
    .B1(_21816_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2290]),
    .C1(_23097_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2339]),
    .ZN(_25532_));
 AOI22_X2 _56762_ (.A1(_10956_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2192]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2045]),
    .B2(_22911_),
    .ZN(_25533_));
 AND4_X4 _56763_ (.A1(_25524_),
    .A2(_25530_),
    .A3(_25532_),
    .A4(_25533_),
    .ZN(_25534_));
 NAND3_X1 _56764_ (.A1(_23340_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1408]),
    .A3(_23051_),
    .ZN(_25535_));
 AND3_X1 _56765_ (.A1(_23733_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1261]),
    .A3(_23701_),
    .ZN(_25536_));
 AOI221_X4 _56766_ (.A(_25536_),
    .B1(_11060_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1310]),
    .C1(_22282_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1359]),
    .ZN(_25537_));
 AOI22_X2 _56767_ (.A1(_23315_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1555]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1506]),
    .B2(_23095_),
    .ZN(_25538_));
 AOI22_X4 _56768_ (.A1(_23325_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1212]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1457]),
    .B2(_23326_),
    .ZN(_25539_));
 AND4_X4 _56769_ (.A1(_25535_),
    .A2(_25537_),
    .A3(_25538_),
    .A4(_25539_),
    .ZN(_25540_));
 NAND3_X1 _56770_ (.A1(_22242_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [673]),
    .A3(_11127_),
    .ZN(_25541_));
 AND3_X1 _56771_ (.A1(_23230_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [428]),
    .A3(_23255_),
    .ZN(_25542_));
 AOI221_X4 _56772_ (.A(_25542_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [526]),
    .B2(_11152_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [575]),
    .C2(_11147_),
    .ZN(_25543_));
 AND3_X1 _56773_ (.A1(_23408_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [722]),
    .A3(_23255_),
    .ZN(_25544_));
 AOI221_X4 _56774_ (.A(_25544_),
    .B1(_23515_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [624]),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [771]),
    .C2(_22597_),
    .ZN(_25545_));
 NAND3_X1 _56775_ (.A1(_10869_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [477]),
    .A3(_11127_),
    .ZN(_25546_));
 AND4_X4 _56776_ (.A1(_25541_),
    .A2(_25543_),
    .A3(_25545_),
    .A4(_25546_),
    .ZN(_25547_));
 NAND4_X1 _56777_ (.A1(_25522_),
    .A2(_25534_),
    .A3(_25540_),
    .A4(_25547_),
    .ZN(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [36]));
 NAND3_X2 _56778_ (.A1(_23194_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2389]),
    .A3(_23143_),
    .ZN(_25548_));
 AND3_X1 _56779_ (.A1(_10866_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2830]),
    .A3(_10787_),
    .ZN(_25549_));
 AOI221_X2 _56780_ (.A(_25549_),
    .B1(_10851_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2879]),
    .C1(_10773_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2928]),
    .ZN(_25550_));
 NAND3_X1 _56781_ (.A1(_23204_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2487]),
    .A3(_23422_),
    .ZN(_25551_));
 NAND3_X1 _56782_ (.A1(_23421_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2536]),
    .A3(_23422_),
    .ZN(_25552_));
 AND4_X1 _56783_ (.A1(_25548_),
    .A2(_25550_),
    .A3(_25551_),
    .A4(_25552_),
    .ZN(_25553_));
 NAND3_X2 _56784_ (.A1(_23080_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3026]),
    .A3(_23037_),
    .ZN(_25554_));
 AOI22_X2 _56785_ (.A1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2781]),
    .A2(_23625_),
    .B1(_10839_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2977]),
    .ZN(_25555_));
 NAND3_X1 _56786_ (.A1(_24186_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3075]),
    .A3(_23673_),
    .ZN(_25556_));
 NAND3_X2 _56787_ (.A1(_23236_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3124]),
    .A3(_23673_),
    .ZN(_25557_));
 AND4_X4 _56788_ (.A1(_25554_),
    .A2(_25555_),
    .A3(_25556_),
    .A4(_25557_),
    .ZN(_25558_));
 NAND3_X1 _56789_ (.A1(_23426_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2438]),
    .A3(_23422_),
    .ZN(_25559_));
 AOI22_X2 _56790_ (.A1(_23373_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2732]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2683]),
    .B2(_23374_),
    .ZN(_25560_));
 NAND3_X1 _56791_ (.A1(_23434_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2634]),
    .A3(_23427_),
    .ZN(_25561_));
 NAND3_X1 _56792_ (.A1(_23221_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2585]),
    .A3(_23427_),
    .ZN(_25562_));
 AND4_X4 _56793_ (.A1(_25559_),
    .A2(_25560_),
    .A3(_25561_),
    .A4(_25562_),
    .ZN(_25563_));
 AND3_X2 _56794_ (.A1(_25553_),
    .A2(_25558_),
    .A3(_25563_),
    .ZN(_25564_));
 AOI22_X4 _56795_ (.A1(_23622_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [576]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [527]),
    .B2(_11153_),
    .ZN(_25565_));
 AOI22_X4 _56796_ (.A1(_23610_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [429]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [478]),
    .B2(_11159_),
    .ZN(_25566_));
 OAI211_X4 _56797_ (.A(_25565_),
    .B(_25566_),
    .C1(_22661_),
    .C2(_11137_),
    .ZN(_25567_));
 NAND3_X1 _56798_ (.A1(_23560_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [772]),
    .A3(_23060_),
    .ZN(_25568_));
 OAI221_X2 _56799_ (.A(_25568_),
    .B1(_11132_),
    .B2(_22640_),
    .C1(_11142_),
    .C2(_22684_),
    .ZN(_25569_));
 AOI22_X4 _56800_ (.A1(_23325_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1213]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1262]),
    .B2(_23048_),
    .ZN(_25570_));
 NAND3_X2 _56801_ (.A1(_23140_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1311]),
    .A3(_23566_),
    .ZN(_25571_));
 NAND3_X2 _56802_ (.A1(_23200_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1360]),
    .A3(_23274_),
    .ZN(_25572_));
 NAND3_X2 _56803_ (.A1(_22958_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1458]),
    .A3(_23277_),
    .ZN(_25573_));
 NAND4_X4 _56804_ (.A1(_25570_),
    .A2(_25571_),
    .A3(_25572_),
    .A4(_25573_),
    .ZN(_25574_));
 NAND3_X2 _56805_ (.A1(_22950_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1556]),
    .A3(_22945_),
    .ZN(_25575_));
 NAND3_X2 _56806_ (.A1(_23127_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1507]),
    .A3(_24026_),
    .ZN(_25576_));
 NAND3_X2 _56807_ (.A1(_23011_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1409]),
    .A3(_11037_),
    .ZN(_25577_));
 NAND3_X4 _56808_ (.A1(_25575_),
    .A2(_25576_),
    .A3(_25577_),
    .ZN(_25578_));
 NOR4_X4 _56809_ (.A1(_25567_),
    .A2(_25569_),
    .A3(_25574_),
    .A4(_25578_),
    .ZN(_25579_));
 AOI22_X4 _56810_ (.A1(_23290_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1752]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1703]),
    .B2(_23591_),
    .ZN(_25580_));
 AOI22_X4 _56811_ (.A1(_23595_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1605]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1654]),
    .B2(_23604_),
    .ZN(_25581_));
 OAI211_X4 _56812_ (.A(_25580_),
    .B(_25581_),
    .C1(_22076_),
    .C2(_11004_),
    .ZN(_25582_));
 NAND3_X4 _56813_ (.A1(_23536_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1850]),
    .A3(_23009_),
    .ZN(_25583_));
 OAI221_X2 _56814_ (.A(_25583_),
    .B1(_10994_),
    .B2(_22038_),
    .C1(_10984_),
    .C2(_21993_),
    .ZN(_25584_));
 AOI22_X4 _56815_ (.A1(_23485_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1997]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2046]),
    .B2(_22911_),
    .ZN(_25585_));
 NAND3_X4 _56816_ (.A1(_23200_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2144]),
    .A3(_22964_),
    .ZN(_25586_));
 OAI211_X4 _56817_ (.A(_25585_),
    .B(_25586_),
    .C1(_21929_),
    .C2(_10969_),
    .ZN(_25587_));
 NAND3_X2 _56818_ (.A1(_23076_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2340]),
    .A3(_23894_),
    .ZN(_25588_));
 NAND3_X2 _56819_ (.A1(_22961_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2291]),
    .A3(_23832_),
    .ZN(_25589_));
 NAND3_X1 _56820_ (.A1(_23839_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2193]),
    .A3(_23081_),
    .ZN(_25590_));
 NAND3_X2 _56821_ (.A1(_23575_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2242]),
    .A3(_23600_),
    .ZN(_25591_));
 NAND4_X4 _56822_ (.A1(_25588_),
    .A2(_25589_),
    .A3(_25590_),
    .A4(_25591_),
    .ZN(_25592_));
 NOR4_X4 _56823_ (.A1(_25582_),
    .A2(_25584_),
    .A3(_25587_),
    .A4(_25592_),
    .ZN(_25593_));
 AOI22_X4 _56824_ (.A1(_23331_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1164]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1115]),
    .B2(_23333_),
    .ZN(_25594_));
 NAND3_X2 _56825_ (.A1(_22998_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1066]),
    .A3(_23880_),
    .ZN(_25595_));
 OAI211_X4 _56826_ (.A(_25594_),
    .B(_25595_),
    .C1(_22488_),
    .C2(_11096_),
    .ZN(_25596_));
 AOI22_X4 _56827_ (.A1(_11206_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [37]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [86]),
    .B2(_23490_),
    .ZN(_25597_));
 NAND3_X4 _56828_ (.A1(_23020_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [184]),
    .A3(_11176_),
    .ZN(_25598_));
 OAI211_X4 _56829_ (.A(_25597_),
    .B(_25598_),
    .C1(_22855_),
    .C2(_11201_),
    .ZN(_25599_));
 NAND3_X2 _56830_ (.A1(_22955_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [968]),
    .A3(_22970_),
    .ZN(_25600_));
 NAND3_X2 _56831_ (.A1(_23036_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [870]),
    .A3(_22976_),
    .ZN(_25601_));
 NAND3_X2 _56832_ (.A1(_23078_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [919]),
    .A3(_23891_),
    .ZN(_25602_));
 NAND3_X2 _56833_ (.A1(_23085_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [821]),
    .A3(_23547_),
    .ZN(_25603_));
 NAND4_X4 _56834_ (.A1(_25600_),
    .A2(_25601_),
    .A3(_25602_),
    .A4(_25603_),
    .ZN(_25604_));
 NAND3_X1 _56835_ (.A1(_23076_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [380]),
    .A3(_23835_),
    .ZN(_25605_));
 NAND3_X1 _56836_ (.A1(_22978_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [282]),
    .A3(_23196_),
    .ZN(_25606_));
 NAND3_X1 _56837_ (.A1(_23839_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [233]),
    .A3(_23086_),
    .ZN(_25607_));
 NAND3_X1 _56838_ (.A1(_23280_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [331]),
    .A3(_23086_),
    .ZN(_25608_));
 NAND4_X2 _56839_ (.A1(_25605_),
    .A2(_25606_),
    .A3(_25607_),
    .A4(_25608_),
    .ZN(_25609_));
 NOR4_X4 _56840_ (.A1(_25596_),
    .A2(_25599_),
    .A3(_25604_),
    .A4(_25609_),
    .ZN(_25610_));
 NAND4_X1 _56841_ (.A1(_25564_),
    .A2(net2),
    .A3(_25593_),
    .A4(_25610_),
    .ZN(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [37]));
 NAND3_X2 _56842_ (.A1(_22953_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2145]),
    .A3(_22913_),
    .ZN(_25611_));
 NAND3_X2 _56843_ (.A1(_10878_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1998]),
    .A3(_22913_),
    .ZN(_25612_));
 NAND2_X4 _56844_ (.A1(_25611_),
    .A2(_25612_),
    .ZN(_25613_));
 AOI221_X4 _56845_ (.A(_25613_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [920]),
    .B2(_23265_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [871]),
    .C2(_22544_),
    .ZN(_25614_));
 OAI22_X4 _56846_ (.A1(_21812_),
    .A2(_10937_),
    .B1(_11009_),
    .B2(_22101_),
    .ZN(_25615_));
 AOI221_X2 _56847_ (.A(_25615_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2439]),
    .B2(_10921_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1655]),
    .C2(_23604_),
    .ZN(_25616_));
 OAI22_X4 _56848_ (.A1(_10897_),
    .A2(_21623_),
    .B1(_22792_),
    .B2(_11187_),
    .ZN(_25617_));
 AOI221_X2 _56849_ (.A(_25617_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3076]),
    .B2(_23225_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [87]),
    .C2(_23714_),
    .ZN(_25618_));
 NAND3_X4 _56850_ (.A1(_22907_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [430]),
    .A3(_23510_),
    .ZN(_25619_));
 NAND3_X4 _56851_ (.A1(_23153_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1410]),
    .A3(_23848_),
    .ZN(_25620_));
 NAND2_X2 _56852_ (.A1(_25619_),
    .A2(_25620_),
    .ZN(_25621_));
 AOI221_X4 _56853_ (.A(_25621_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1312]),
    .B2(_11060_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [136]),
    .C2(_22827_),
    .ZN(_25622_));
 AND4_X1 _56854_ (.A1(_25614_),
    .A2(net20),
    .A3(net19),
    .A4(_25622_),
    .ZN(_25623_));
 AOI22_X4 _56855_ (.A1(_23587_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2537]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2831]),
    .B2(_21536_),
    .ZN(_25624_));
 NAND3_X2 _56856_ (.A1(_22242_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1851]),
    .A3(_10990_),
    .ZN(_25625_));
 OAI211_X4 _56857_ (.A(_25624_),
    .B(_25625_),
    .C1(_21996_),
    .C2(_10984_),
    .ZN(_25626_));
 AOI22_X4 _56858_ (.A1(_23591_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1704]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2047]),
    .B2(_22911_),
    .ZN(_25627_));
 OAI221_X2 _56859_ (.A(_25627_),
    .B1(_10852_),
    .B2(_21532_),
    .C1(_21732_),
    .C2(_10917_),
    .ZN(_25628_));
 NAND3_X4 _56860_ (.A1(_24045_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2929]),
    .A3(_23128_),
    .ZN(_25629_));
 NAND3_X2 _56861_ (.A1(_23192_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1802]),
    .A3(_22956_),
    .ZN(_25630_));
 NAND3_X2 _56862_ (.A1(_23888_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2292]),
    .A3(_22964_),
    .ZN(_25631_));
 NAND3_X2 _56863_ (.A1(_23025_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2096]),
    .A3(_22964_),
    .ZN(_25632_));
 NAND4_X4 _56864_ (.A1(_25629_),
    .A2(_25630_),
    .A3(_25631_),
    .A4(_25632_),
    .ZN(_25633_));
 NAND3_X2 _56865_ (.A1(_23192_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2194]),
    .A3(_24052_),
    .ZN(_25634_));
 NAND3_X4 _56866_ (.A1(_23022_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1606]),
    .A3(_23141_),
    .ZN(_25635_));
 NAND3_X2 _56867_ (.A1(_22961_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1900]),
    .A3(_23830_),
    .ZN(_25636_));
 NAND3_X2 _56868_ (.A1(_22978_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2243]),
    .A3(_23832_),
    .ZN(_25637_));
 NAND4_X4 _56869_ (.A1(_25634_),
    .A2(_25635_),
    .A3(_25636_),
    .A4(_25637_),
    .ZN(_25638_));
 NOR4_X4 _56870_ (.A1(_25626_),
    .A2(_25628_),
    .A3(_25633_),
    .A4(_25638_),
    .ZN(_25639_));
 NAND3_X2 _56871_ (.A1(_23810_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1557]),
    .A3(_23701_),
    .ZN(_25640_));
 OAI21_X4 _56872_ (.A(_25640_),
    .B1(_11042_),
    .B2(_22226_),
    .ZN(_25641_));
 AOI221_X2 _56873_ (.A(_25641_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1263]),
    .B2(_11065_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [724]),
    .C2(_23092_),
    .ZN(_25642_));
 NAND3_X2 _56874_ (.A1(_23309_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [234]),
    .A3(_22937_),
    .ZN(_25643_));
 OAI21_X4 _56875_ (.A(_25643_),
    .B1(_11171_),
    .B2(_22755_),
    .ZN(_25644_));
 AOI221_X1 _56876_ (.A(_25644_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1459]),
    .B2(_22232_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [38]),
    .C2(_23164_),
    .ZN(_25645_));
 NAND3_X2 _56877_ (.A1(_23215_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2635]),
    .A3(_23310_),
    .ZN(_25646_));
 OAI21_X4 _56878_ (.A(_25646_),
    .B1(_10888_),
    .B2(_21594_),
    .ZN(_25647_));
 AOI221_X2 _56879_ (.A(_25647_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1361]),
    .B2(_11054_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [577]),
    .C2(_11147_),
    .ZN(_25648_));
 NAND3_X1 _56880_ (.A1(_23242_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2978]),
    .A3(_22999_),
    .ZN(_25649_));
 NAND3_X1 _56881_ (.A1(_23390_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3125]),
    .A3(_23122_),
    .ZN(_25650_));
 NAND3_X1 _56882_ (.A1(_23303_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3027]),
    .A3(_23122_),
    .ZN(_25651_));
 NAND3_X1 _56883_ (.A1(_22967_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2782]),
    .A3(_23122_),
    .ZN(_25652_));
 AND4_X4 _56884_ (.A1(_25649_),
    .A2(_25650_),
    .A3(_25651_),
    .A4(_25652_),
    .ZN(_25653_));
 AND4_X2 _56885_ (.A1(_25642_),
    .A2(_25645_),
    .A3(_25648_),
    .A4(_25653_),
    .ZN(_25654_));
 AOI22_X4 _56886_ (.A1(_11196_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [185]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [332]),
    .B2(_22903_),
    .ZN(_25655_));
 NAND3_X2 _56887_ (.A1(_22998_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1067]),
    .A3(_23880_),
    .ZN(_25656_));
 OAI211_X4 _56888_ (.A(_25655_),
    .B(_25656_),
    .C1(_22405_),
    .C2(_11076_),
    .ZN(_25657_));
 AOI22_X4 _56889_ (.A1(_23267_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [822]),
    .B1(_23333_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1116]),
    .ZN(_25658_));
 NAND3_X2 _56890_ (.A1(_22968_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2390]),
    .A3(_23014_),
    .ZN(_25659_));
 OAI211_X4 _56891_ (.A(_25658_),
    .B(_25659_),
    .C1(_21671_),
    .C2(_10908_),
    .ZN(_25660_));
 AOI22_X2 _56892_ (.A1(_11153_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [528]),
    .B1(_11159_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [479]),
    .ZN(_25661_));
 NAND3_X2 _56893_ (.A1(_22975_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [675]),
    .A3(_23201_),
    .ZN(_25662_));
 OAI211_X4 _56894_ (.A(_25661_),
    .B(_25662_),
    .C1(_11121_),
    .C2(_22622_),
    .ZN(_25663_));
 NAND3_X1 _56895_ (.A1(_23200_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [969]),
    .A3(_22973_),
    .ZN(_25664_));
 NAND3_X2 _56896_ (.A1(_23271_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1018]),
    .A3(_23891_),
    .ZN(_25665_));
 NAND3_X4 _56897_ (.A1(_23839_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [626]),
    .A3(_23208_),
    .ZN(_25666_));
 NAND3_X2 _56898_ (.A1(_23207_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1214]),
    .A3(_23205_),
    .ZN(_25667_));
 NAND4_X4 _56899_ (.A1(_25664_),
    .A2(_25665_),
    .A3(_25666_),
    .A4(_25667_),
    .ZN(_25668_));
 NOR4_X4 _56900_ (.A1(_25657_),
    .A2(_25660_),
    .A3(_25663_),
    .A4(_25668_),
    .ZN(_25669_));
 NAND4_X1 _56901_ (.A1(_25623_),
    .A2(_25639_),
    .A3(_25654_),
    .A4(_25669_),
    .ZN(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [38]));
 AND3_X1 _56902_ (.A1(_23721_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [137]),
    .A3(_23643_),
    .ZN(_25670_));
 AOI221_X4 _56903_ (.A(_25670_),
    .B1(_11205_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [39]),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [186]),
    .C2(_11196_),
    .ZN(_25671_));
 NAND3_X1 _56904_ (.A1(_23215_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1068]),
    .A3(_23938_),
    .ZN(_25672_));
 OAI221_X2 _56905_ (.A(_25672_),
    .B1(_11086_),
    .B2(_22430_),
    .C1(_11076_),
    .C2(_22407_),
    .ZN(_25673_));
 AOI221_X4 _56906_ (.A(_25673_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1019]),
    .B2(_23104_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [872]),
    .C2(_22544_),
    .ZN(_25674_));
 AND3_X1 _56907_ (.A1(_22942_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [333]),
    .A3(_23159_),
    .ZN(_25675_));
 AOI221_X4 _56908_ (.A(_25675_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [284]),
    .B2(_22777_),
    .C1(_23615_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [382]),
    .ZN(_25676_));
 AOI22_X2 _56909_ (.A1(_23248_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [235]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [88]),
    .B2(_23490_),
    .ZN(_25677_));
 AND4_X4 _56910_ (.A1(_25671_),
    .A2(_25674_),
    .A3(_25676_),
    .A4(_25677_),
    .ZN(_25678_));
 NAND3_X1 _56911_ (.A1(_23215_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1852]),
    .A3(_10987_),
    .ZN(_25679_));
 OAI221_X2 _56912_ (.A(_25679_),
    .B1(_10994_),
    .B2(_22040_),
    .C1(_10984_),
    .C2(_21998_),
    .ZN(_25680_));
 AOI221_X4 _56913_ (.A(_25680_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1803]),
    .B2(_11002_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1656]),
    .C2(_23396_),
    .ZN(_25681_));
 NAND3_X1 _56914_ (.A1(_23245_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2342]),
    .A3(_10941_),
    .ZN(_25682_));
 NAND3_X1 _56915_ (.A1(_22241_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2244]),
    .A3(_10941_),
    .ZN(_25683_));
 NAND3_X1 _56916_ (.A1(_23367_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2195]),
    .A3(_23553_),
    .ZN(_25684_));
 NAND3_X1 _56917_ (.A1(_10818_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2293]),
    .A3(_23388_),
    .ZN(_25685_));
 AND4_X2 _56918_ (.A1(_25682_),
    .A2(_25683_),
    .A3(_25684_),
    .A4(_25685_),
    .ZN(_25686_));
 AND3_X1 _56919_ (.A1(_23173_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1705]),
    .A3(_23662_),
    .ZN(_25687_));
 AOI221_X4 _56920_ (.A(_25687_),
    .B1(_11025_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1607]),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1754]),
    .C2(_22078_),
    .ZN(_25688_));
 NAND3_X1 _56921_ (.A1(_10877_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1999]),
    .A3(_10939_),
    .ZN(_25689_));
 OAI21_X1 _56922_ (.A(_25689_),
    .B1(_10973_),
    .B2(_21957_),
    .ZN(_25690_));
 AOI221_X4 _56923_ (.A(_25690_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2146]),
    .B2(_10961_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2097]),
    .C2(_21900_),
    .ZN(_25691_));
 AND4_X4 _56924_ (.A1(_25681_),
    .A2(_25686_),
    .A3(_25688_),
    .A4(_25691_),
    .ZN(_25692_));
 NAND3_X1 _56925_ (.A1(_23309_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2587]),
    .A3(_23669_),
    .ZN(_25693_));
 OAI221_X2 _56926_ (.A(_25693_),
    .B1(_10897_),
    .B2(_21625_),
    .C1(_10888_),
    .C2(_21597_),
    .ZN(_25694_));
 AOI221_X2 _56927_ (.A(_25694_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2636]),
    .B2(_23627_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2440]),
    .C2(_10922_),
    .ZN(_25695_));
 NAND3_X1 _56928_ (.A1(_23434_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3028]),
    .A3(_23673_),
    .ZN(_25696_));
 AOI22_X1 _56929_ (.A1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2783]),
    .A2(_21289_),
    .B1(_22918_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2979]),
    .ZN(_25697_));
 NAND3_X1 _56930_ (.A1(_23240_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3077]),
    .A3(_23360_),
    .ZN(_25698_));
 NAND3_X1 _56931_ (.A1(_10804_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3126]),
    .A3(_22990_),
    .ZN(_25699_));
 AND4_X2 _56932_ (.A1(_25696_),
    .A2(_25697_),
    .A3(_25698_),
    .A4(_25699_),
    .ZN(_25700_));
 NAND3_X2 _56933_ (.A1(_22967_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2391]),
    .A3(_23304_),
    .ZN(_25701_));
 OAI221_X2 _56934_ (.A(_25701_),
    .B1(_10917_),
    .B2(_21734_),
    .C1(_10913_),
    .C2(_21700_),
    .ZN(_25702_));
 AND3_X1 _56935_ (.A1(_23035_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2832]),
    .A3(_23122_),
    .ZN(_25703_));
 AND3_X1 _56936_ (.A1(_22954_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2930]),
    .A3(_10789_),
    .ZN(_25704_));
 AND3_X1 _56937_ (.A1(_10857_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2881]),
    .A3(_10789_),
    .ZN(_25705_));
 NOR4_X1 _56938_ (.A1(_25702_),
    .A2(_25703_),
    .A3(_25704_),
    .A4(_25705_),
    .ZN(_25706_));
 AND3_X2 _56939_ (.A1(_25695_),
    .A2(_25700_),
    .A3(_25706_),
    .ZN(_25707_));
 NAND3_X1 _56940_ (.A1(_23385_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [676]),
    .A3(_23237_),
    .ZN(_25708_));
 AND3_X1 _56941_ (.A1(_10811_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [725]),
    .A3(_11123_),
    .ZN(_25709_));
 AOI221_X2 _56942_ (.A(_25709_),
    .B1(_11141_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [627]),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [774]),
    .C2(_22597_),
    .ZN(_25710_));
 AOI22_X2 _56943_ (.A1(_11147_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [578]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [529]),
    .B2(_23689_),
    .ZN(_25711_));
 AOI22_X4 _56944_ (.A1(_22733_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [431]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [480]),
    .B2(_11158_),
    .ZN(_25712_));
 AND4_X4 _56945_ (.A1(_25708_),
    .A2(_25710_),
    .A3(_25711_),
    .A4(_25712_),
    .ZN(_25713_));
 NAND3_X1 _56946_ (.A1(_22241_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1460]),
    .A3(_23693_),
    .ZN(_25714_));
 NAND3_X1 _56947_ (.A1(_23390_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1558]),
    .A3(_23608_),
    .ZN(_25715_));
 NAND3_X1 _56948_ (.A1(_23296_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1411]),
    .A3(_23608_),
    .ZN(_25716_));
 NAND3_X1 _56949_ (.A1(_10818_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1509]),
    .A3(_23608_),
    .ZN(_25717_));
 AND4_X4 _56950_ (.A1(_25714_),
    .A2(_25715_),
    .A3(_25716_),
    .A4(_25717_),
    .ZN(_25718_));
 AND3_X1 _56951_ (.A1(_23083_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [823]),
    .A3(_23460_),
    .ZN(_25719_));
 AOI221_X4 _56952_ (.A(_25719_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [921]),
    .B2(_11106_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [970]),
    .C2(_11100_),
    .ZN(_25720_));
 NAND3_X1 _56953_ (.A1(_23083_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1215]),
    .A3(_23701_),
    .ZN(_25721_));
 NAND3_X1 _56954_ (.A1(_23176_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1264]),
    .A3(_23701_),
    .ZN(_25722_));
 NAND2_X1 _56955_ (.A1(_25721_),
    .A2(_25722_),
    .ZN(_25723_));
 AOI221_X4 _56956_ (.A(_25723_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1313]),
    .B2(_11059_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1362]),
    .C2(_23748_),
    .ZN(_25724_));
 AND4_X4 _56957_ (.A1(_25713_),
    .A2(_25718_),
    .A3(_25720_),
    .A4(_25724_),
    .ZN(_25725_));
 NAND4_X4 _56958_ (.A1(_25678_),
    .A2(_25692_),
    .A3(_25707_),
    .A4(_25725_),
    .ZN(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [39]));
 OAI22_X4 _56959_ (.A1(_22277_),
    .A2(_11051_),
    .B1(_11070_),
    .B2(_22383_),
    .ZN(_25726_));
 OAI22_X4 _56960_ (.A1(_11032_),
    .A2(_22207_),
    .B1(_22228_),
    .B2(_11042_),
    .ZN(_25727_));
 AOI211_X2 _56961_ (.A(_25726_),
    .B(_25727_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1461]),
    .C2(_23326_),
    .ZN(_25728_));
 NAND3_X1 _56962_ (.A1(_23217_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1167]),
    .A3(_23938_),
    .ZN(_25729_));
 OAI221_X2 _56963_ (.A(_25729_),
    .B1(_11086_),
    .B2(_22432_),
    .C1(_11095_),
    .C2(_22491_),
    .ZN(_25730_));
 AOI221_X2 _56964_ (.A(_25730_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1069]),
    .B2(_22435_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [873]),
    .C2(_22544_),
    .ZN(_25731_));
 AND3_X2 _56965_ (.A1(_23382_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [824]),
    .A3(_23494_),
    .ZN(_25732_));
 AOI221_X2 _56966_ (.A(_25732_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [922]),
    .B2(_23265_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [971]),
    .C2(_23047_),
    .ZN(_25733_));
 AND3_X1 _56967_ (.A1(_23806_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1265]),
    .A3(_23848_),
    .ZN(_25734_));
 AOI221_X4 _56968_ (.A(_25734_),
    .B1(_11060_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1314]),
    .C1(_22282_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1363]),
    .ZN(_25735_));
 AND4_X4 _56969_ (.A1(_25728_),
    .A2(_25731_),
    .A3(_25733_),
    .A4(_25735_),
    .ZN(_25736_));
 AND3_X1 _56970_ (.A1(_22953_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2931]),
    .A3(_23498_),
    .ZN(_25737_));
 AOI221_X4 _56971_ (.A(_25737_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2882]),
    .B2(_10851_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2833]),
    .C2(_21536_),
    .ZN(_25738_));
 NAND3_X1 _56972_ (.A1(_23284_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2343]),
    .A3(_23657_),
    .ZN(_25739_));
 NAND3_X1 _56973_ (.A1(_23751_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2294]),
    .A3(_23657_),
    .ZN(_25740_));
 NAND2_X1 _56974_ (.A1(_25739_),
    .A2(_25740_),
    .ZN(_25741_));
 AOI221_X2 _56975_ (.A(_25741_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2245]),
    .B2(_10950_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2196]),
    .C2(_23660_),
    .ZN(_25742_));
 NAND3_X1 _56976_ (.A1(_23339_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2980]),
    .A3(_22990_),
    .ZN(_25743_));
 AOI22_X2 _56977_ (.A1(_23224_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3127]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3078]),
    .B2(_23225_),
    .ZN(_25744_));
 NAND3_X1 _56978_ (.A1(_10879_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2784]),
    .A3(_22999_),
    .ZN(_25745_));
 NAND3_X1 _56979_ (.A1(_23757_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3029]),
    .A3(_23122_),
    .ZN(_25746_));
 AND4_X4 _56980_ (.A1(_25743_),
    .A2(_25744_),
    .A3(_25745_),
    .A4(_25746_),
    .ZN(_25747_));
 NAND3_X1 _56981_ (.A1(_23230_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2000]),
    .A3(_22962_),
    .ZN(_25748_));
 NAND3_X1 _56982_ (.A1(_23176_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2049]),
    .A3(_23169_),
    .ZN(_25749_));
 NAND2_X1 _56983_ (.A1(_25748_),
    .A2(_25749_),
    .ZN(_25750_));
 AOI221_X4 _56984_ (.A(_25750_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2098]),
    .B2(_10968_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2147]),
    .C2(_23736_),
    .ZN(_25751_));
 AND4_X2 _56985_ (.A1(_25738_),
    .A2(net18),
    .A3(_25747_),
    .A4(_25751_),
    .ZN(_25752_));
 AND3_X1 _56986_ (.A1(_23382_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [432]),
    .A3(_23512_),
    .ZN(_25753_));
 AOI221_X4 _56987_ (.A(_25753_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [530]),
    .B2(_11152_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [579]),
    .C2(_11147_),
    .ZN(_25754_));
 NAND3_X1 _56988_ (.A1(_23339_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [236]),
    .A3(_23246_),
    .ZN(_25755_));
 AND3_X1 _56989_ (.A1(_10901_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [285]),
    .A3(_11185_),
    .ZN(_25756_));
 AOI221_X2 _56990_ (.A(_25756_),
    .B1(_11181_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [334]),
    .C1(_11170_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [383]),
    .ZN(_25757_));
 AOI22_X2 _56991_ (.A1(_22806_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [187]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [138]),
    .B2(_23453_),
    .ZN(_25758_));
 AOI22_X2 _56992_ (.A1(_23164_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [40]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [89]),
    .B2(_11211_),
    .ZN(_25759_));
 AND4_X4 _56993_ (.A1(_25755_),
    .A2(_25757_),
    .A3(_25758_),
    .A4(_25759_),
    .ZN(_25760_));
 AND3_X1 _56994_ (.A1(_23524_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [726]),
    .A3(_23255_),
    .ZN(_25761_));
 AOI221_X4 _56995_ (.A(_25761_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [677]),
    .B2(_22642_),
    .C1(_22597_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [775]),
    .ZN(_25762_));
 AOI22_X2 _56996_ (.A1(_23106_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [628]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [481]),
    .B2(_11159_),
    .ZN(_25763_));
 AND4_X4 _56997_ (.A1(_25754_),
    .A2(_25760_),
    .A3(_25762_),
    .A4(_25763_),
    .ZN(_25764_));
 AND3_X1 _56998_ (.A1(_23751_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1902]),
    .A3(_23519_),
    .ZN(_25765_));
 AOI221_X4 _56999_ (.A(_25765_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1853]),
    .B2(_22044_),
    .C1(_23584_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1951]),
    .ZN(_25766_));
 NAND3_X1 _57000_ (.A1(_22987_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2539]),
    .A3(_10892_),
    .ZN(_25767_));
 AOI22_X1 _57001_ (.A1(_10929_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2392]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2441]),
    .B2(_23301_),
    .ZN(_25768_));
 NAND3_X1 _57002_ (.A1(_22523_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2490]),
    .A3(_23119_),
    .ZN(_25769_));
 NAND3_X1 _57003_ (.A1(_23757_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2637]),
    .A3(_23119_),
    .ZN(_25770_));
 AND4_X1 _57004_ (.A1(_25767_),
    .A2(_25768_),
    .A3(_25769_),
    .A4(_25770_),
    .ZN(_25771_));
 AOI22_X2 _57005_ (.A1(_23290_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1755]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1706]),
    .B2(_22105_),
    .ZN(_25772_));
 NAND3_X1 _57006_ (.A1(_23339_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1804]),
    .A3(_23393_),
    .ZN(_25773_));
 AOI22_X2 _57007_ (.A1(_23595_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1608]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1657]),
    .B2(_23396_),
    .ZN(_25774_));
 AND3_X4 _57008_ (.A1(_25772_),
    .A2(_25773_),
    .A3(_25774_),
    .ZN(_25775_));
 AND3_X1 _57009_ (.A1(_23309_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2588]),
    .A3(_23310_),
    .ZN(_25776_));
 AOI221_X4 _57010_ (.A(_25776_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2686]),
    .B2(_21600_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2735]),
    .C2(_21573_),
    .ZN(_25777_));
 AND4_X2 _57011_ (.A1(_25766_),
    .A2(_25771_),
    .A3(_25775_),
    .A4(_25777_),
    .ZN(_25778_));
 NAND4_X2 _57012_ (.A1(_25736_),
    .A2(_25752_),
    .A3(_25764_),
    .A4(_25778_),
    .ZN(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [40]));
 NAND3_X1 _57013_ (.A1(_22897_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [776]),
    .A3(_23055_),
    .ZN(_25779_));
 NAND3_X4 _57014_ (.A1(_22907_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [433]),
    .A3(_23504_),
    .ZN(_25780_));
 NAND2_X1 _57015_ (.A1(_25779_),
    .A2(_25780_),
    .ZN(_25781_));
 AOI221_X2 _57016_ (.A(_25781_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [678]),
    .B2(_23107_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [629]),
    .C2(_23106_),
    .ZN(_25782_));
 NAND3_X4 _57017_ (.A1(_23166_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [580]),
    .A3(_23161_),
    .ZN(_25783_));
 OAI21_X4 _57018_ (.A(_25783_),
    .B1(_10917_),
    .B2(_21736_),
    .ZN(_25784_));
 AOI221_X4 _57019_ (.A(_25784_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2148]),
    .B2(_23736_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2099]),
    .C2(_21900_),
    .ZN(_25785_));
 NAND3_X1 _57020_ (.A1(_23982_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [531]),
    .A3(_23237_),
    .ZN(_25786_));
 NAND3_X1 _57021_ (.A1(_23240_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [727]),
    .A3(_11126_),
    .ZN(_25787_));
 NAND3_X4 _57022_ (.A1(_22997_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3030]),
    .A3(_22999_),
    .ZN(_25788_));
 NAND3_X1 _57023_ (.A1(_23113_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [482]),
    .A3(_23346_),
    .ZN(_25789_));
 AND4_X4 _57024_ (.A1(_25786_),
    .A2(_25787_),
    .A3(_25788_),
    .A4(_25789_),
    .ZN(_25790_));
 NAND3_X2 _57025_ (.A1(_23509_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1756]),
    .A3(_22921_),
    .ZN(_25791_));
 NAND3_X2 _57026_ (.A1(_23806_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2050]),
    .A3(_23657_),
    .ZN(_25792_));
 NAND2_X4 _57027_ (.A1(_25791_),
    .A2(_25792_),
    .ZN(_25793_));
 AOI221_X4 _57028_ (.A(_25793_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2393]),
    .B2(_10928_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1609]),
    .C2(_23395_),
    .ZN(_25794_));
 AND4_X1 _57029_ (.A1(net17),
    .A2(_25785_),
    .A3(_25790_),
    .A4(_25794_),
    .ZN(_25795_));
 NAND3_X1 _57030_ (.A1(_23810_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2736]),
    .A3(_23012_),
    .ZN(_25796_));
 OAI21_X1 _57031_ (.A(_25796_),
    .B1(_10897_),
    .B2(_21628_),
    .ZN(_25797_));
 AOI221_X2 _57032_ (.A(_25797_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2638]),
    .B2(_10902_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2246]),
    .C2(_10950_),
    .ZN(_25798_));
 NAND3_X1 _57033_ (.A1(_10778_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [188]),
    .A3(_22937_),
    .ZN(_25799_));
 OAI21_X2 _57034_ (.A(_25799_),
    .B1(_11201_),
    .B2(_22857_),
    .ZN(_25800_));
 AOI221_X4 _57035_ (.A(_25800_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2785]),
    .B2(_21289_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3079]),
    .C2(_23225_),
    .ZN(_25801_));
 NAND3_X2 _57036_ (.A1(_23518_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2197]),
    .A3(_23231_),
    .ZN(_25802_));
 NAND3_X4 _57037_ (.A1(_23518_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2589]),
    .A3(_23012_),
    .ZN(_25803_));
 NAND2_X4 _57038_ (.A1(_25802_),
    .A2(_25803_),
    .ZN(_25804_));
 AOI221_X4 _57039_ (.A(_25804_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1511]),
    .B2(_22210_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1462]),
    .C2(_23326_),
    .ZN(_25805_));
 NAND3_X1 _57040_ (.A1(_10856_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2883]),
    .A3(_23794_),
    .ZN(_25806_));
 NAND3_X1 _57041_ (.A1(_23176_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2834]),
    .A3(_23174_),
    .ZN(_25807_));
 NAND2_X2 _57042_ (.A1(_25806_),
    .A2(_25807_),
    .ZN(_25808_));
 AOI221_X4 _57043_ (.A(_25808_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1707]),
    .B2(_11012_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2981]),
    .C2(_22918_),
    .ZN(_25809_));
 AND4_X2 _57044_ (.A1(_25798_),
    .A2(_25801_),
    .A3(_25805_),
    .A4(_25809_),
    .ZN(_25810_));
 NAND3_X4 _57045_ (.A1(_23492_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2344]),
    .A3(_22913_),
    .ZN(_25811_));
 NAND3_X2 _57046_ (.A1(_23721_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [923]),
    .A3(_23494_),
    .ZN(_25812_));
 NAND2_X4 _57047_ (.A1(_25811_),
    .A2(_25812_),
    .ZN(_25813_));
 AOI221_X2 _57048_ (.A(_25813_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1364]),
    .B2(_23748_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1266]),
    .C2(_23048_),
    .ZN(_25814_));
 NAND3_X1 _57049_ (.A1(_23158_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [972]),
    .A3(_23804_),
    .ZN(_25815_));
 NAND3_X1 _57050_ (.A1(_23733_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [874]),
    .A3(_23804_),
    .ZN(_25816_));
 NAND2_X1 _57051_ (.A1(_25815_),
    .A2(_25816_),
    .ZN(_25817_));
 AOI221_X4 _57052_ (.A(_25817_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1070]),
    .B2(_11090_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [825]),
    .C2(_11114_),
    .ZN(_25818_));
 NAND3_X1 _57053_ (.A1(_23810_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1952]),
    .A3(_23662_),
    .ZN(_25819_));
 NAND3_X2 _57054_ (.A1(_23168_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1854]),
    .A3(_23662_),
    .ZN(_25820_));
 NAND2_X4 _57055_ (.A1(_25819_),
    .A2(_25820_),
    .ZN(_25821_));
 AOI221_X2 _57056_ (.A(_25821_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1658]),
    .B2(_11019_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1315]),
    .C2(_11060_),
    .ZN(_25822_));
 NAND3_X1 _57057_ (.A1(_23459_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [384]),
    .A3(_23258_),
    .ZN(_25823_));
 NAND3_X4 _57058_ (.A1(_23408_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1903]),
    .A3(_23402_),
    .ZN(_25824_));
 NAND2_X1 _57059_ (.A1(_25823_),
    .A2(_25824_),
    .ZN(_25825_));
 AOI221_X2 _57060_ (.A(_25825_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1217]),
    .B2(_11069_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [286]),
    .C2(_23446_),
    .ZN(_25826_));
 AND4_X4 _57061_ (.A1(net13),
    .A2(_25818_),
    .A3(_25822_),
    .A4(_25826_),
    .ZN(_25827_));
 AND3_X1 _57062_ (.A1(_10803_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1168]),
    .A3(_11080_),
    .ZN(_25828_));
 AOI21_X4 _57063_ (.A(_25828_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1119]),
    .B2(_23333_),
    .ZN(_25829_));
 OAI221_X2 _57064_ (.A(_25829_),
    .B1(_21409_),
    .B2(_10801_),
    .C1(_21501_),
    .C2(_10774_),
    .ZN(_25830_));
 NAND3_X4 _57065_ (.A1(_23054_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1560]),
    .A3(_22945_),
    .ZN(_25831_));
 NAND3_X4 _57066_ (.A1(_23127_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [335]),
    .A3(_11176_),
    .ZN(_25832_));
 NAND3_X2 _57067_ (.A1(_23062_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2442]),
    .A3(_23068_),
    .ZN(_25833_));
 NAND3_X4 _57068_ (.A1(_23192_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1413]),
    .A3(_23566_),
    .ZN(_25834_));
 NAND4_X4 _57069_ (.A1(_25831_),
    .A2(_25832_),
    .A3(_25833_),
    .A4(_25834_),
    .ZN(_25835_));
 NAND3_X2 _57070_ (.A1(_22955_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2540]),
    .A3(_23134_),
    .ZN(_25836_));
 NAND3_X2 _57071_ (.A1(_22972_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2295]),
    .A3(_22964_),
    .ZN(_25837_));
 NAND3_X2 _57072_ (.A1(_23271_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1805]),
    .A3(_23146_),
    .ZN(_25838_));
 NAND3_X2 _57073_ (.A1(_23085_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2001]),
    .A3(_23081_),
    .ZN(_25839_));
 NAND4_X4 _57074_ (.A1(_25836_),
    .A2(_25837_),
    .A3(_25838_),
    .A4(_25839_),
    .ZN(_25840_));
 NAND3_X1 _57075_ (.A1(_10844_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [237]),
    .A3(_23835_),
    .ZN(_25841_));
 NAND3_X1 _57076_ (.A1(_23837_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [41]),
    .A3(_23196_),
    .ZN(_25842_));
 NAND3_X4 _57077_ (.A1(_23839_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1021]),
    .A3(_23547_),
    .ZN(_25843_));
 NAND3_X1 _57078_ (.A1(_23426_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [90]),
    .A3(_23086_),
    .ZN(_25844_));
 NAND4_X2 _57079_ (.A1(_25841_),
    .A2(_25842_),
    .A3(_25843_),
    .A4(_25844_),
    .ZN(_25845_));
 NOR4_X1 _57080_ (.A1(_25830_),
    .A2(_25835_),
    .A3(_25840_),
    .A4(_25845_),
    .ZN(_25846_));
 NAND4_X1 _57081_ (.A1(_25795_),
    .A2(_25810_),
    .A3(_25827_),
    .A4(_25846_),
    .ZN(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [41]));
 NAND3_X2 _57082_ (.A1(_22897_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [777]),
    .A3(_23055_),
    .ZN(_25847_));
 NAND3_X2 _57083_ (.A1(_10829_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [679]),
    .A3(_23504_),
    .ZN(_25848_));
 NAND2_X4 _57084_ (.A1(_25847_),
    .A2(_25848_),
    .ZN(_25849_));
 AOI221_X4 _57085_ (.A(_25849_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1463]),
    .B2(_22232_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1218]),
    .C2(_23103_),
    .ZN(_25850_));
 NAND3_X1 _57086_ (.A1(_23166_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1365]),
    .A3(_23848_),
    .ZN(_25851_));
 OAI21_X2 _57087_ (.A(_25851_),
    .B1(_11051_),
    .B2(_22279_),
    .ZN(_25852_));
 AOI221_X4 _57088_ (.A(_25852_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1561]),
    .B2(_11031_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1512]),
    .C2(_23095_),
    .ZN(_25853_));
 NAND3_X1 _57089_ (.A1(_23733_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2443]),
    .A3(_23669_),
    .ZN(_25854_));
 OAI21_X1 _57090_ (.A(_25854_),
    .B1(_10903_),
    .B2(_21651_),
    .ZN(_25855_));
 AOI221_X4 _57091_ (.A(_25855_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2492]),
    .B2(_10916_),
    .C1(net1391),
    .C2(_23092_),
    .ZN(_25856_));
 NAND3_X4 _57092_ (.A1(_22915_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [483]),
    .A3(_23510_),
    .ZN(_25857_));
 NAND3_X1 _57093_ (.A1(_23806_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2835]),
    .A3(_23794_),
    .ZN(_25858_));
 NAND2_X1 _57094_ (.A1(_25857_),
    .A2(_25858_),
    .ZN(_25859_));
 AOI221_X4 _57095_ (.A(_25859_),
    .B1(_23300_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2394]),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2933]),
    .C2(_21466_),
    .ZN(_25860_));
 AND4_X1 _57096_ (.A1(_25850_),
    .A2(_25853_),
    .A3(_25856_),
    .A4(_25860_),
    .ZN(_25861_));
 NAND3_X2 _57097_ (.A1(_23810_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1953]),
    .A3(_23519_),
    .ZN(_25862_));
 OAI21_X4 _57098_ (.A(_25862_),
    .B1(_10994_),
    .B2(_22043_),
    .ZN(_25863_));
 AOI221_X2 _57099_ (.A(_25863_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1806]),
    .B2(_11002_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1267]),
    .C2(_23048_),
    .ZN(_25864_));
 NAND3_X2 _57100_ (.A1(_23509_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [581]),
    .A3(_23510_),
    .ZN(_25865_));
 NAND3_X2 _57101_ (.A1(_23518_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [630]),
    .A3(_23512_),
    .ZN(_25866_));
 NAND2_X4 _57102_ (.A1(_25865_),
    .A2(_25866_),
    .ZN(_25867_));
 AOI221_X4 _57103_ (.A(_25867_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1855]),
    .B2(_22044_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1316]),
    .C2(_23262_),
    .ZN(_25868_));
 NAND3_X1 _57104_ (.A1(_23487_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2737]),
    .A3(_23481_),
    .ZN(_25869_));
 NAND3_X4 _57105_ (.A1(_23230_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2786]),
    .A3(_23174_),
    .ZN(_25870_));
 NAND2_X1 _57106_ (.A1(_25869_),
    .A2(_25870_),
    .ZN(_25871_));
 AOI221_X2 _57107_ (.A(_25871_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2688]),
    .B2(_21601_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2100]),
    .C2(_21900_),
    .ZN(_25872_));
 NAND3_X1 _57108_ (.A1(_23524_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3080]),
    .A3(_23794_),
    .ZN(_25873_));
 NAND3_X1 _57109_ (.A1(_23168_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3031]),
    .A3(_23174_),
    .ZN(_25874_));
 NAND2_X2 _57110_ (.A1(_25873_),
    .A2(_25874_),
    .ZN(_25875_));
 AOI221_X4 _57111_ (.A(_25875_),
    .B1(_11190_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [238]),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [385]),
    .C2(_11170_),
    .ZN(_25876_));
 AND4_X2 _57112_ (.A1(_25864_),
    .A2(_25868_),
    .A3(_25872_),
    .A4(_25876_),
    .ZN(_25877_));
 AOI22_X4 _57113_ (.A1(_23331_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1169]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1708]),
    .B2(_23591_),
    .ZN(_25878_));
 NAND3_X2 _57114_ (.A1(_22944_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2296]),
    .A3(_23554_),
    .ZN(_25879_));
 OAI211_X4 _57115_ (.A(_25878_),
    .B(_25879_),
    .C1(_21814_),
    .C2(_10937_),
    .ZN(_25880_));
 NAND3_X1 _57116_ (.A1(_23004_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [973]),
    .A3(_23880_),
    .ZN(_25881_));
 NAND3_X2 _57117_ (.A1(_23377_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [875]),
    .A3(_23882_),
    .ZN(_25882_));
 NAND3_X2 _57118_ (.A1(_10858_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [924]),
    .A3(_23882_),
    .ZN(_25883_));
 NAND3_X2 _57119_ (.A1(_23133_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [826]),
    .A3(_22970_),
    .ZN(_25884_));
 NAND4_X4 _57120_ (.A1(_25881_),
    .A2(_25882_),
    .A3(_25883_),
    .A4(_25884_),
    .ZN(_25885_));
 NAND3_X4 _57121_ (.A1(_23067_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3129]),
    .A3(_23033_),
    .ZN(_25886_));
 NAND3_X1 _57122_ (.A1(_22972_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1120]),
    .A3(_22973_),
    .ZN(_25887_));
 NAND3_X2 _57123_ (.A1(_23276_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1022]),
    .A3(_22976_),
    .ZN(_25888_));
 NAND3_X2 _57124_ (.A1(_23071_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1071]),
    .A3(_23891_),
    .ZN(_25889_));
 NAND4_X4 _57125_ (.A1(_25886_),
    .A2(_25887_),
    .A3(_25888_),
    .A4(_25889_),
    .ZN(_25890_));
 NAND3_X2 _57126_ (.A1(_22955_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2149]),
    .A3(_23894_),
    .ZN(_25891_));
 NAND3_X2 _57127_ (.A1(_23271_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2198]),
    .A3(_23832_),
    .ZN(_25892_));
 NAND3_X1 _57128_ (.A1(_23080_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2247]),
    .A3(_23081_),
    .ZN(_25893_));
 NAND3_X2 _57129_ (.A1(_23426_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1659]),
    .A3(_23576_),
    .ZN(_25894_));
 NAND4_X4 _57130_ (.A1(_25891_),
    .A2(_25892_),
    .A3(_25893_),
    .A4(_25894_),
    .ZN(_25895_));
 NOR4_X1 _57131_ (.A1(_25880_),
    .A2(_25885_),
    .A3(_25890_),
    .A4(_25895_),
    .ZN(_25896_));
 AND3_X1 _57132_ (.A1(_23041_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [91]),
    .A3(_22938_),
    .ZN(_25897_));
 AOI21_X4 _57133_ (.A(_25897_),
    .B1(_11206_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [42]),
    .ZN(_25898_));
 OAI221_X2 _57134_ (.A(_25898_),
    .B1(_10840_),
    .B2(_21463_),
    .C1(_21675_),
    .C2(_10908_),
    .ZN(_25899_));
 AOI22_X4 _57135_ (.A1(_22903_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [336]),
    .B1(_23446_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [287]),
    .ZN(_25900_));
 NAND3_X2 _57136_ (.A1(_23016_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [140]),
    .A3(_23187_),
    .ZN(_25901_));
 OAI211_X4 _57137_ (.A(_25900_),
    .B(_25901_),
    .C1(_11197_),
    .C2(_22826_),
    .ZN(_25902_));
 NAND3_X4 _57138_ (.A1(_23133_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1610]),
    .A3(_22956_),
    .ZN(_25903_));
 NAND3_X2 _57139_ (.A1(_23194_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [434]),
    .A3(_23201_),
    .ZN(_25904_));
 NAND3_X4 _57140_ (.A1(_23078_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2884]),
    .A3(_23037_),
    .ZN(_25905_));
 NAND3_X4 _57141_ (.A1(_23039_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [532]),
    .A3(_23208_),
    .ZN(_25906_));
 NAND4_X4 _57142_ (.A1(_25903_),
    .A2(_25904_),
    .A3(_25905_),
    .A4(_25906_),
    .ZN(_25907_));
 NAND3_X2 _57143_ (.A1(_23200_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1757]),
    .A3(_23141_),
    .ZN(_25908_));
 NAND3_X4 _57144_ (.A1(_23421_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2541]),
    .A3(_23029_),
    .ZN(_25909_));
 NAND3_X2 _57145_ (.A1(_23042_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2051]),
    .A3(_23081_),
    .ZN(_25910_));
 NAND3_X2 _57146_ (.A1(_23207_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2002]),
    .A3(_23600_),
    .ZN(_25911_));
 NAND4_X4 _57147_ (.A1(_25908_),
    .A2(_25909_),
    .A3(_25910_),
    .A4(_25911_),
    .ZN(_25912_));
 NOR4_X2 _57148_ (.A1(_25899_),
    .A2(_25902_),
    .A3(_25907_),
    .A4(_25912_),
    .ZN(_25913_));
 NAND4_X1 _57149_ (.A1(_25861_),
    .A2(_25877_),
    .A3(_25896_),
    .A4(_25913_),
    .ZN(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [42]));
 NAND3_X1 _57150_ (.A1(_23438_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1464]),
    .A3(_23931_),
    .ZN(_25914_));
 AOI22_X1 _57151_ (.A1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1415]),
    .A2(_23094_),
    .B1(_23103_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1219]),
    .ZN(_25915_));
 NAND3_X1 _57152_ (.A1(_24262_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1562]),
    .A3(_23931_),
    .ZN(_25916_));
 NAND3_X1 _57153_ (.A1(_24186_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1513]),
    .A3(_23412_),
    .ZN(_25917_));
 AND4_X4 _57154_ (.A1(_25914_),
    .A2(_25915_),
    .A3(_25916_),
    .A4(_25917_),
    .ZN(_25918_));
 NAND3_X1 _57155_ (.A1(_10842_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1023]),
    .A3(_23938_),
    .ZN(_25919_));
 OAI221_X2 _57156_ (.A(_25919_),
    .B1(_11086_),
    .B2(_22434_),
    .C1(_11076_),
    .C2(_22409_),
    .ZN(_25920_));
 AOI221_X4 _57157_ (.A(_25920_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1072]),
    .B2(_22435_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [827]),
    .C2(_23267_),
    .ZN(_25921_));
 AND3_X1 _57158_ (.A1(_23158_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [974]),
    .A3(_23494_),
    .ZN(_25922_));
 AOI221_X4 _57159_ (.A(_25922_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [925]),
    .B2(_23265_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [876]),
    .C2(_22544_),
    .ZN(_25923_));
 AND3_X1 _57160_ (.A1(_23806_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1268]),
    .A3(_23848_),
    .ZN(_25924_));
 AOI221_X4 _57161_ (.A(_25924_),
    .B1(_11060_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1317]),
    .C1(_22282_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1366]),
    .ZN(_25925_));
 AND4_X4 _57162_ (.A1(_25918_),
    .A2(_25921_),
    .A3(_25923_),
    .A4(_25925_),
    .ZN(_25926_));
 AND3_X1 _57163_ (.A1(_22915_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2052]),
    .A3(_22913_),
    .ZN(_25927_));
 AOI221_X4 _57164_ (.A(_25927_),
    .B1(_21900_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2101]),
    .C1(_10962_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2150]),
    .ZN(_25928_));
 NAND3_X1 _57165_ (.A1(_10798_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2738]),
    .A3(_10890_),
    .ZN(_25929_));
 OAI221_X2 _57166_ (.A(_25929_),
    .B1(_10897_),
    .B2(_21631_),
    .C1(_10908_),
    .C2(_21677_),
    .ZN(_25930_));
 AOI221_X1 _57167_ (.A(_25930_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2640]),
    .B2(_10902_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2395]),
    .C2(_23300_),
    .ZN(_25931_));
 AND3_X1 _57168_ (.A1(_23168_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2248]),
    .A3(_22962_),
    .ZN(_25932_));
 AOI221_X4 _57169_ (.A(_25932_),
    .B1(_21816_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2297]),
    .C1(_23097_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2346]),
    .ZN(_25933_));
 AOI22_X4 _57170_ (.A1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2199]),
    .A2(_10956_),
    .B1(_23485_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2003]),
    .ZN(_25934_));
 AND4_X2 _57171_ (.A1(_25928_),
    .A2(_25931_),
    .A3(_25933_),
    .A4(_25934_),
    .ZN(_25935_));
 AND3_X1 _57172_ (.A1(_22942_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [729]),
    .A3(_23512_),
    .ZN(_25936_));
 AOI221_X4 _57173_ (.A(_25936_),
    .B1(_23515_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [631]),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [778]),
    .C2(_23638_),
    .ZN(_25937_));
 NAND3_X2 _57174_ (.A1(_10779_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [190]),
    .A3(_22938_),
    .ZN(_25938_));
 OAI21_X4 _57175_ (.A(_25938_),
    .B1(_11201_),
    .B2(_22859_),
    .ZN(_25939_));
 NAND3_X2 _57176_ (.A1(_22522_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [533]),
    .A3(_11125_),
    .ZN(_25940_));
 NAND3_X2 _57177_ (.A1(_23041_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [484]),
    .A3(_11125_),
    .ZN(_25941_));
 OAI211_X4 _57178_ (.A(_25940_),
    .B(_25941_),
    .C1(_11148_),
    .C2(_22696_),
    .ZN(_25942_));
 AOI211_X1 _57179_ (.A(_25939_),
    .B(_25942_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [43]),
    .C2(_11206_),
    .ZN(_25943_));
 OAI22_X4 _57180_ (.A1(_11191_),
    .A2(_22805_),
    .B1(_22893_),
    .B2(_11212_),
    .ZN(_25944_));
 OAI22_X2 _57181_ (.A1(_11171_),
    .A2(_22757_),
    .B1(_22776_),
    .B2(_11182_),
    .ZN(_25945_));
 AOI211_X2 _57182_ (.A(_25944_),
    .B(_25945_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [288]),
    .C2(_23446_),
    .ZN(_25946_));
 AOI22_X4 _57183_ (.A1(_23610_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [435]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [680]),
    .B2(_23107_),
    .ZN(_25947_));
 AND4_X4 _57184_ (.A1(_25937_),
    .A2(_25943_),
    .A3(_25946_),
    .A4(_25947_),
    .ZN(_25948_));
 AND3_X1 _57185_ (.A1(_23751_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1905]),
    .A3(_23519_),
    .ZN(_25949_));
 AOI221_X4 _57186_ (.A(_25949_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1856]),
    .B2(_22044_),
    .C1(_23584_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1954]),
    .ZN(_25950_));
 OAI22_X2 _57187_ (.A1(_11026_),
    .A2(_22183_),
    .B1(_22156_),
    .B2(_11020_),
    .ZN(_25951_));
 OAI22_X2 _57188_ (.A1(_11009_),
    .A2(_22103_),
    .B1(_22131_),
    .B2(_11013_),
    .ZN(_25952_));
 AOI211_X2 _57189_ (.A(_25951_),
    .B(_25952_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1807]),
    .C2(_11003_),
    .ZN(_25953_));
 NAND3_X1 _57190_ (.A1(_23245_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3130]),
    .A3(_23360_),
    .ZN(_25954_));
 NAND3_X1 _57191_ (.A1(_23240_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3081]),
    .A3(_22990_),
    .ZN(_25955_));
 NAND2_X2 _57192_ (.A1(_25954_),
    .A2(_25955_),
    .ZN(_25956_));
 AND3_X1 _57193_ (.A1(_22932_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2983]),
    .A3(_23122_),
    .ZN(_25957_));
 AND3_X1 _57194_ (.A1(_23303_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3032]),
    .A3(_10789_),
    .ZN(_25958_));
 NOR3_X4 _57195_ (.A1(_25956_),
    .A2(_25957_),
    .A3(_25958_),
    .ZN(_25959_));
 OAI22_X2 _57196_ (.A1(_10913_),
    .A2(_21702_),
    .B1(_21740_),
    .B2(_10917_),
    .ZN(_25960_));
 NAND3_X1 _57197_ (.A1(_22954_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2934]),
    .A3(_22928_),
    .ZN(_25961_));
 OAI21_X2 _57198_ (.A(_25961_),
    .B1(_10852_),
    .B2(_21535_),
    .ZN(_25962_));
 NAND3_X1 _57199_ (.A1(_23084_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2787]),
    .A3(_22928_),
    .ZN(_25963_));
 OAI21_X2 _57200_ (.A(_25963_),
    .B1(_10864_),
    .B2(_21568_),
    .ZN(_25964_));
 AND3_X1 _57201_ (.A1(_23041_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2444]),
    .A3(_10891_),
    .ZN(_25965_));
 NOR4_X1 _57202_ (.A1(_25960_),
    .A2(_25962_),
    .A3(_25964_),
    .A4(_25965_),
    .ZN(_25966_));
 AND4_X1 _57203_ (.A1(_25950_),
    .A2(net12),
    .A3(_25959_),
    .A4(_25966_),
    .ZN(_25967_));
 NAND4_X2 _57204_ (.A1(_25926_),
    .A2(_25935_),
    .A3(_25948_),
    .A4(_25967_),
    .ZN(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [43]));
 AND3_X1 _57205_ (.A1(_23721_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2886]),
    .A3(_10788_),
    .ZN(_25968_));
 AOI221_X4 _57206_ (.A(_25968_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2837]),
    .B2(_21536_),
    .C1(_23213_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2935]),
    .ZN(_25969_));
 NAND3_X1 _57207_ (.A1(_24186_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3082]),
    .A3(_23673_),
    .ZN(_25970_));
 AOI22_X4 _57208_ (.A1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2788]),
    .A2(_21289_),
    .B1(_22918_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2984]),
    .ZN(_25971_));
 NAND3_X1 _57209_ (.A1(_10804_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3131]),
    .A3(_22990_),
    .ZN(_25972_));
 NAND3_X1 _57210_ (.A1(_22241_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3033]),
    .A3(_22990_),
    .ZN(_25973_));
 AND4_X2 _57211_ (.A1(_25970_),
    .A2(_25971_),
    .A3(_25972_),
    .A4(_25973_),
    .ZN(_25974_));
 AND3_X1 _57212_ (.A1(_23382_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2004]),
    .A3(_23657_),
    .ZN(_25975_));
 AOI221_X4 _57213_ (.A(_25975_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2102]),
    .B2(_22910_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2151]),
    .C2(_10962_),
    .ZN(_25976_));
 NAND3_X1 _57214_ (.A1(_24186_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2298]),
    .A3(_23600_),
    .ZN(_25977_));
 AOI22_X2 _57215_ (.A1(_10956_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2200]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2053]),
    .B2(_21937_),
    .ZN(_25978_));
 NAND3_X1 _57216_ (.A1(_22997_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2249]),
    .A3(_23553_),
    .ZN(_25979_));
 NAND3_X1 _57217_ (.A1(_10804_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2347]),
    .A3(_23388_),
    .ZN(_25980_));
 AND4_X4 _57218_ (.A1(_25977_),
    .A2(_25978_),
    .A3(_25979_),
    .A4(_25980_),
    .ZN(_25981_));
 AND4_X2 _57219_ (.A1(_25969_),
    .A2(_25974_),
    .A3(_25976_),
    .A4(_25981_),
    .ZN(_25982_));
 AND3_X1 _57220_ (.A1(_22920_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [338]),
    .A3(_23643_),
    .ZN(_25983_));
 AOI221_X4 _57221_ (.A(_25983_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [289]),
    .B2(_22777_),
    .C1(_23615_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [387]),
    .ZN(_25984_));
 NAND3_X1 _57222_ (.A1(_23982_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [142]),
    .A3(_23246_),
    .ZN(_25985_));
 AOI22_X2 _57223_ (.A1(_23164_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [44]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [93]),
    .B2(_11211_),
    .ZN(_25986_));
 NAND3_X1 _57224_ (.A1(_23367_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [240]),
    .A3(_23250_),
    .ZN(_25987_));
 NAND3_X1 _57225_ (.A1(_23003_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [191]),
    .A3(_23250_),
    .ZN(_25988_));
 AND4_X4 _57226_ (.A1(_25985_),
    .A2(_25986_),
    .A3(_25987_),
    .A4(_25988_),
    .ZN(_25989_));
 NAND3_X1 _57227_ (.A1(_23982_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [926]),
    .A3(_23321_),
    .ZN(_25990_));
 AOI22_X2 _57228_ (.A1(_23267_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [828]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [877]),
    .B2(_22544_),
    .ZN(_25991_));
 NAND3_X1 _57229_ (.A1(_23003_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [975]),
    .A3(_11081_),
    .ZN(_25992_));
 NAND3_X1 _57230_ (.A1(_23757_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1073]),
    .A3(_23879_),
    .ZN(_25993_));
 AND4_X4 _57231_ (.A1(_25990_),
    .A2(_25991_),
    .A3(_25992_),
    .A4(_25993_),
    .ZN(_25994_));
 NAND3_X1 _57232_ (.A1(_24262_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1171]),
    .A3(_23329_),
    .ZN(_25995_));
 NAND3_X1 _57233_ (.A1(_23328_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1024]),
    .A3(_23329_),
    .ZN(_25996_));
 NAND3_X1 _57234_ (.A1(_23240_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1122]),
    .A3(_23329_),
    .ZN(_25997_));
 AND3_X4 _57235_ (.A1(_25995_),
    .A2(_25996_),
    .A3(_25997_),
    .ZN(_25998_));
 AND4_X4 _57236_ (.A1(_25984_),
    .A2(_25989_),
    .A3(_25994_),
    .A4(_25998_),
    .ZN(_25999_));
 AOI22_X4 _57237_ (.A1(_23638_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [779]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [730]),
    .B2(_23092_),
    .ZN(_26000_));
 NAND3_X1 _57238_ (.A1(_22242_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [681]),
    .A3(_22995_),
    .ZN(_26001_));
 NAND3_X2 _57239_ (.A1(_23368_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [632]),
    .A3(_23057_),
    .ZN(_26002_));
 NAND3_X2 _57240_ (.A1(_23114_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [485]),
    .A3(_23057_),
    .ZN(_26003_));
 NAND4_X4 _57241_ (.A1(_26000_),
    .A2(_26001_),
    .A3(_26002_),
    .A4(_26003_),
    .ZN(_26004_));
 AOI22_X4 _57242_ (.A1(_23315_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1563]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1514]),
    .B2(_23095_),
    .ZN(_26005_));
 NAND3_X2 _57243_ (.A1(_23059_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1416]),
    .A3(_24026_),
    .ZN(_26006_));
 NAND3_X2 _57244_ (.A1(_22968_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1220]),
    .A3(_11037_),
    .ZN(_26007_));
 NAND3_X2 _57245_ (.A1(_24029_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1465]),
    .A3(_23566_),
    .ZN(_26008_));
 NAND4_X4 _57246_ (.A1(_26005_),
    .A2(_26006_),
    .A3(_26007_),
    .A4(_26008_),
    .ZN(_26009_));
 NAND3_X2 _57247_ (.A1(_23036_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1269]),
    .A3(_23274_),
    .ZN(_26010_));
 NAND3_X2 _57248_ (.A1(_23025_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1318]),
    .A3(_23277_),
    .ZN(_26011_));
 OAI211_X4 _57249_ (.A(_26010_),
    .B(_26011_),
    .C1(_11055_),
    .C2(_22310_),
    .ZN(_26012_));
 NAND3_X2 _57250_ (.A1(_23421_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [583]),
    .A3(_23072_),
    .ZN(_26013_));
 NAND3_X2 _57251_ (.A1(_23085_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [436]),
    .A3(_23208_),
    .ZN(_26014_));
 OAI211_X4 _57252_ (.A(_26013_),
    .B(_26014_),
    .C1(_11154_),
    .C2(_22721_),
    .ZN(_26015_));
 NOR4_X4 _57253_ (.A1(_26004_),
    .A2(_26009_),
    .A3(_26012_),
    .A4(_26015_),
    .ZN(_26016_));
 AND3_X1 _57254_ (.A1(_23751_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1906]),
    .A3(_23519_),
    .ZN(_26017_));
 AOI221_X4 _57255_ (.A(_26017_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1857]),
    .B2(_22044_),
    .C1(_23584_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1955]),
    .ZN(_26018_));
 NAND3_X1 _57256_ (.A1(_22241_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2641]),
    .A3(_10892_),
    .ZN(_26019_));
 AOI22_X1 _57257_ (.A1(_10929_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2396]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2445]),
    .B2(_23301_),
    .ZN(_26020_));
 NAND3_X1 _57258_ (.A1(_22523_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2494]),
    .A3(_23119_),
    .ZN(_26021_));
 NAND3_X1 _57259_ (.A1(_23003_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2543]),
    .A3(_23119_),
    .ZN(_26022_));
 AND4_X2 _57260_ (.A1(_26019_),
    .A2(_26020_),
    .A3(_26021_),
    .A4(_26022_),
    .ZN(_26023_));
 NAND3_X1 _57261_ (.A1(_23242_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1808]),
    .A3(_10989_),
    .ZN(_26024_));
 AOI22_X2 _57262_ (.A1(_23395_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1612]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1661]),
    .B2(_11019_),
    .ZN(_26025_));
 NAND3_X1 _57263_ (.A1(_23019_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1759]),
    .A3(_23398_),
    .ZN(_26026_));
 NAND3_X1 _57264_ (.A1(_23306_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1710]),
    .A3(_23398_),
    .ZN(_26027_));
 AND4_X4 _57265_ (.A1(_26024_),
    .A2(_26025_),
    .A3(_26026_),
    .A4(_26027_),
    .ZN(_26028_));
 AND3_X1 _57266_ (.A1(_23408_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2690]),
    .A3(_23310_),
    .ZN(_26029_));
 AOI221_X4 _57267_ (.A(_26029_),
    .B1(_21654_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2592]),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2739]),
    .C2(_21573_),
    .ZN(_26030_));
 AND4_X4 _57268_ (.A1(_26018_),
    .A2(_26023_),
    .A3(_26028_),
    .A4(_26030_),
    .ZN(_26031_));
 NAND4_X4 _57269_ (.A1(_25982_),
    .A2(_25999_),
    .A3(net1),
    .A4(_26031_),
    .ZN(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [44]));
 NAND3_X1 _57270_ (.A1(_23221_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [633]),
    .A3(_23237_),
    .ZN(_26032_));
 NAND3_X1 _57271_ (.A1(_10780_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [976]),
    .A3(_23317_),
    .ZN(_26033_));
 NAND3_X1 _57272_ (.A1(_23385_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [682]),
    .A3(_23237_),
    .ZN(_26034_));
 NAND3_X4 _57273_ (.A1(_23982_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1319]),
    .A3(_23412_),
    .ZN(_26035_));
 AND4_X4 _57274_ (.A1(_26032_),
    .A2(_26033_),
    .A3(_26034_),
    .A4(_26035_),
    .ZN(_26036_));
 NAND3_X2 _57275_ (.A1(_23150_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1564]),
    .A3(_11035_),
    .ZN(_26037_));
 NAND3_X4 _57276_ (.A1(_22915_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [878]),
    .A3(_22905_),
    .ZN(_26038_));
 NAND2_X4 _57277_ (.A1(_26037_),
    .A2(_26038_),
    .ZN(_26039_));
 AOI221_X4 _57278_ (.A(_26039_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1809]),
    .B2(_11002_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1613]),
    .C2(_23395_),
    .ZN(_26040_));
 NAND3_X4 _57279_ (.A1(_22920_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [731]),
    .A3(_23151_),
    .ZN(_26041_));
 NAND3_X2 _57280_ (.A1(_23775_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [486]),
    .A3(_23510_),
    .ZN(_26042_));
 NAND2_X4 _57281_ (.A1(_26041_),
    .A2(_26042_),
    .ZN(_26043_));
 AOI221_X4 _57282_ (.A(_26043_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [535]),
    .B2(_11152_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2348]),
    .C2(_23097_),
    .ZN(_26044_));
 NAND3_X1 _57283_ (.A1(_22942_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2299]),
    .A3(_22913_),
    .ZN(_26045_));
 NAND3_X4 _57284_ (.A1(_23806_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1270]),
    .A3(_23848_),
    .ZN(_26046_));
 NAND2_X1 _57285_ (.A1(_26045_),
    .A2(_26046_),
    .ZN(_26047_));
 AOI221_X4 _57286_ (.A(_26047_),
    .B1(_10955_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2201]),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2152]),
    .C2(_10962_),
    .ZN(_26048_));
 AND4_X1 _57287_ (.A1(_26036_),
    .A2(_26040_),
    .A3(_26044_),
    .A4(_26048_),
    .ZN(_26049_));
 NAND3_X1 _57288_ (.A1(_23150_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2740]),
    .A3(_23481_),
    .ZN(_26050_));
 NAND3_X1 _57289_ (.A1(_23150_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3132]),
    .A3(_10788_),
    .ZN(_26051_));
 NAND2_X1 _57290_ (.A1(_26050_),
    .A2(_26051_),
    .ZN(_26052_));
 AOI221_X2 _57291_ (.A(_26052_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2691]),
    .B2(_23374_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [437]),
    .C2(_23610_),
    .ZN(_26053_));
 NAND3_X4 _57292_ (.A1(_23509_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [192]),
    .A3(_23643_),
    .ZN(_26054_));
 NAND3_X1 _57293_ (.A1(_23806_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2054]),
    .A3(_23231_),
    .ZN(_26055_));
 NAND2_X2 _57294_ (.A1(_26054_),
    .A2(_26055_),
    .ZN(_26056_));
 AOI221_X4 _57295_ (.A(_26056_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2103]),
    .B2(_23233_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1760]),
    .C2(_22078_),
    .ZN(_26057_));
 NAND3_X4 _57296_ (.A1(_24467_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1858]),
    .A3(_22923_),
    .ZN(_26058_));
 NAND3_X1 _57297_ (.A1(_24467_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3034]),
    .A3(_23174_),
    .ZN(_26059_));
 NAND2_X1 _57298_ (.A1(_26058_),
    .A2(_26059_),
    .ZN(_26060_));
 AOI221_X2 _57299_ (.A(_26060_),
    .B1(_23225_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3083]),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2789]),
    .C2(_21289_),
    .ZN(_26061_));
 NAND3_X1 _57300_ (.A1(_10856_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2887]),
    .A3(_23794_),
    .ZN(_26062_));
 NAND3_X1 _57301_ (.A1(_23176_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2838]),
    .A3(_23174_),
    .ZN(_26063_));
 NAND2_X1 _57302_ (.A1(_26062_),
    .A2(_26063_),
    .ZN(_26064_));
 AOI221_X4 _57303_ (.A(_26064_),
    .B1(_22918_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2985]),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2936]),
    .C2(_21466_),
    .ZN(_26065_));
 AND4_X4 _57304_ (.A1(_26053_),
    .A2(_26057_),
    .A3(_26061_),
    .A4(_26065_),
    .ZN(_26066_));
 AND3_X1 _57305_ (.A1(_10817_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1907]),
    .A3(_22934_),
    .ZN(_26067_));
 AOI21_X4 _57306_ (.A(_26067_),
    .B1(_23584_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1956]),
    .ZN(_26068_));
 OAI221_X2 _57307_ (.A(_26068_),
    .B1(_22230_),
    .B2(_11042_),
    .C1(_22312_),
    .C2(_11055_),
    .ZN(_26069_));
 NAND3_X1 _57308_ (.A1(_23008_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2397]),
    .A3(_23131_),
    .ZN(_26070_));
 NAND3_X1 _57309_ (.A1(_23377_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2446]),
    .A3(_23131_),
    .ZN(_26071_));
 NAND3_X1 _57310_ (.A1(_23016_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2495]),
    .A3(_23014_),
    .ZN(_26072_));
 NAND3_X4 _57311_ (.A1(_24029_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1466]),
    .A3(_23566_),
    .ZN(_26073_));
 NAND4_X2 _57312_ (.A1(_26070_),
    .A2(_26071_),
    .A3(_26072_),
    .A4(_26073_),
    .ZN(_26074_));
 NAND3_X4 _57313_ (.A1(_23067_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1172]),
    .A3(_23882_),
    .ZN(_26075_));
 NAND3_X1 _57314_ (.A1(_23200_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2544]),
    .A3(_23023_),
    .ZN(_26076_));
 NAND3_X1 _57315_ (.A1(_23276_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2593]),
    .A3(_23143_),
    .ZN(_26077_));
 NAND3_X4 _57316_ (.A1(_23271_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1025]),
    .A3(_23891_),
    .ZN(_26078_));
 NAND4_X1 _57317_ (.A1(_26075_),
    .A2(_26076_),
    .A3(_26077_),
    .A4(_26078_),
    .ZN(_26079_));
 NAND3_X2 _57318_ (.A1(_10844_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1417]),
    .A3(_23274_),
    .ZN(_26080_));
 NAND3_X4 _57319_ (.A1(_23837_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [829]),
    .A3(_22976_),
    .ZN(_26081_));
 NAND3_X1 _57320_ (.A1(_23280_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1123]),
    .A3(_23547_),
    .ZN(_26082_));
 NAND3_X2 _57321_ (.A1(_23575_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1074]),
    .A3(_23317_),
    .ZN(_26083_));
 NAND4_X4 _57322_ (.A1(_26080_),
    .A2(_26081_),
    .A3(_26082_),
    .A4(_26083_),
    .ZN(_26084_));
 NOR4_X1 _57323_ (.A1(_26069_),
    .A2(_26074_),
    .A3(_26079_),
    .A4(_26084_),
    .ZN(_26085_));
 NAND3_X4 _57324_ (.A1(_24126_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [780]),
    .A3(_22995_),
    .ZN(_26086_));
 NAND3_X4 _57325_ (.A1(_23114_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1662]),
    .A3(_23116_),
    .ZN(_26087_));
 NAND3_X2 _57326_ (.A1(_10858_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1711]),
    .A3(_23116_),
    .ZN(_26088_));
 NAND3_X4 _57327_ (.A1(_22933_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [241]),
    .A3(_23341_),
    .ZN(_26089_));
 NAND4_X1 _57328_ (.A1(_26086_),
    .A2(_26087_),
    .A3(_26088_),
    .A4(_26089_),
    .ZN(_26090_));
 NAND3_X2 _57329_ (.A1(_22950_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [388]),
    .A3(_22940_),
    .ZN(_26091_));
 NAND3_X2 _57330_ (.A1(_23536_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [290]),
    .A3(_11176_),
    .ZN(_26092_));
 NAND3_X2 _57331_ (.A1(_24050_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [339]),
    .A3(_23187_),
    .ZN(_26093_));
 NAND3_X2 _57332_ (.A1(_23189_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [94]),
    .A3(_23835_),
    .ZN(_26094_));
 NAND4_X4 _57333_ (.A1(_26091_),
    .A2(_26092_),
    .A3(_26093_),
    .A4(_26094_),
    .ZN(_26095_));
 NAND3_X2 _57334_ (.A1(_22955_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [584]),
    .A3(_23063_),
    .ZN(_26096_));
 NAND3_X1 _57335_ (.A1(_23025_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [143]),
    .A3(_22959_),
    .ZN(_26097_));
 NAND3_X1 _57336_ (.A1(_23837_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [45]),
    .A3(_23196_),
    .ZN(_26098_));
 NAND3_X4 _57337_ (.A1(_23080_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2642]),
    .A3(_23043_),
    .ZN(_26099_));
 NAND4_X1 _57338_ (.A1(_26096_),
    .A2(_26097_),
    .A3(_26098_),
    .A4(_26099_),
    .ZN(_26100_));
 NAND3_X1 _57339_ (.A1(_23022_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1221]),
    .A3(_23274_),
    .ZN(_26101_));
 NAND3_X4 _57340_ (.A1(_23837_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2005]),
    .A3(_23832_),
    .ZN(_26102_));
 NAND3_X4 _57341_ (.A1(_23204_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [927]),
    .A3(_23317_),
    .ZN(_26103_));
 NAND3_X4 _57342_ (.A1(_23438_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2250]),
    .A3(_23600_),
    .ZN(_26104_));
 NAND4_X2 _57343_ (.A1(_26101_),
    .A2(_26102_),
    .A3(_26103_),
    .A4(_26104_),
    .ZN(_26105_));
 NOR4_X1 _57344_ (.A1(_26090_),
    .A2(_26095_),
    .A3(_26100_),
    .A4(_26105_),
    .ZN(_26106_));
 NAND4_X1 _57345_ (.A1(_26049_),
    .A2(_26066_),
    .A3(_26085_),
    .A4(_26106_),
    .ZN(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [45]));
 NAND3_X1 _57346_ (.A1(_23288_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [928]),
    .A3(_22905_),
    .ZN(_26107_));
 NAND3_X4 _57347_ (.A1(_10829_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1859]),
    .A3(_22921_),
    .ZN(_26108_));
 NAND2_X1 _57348_ (.A1(_26107_),
    .A2(_26108_),
    .ZN(_26109_));
 AOI221_X4 _57349_ (.A(_26109_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [536]),
    .B2(_23689_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1026]),
    .C2(_23104_),
    .ZN(_26110_));
 NAND3_X1 _57350_ (.A1(_23150_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [781]),
    .A3(_23504_),
    .ZN(_26111_));
 NAND3_X1 _57351_ (.A1(_22900_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [634]),
    .A3(_23504_),
    .ZN(_26112_));
 NAND2_X2 _57352_ (.A1(_26111_),
    .A2(_26112_),
    .ZN(_26113_));
 AOI221_X2 _57353_ (.A(_26113_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1124]),
    .B2(_22410_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1075]),
    .C2(_23632_),
    .ZN(_26114_));
 NAND3_X2 _57354_ (.A1(_23492_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1173]),
    .A3(_22905_),
    .ZN(_26115_));
 NAND3_X2 _57355_ (.A1(_23775_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [487]),
    .A3(_23510_),
    .ZN(_26116_));
 NAND2_X4 _57356_ (.A1(_26115_),
    .A2(_26116_),
    .ZN(_26117_));
 AOI221_X2 _57357_ (.A(_26117_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2986]),
    .B2(_22918_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2202]),
    .C2(_23660_),
    .ZN(_26118_));
 NAND3_X1 _57358_ (.A1(_23153_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1418]),
    .A3(_11035_),
    .ZN(_26119_));
 NAND3_X1 _57359_ (.A1(_10856_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1320]),
    .A3(_23848_),
    .ZN(_26120_));
 NAND2_X2 _57360_ (.A1(_26119_),
    .A2(_26120_),
    .ZN(_26121_));
 AOI221_X4 _57361_ (.A(_26121_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2104]),
    .B2(_23233_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1565]),
    .C2(_23179_),
    .ZN(_26122_));
 AND4_X1 _57362_ (.A1(_26110_),
    .A2(_26114_),
    .A3(_26118_),
    .A4(_26122_),
    .ZN(_26123_));
 AND3_X1 _57363_ (.A1(_23084_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [830]),
    .A3(_22969_),
    .ZN(_26124_));
 AOI21_X4 _57364_ (.A(_26124_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [879]),
    .B2(_23268_),
    .ZN(_26125_));
 OAI221_X2 _57365_ (.A(_26125_),
    .B1(_22861_),
    .B2(_11201_),
    .C1(_22879_),
    .C2(_11207_),
    .ZN(_26126_));
 NAND3_X2 _57366_ (.A1(_24126_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1957]),
    .A3(_22935_),
    .ZN(_26127_));
 NAND3_X1 _57367_ (.A1(_23125_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1761]),
    .A3(_22935_),
    .ZN(_26128_));
 NAND3_X1 _57368_ (.A1(_23059_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1810]),
    .A3(_23009_),
    .ZN(_26129_));
 NAND3_X2 _57369_ (.A1(_23127_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1908]),
    .A3(_23009_),
    .ZN(_26130_));
 NAND4_X4 _57370_ (.A1(_26127_),
    .A2(_26128_),
    .A3(_26129_),
    .A4(_26130_),
    .ZN(_26131_));
 NAND3_X4 _57371_ (.A1(_24045_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [193]),
    .A3(_22951_),
    .ZN(_26132_));
 NAND3_X2 _57372_ (.A1(_23076_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2741]),
    .A3(_23134_),
    .ZN(_26133_));
 NAND3_X4 _57373_ (.A1(_23189_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1663]),
    .A3(_23141_),
    .ZN(_26134_));
 NAND3_X4 _57374_ (.A1(_23025_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1712]),
    .A3(_23830_),
    .ZN(_26135_));
 NAND4_X2 _57375_ (.A1(_26132_),
    .A2(_26133_),
    .A3(_26134_),
    .A4(_26135_),
    .ZN(_26136_));
 NAND3_X4 _57376_ (.A1(_23020_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [585]),
    .A3(_23063_),
    .ZN(_26137_));
 NAND3_X1 _57377_ (.A1(_22972_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2692]),
    .A3(_23023_),
    .ZN(_26138_));
 NAND3_X1 _57378_ (.A1(_23276_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2594]),
    .A3(_23143_),
    .ZN(_26139_));
 NAND3_X2 _57379_ (.A1(_22978_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2643]),
    .A3(_23029_),
    .ZN(_26140_));
 NAND4_X2 _57380_ (.A1(_26137_),
    .A2(_26138_),
    .A3(_26139_),
    .A4(_26140_),
    .ZN(_26141_));
 NOR4_X2 _57381_ (.A1(_26126_),
    .A2(_26131_),
    .A3(_26136_),
    .A4(_26141_),
    .ZN(_26142_));
 AND3_X1 _57382_ (.A1(_10857_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2888]),
    .A3(_10789_),
    .ZN(_26143_));
 AOI21_X1 _57383_ (.A(_26143_),
    .B1(_23213_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2937]),
    .ZN(_26144_));
 OAI221_X2 _57384_ (.A(_26144_),
    .B1(_21570_),
    .B2(_10864_),
    .C1(_21960_),
    .C2(_10973_),
    .ZN(_26145_));
 NAND3_X4 _57385_ (.A1(_23054_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [389]),
    .A3(_22940_),
    .ZN(_26146_));
 NAND3_X2 _57386_ (.A1(_24045_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1369]),
    .A3(_24026_),
    .ZN(_26147_));
 NAND3_X2 _57387_ (.A1(_24045_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2545]),
    .A3(_23014_),
    .ZN(_26148_));
 NAND3_X2 _57388_ (.A1(_23133_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1614]),
    .A3(_22956_),
    .ZN(_26149_));
 NAND4_X4 _57389_ (.A1(_26146_),
    .A2(_26147_),
    .A3(_26148_),
    .A4(_26149_),
    .ZN(_26150_));
 NAND3_X2 _57390_ (.A1(_23011_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [242]),
    .A3(_23187_),
    .ZN(_26151_));
 NAND3_X2 _57391_ (.A1(_23022_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1222]),
    .A3(_23274_),
    .ZN(_26152_));
 NAND3_X2 _57392_ (.A1(_23194_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2398]),
    .A3(_23143_),
    .ZN(_26153_));
 NAND3_X2 _57393_ (.A1(_23071_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [291]),
    .A3(_23196_),
    .ZN(_26154_));
 NAND4_X4 _57394_ (.A1(_26151_),
    .A2(_26152_),
    .A3(_26153_),
    .A4(_26154_),
    .ZN(_26155_));
 NAND3_X2 _57395_ (.A1(_23200_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [977]),
    .A3(_22973_),
    .ZN(_26156_));
 NAND3_X2 _57396_ (.A1(_22975_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [683]),
    .A3(_23072_),
    .ZN(_26157_));
 NAND3_X2 _57397_ (.A1(_23280_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [732]),
    .A3(_23208_),
    .ZN(_26158_));
 NAND3_X2 _57398_ (.A1(_23085_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [438]),
    .A3(_23208_),
    .ZN(_26159_));
 NAND4_X4 _57399_ (.A1(_26156_),
    .A2(_26157_),
    .A3(_26158_),
    .A4(_26159_),
    .ZN(_26160_));
 NOR4_X1 _57400_ (.A1(_26145_),
    .A2(_26150_),
    .A3(_26155_),
    .A4(_26160_),
    .ZN(_26161_));
 NAND3_X4 _57401_ (.A1(_22988_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2153]),
    .A3(_23554_),
    .ZN(_26162_));
 NAND3_X4 _57402_ (.A1(_24126_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3133]),
    .A3(_22991_),
    .ZN(_26163_));
 NAND3_X4 _57403_ (.A1(_22994_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2006]),
    .A3(_23554_),
    .ZN(_26164_));
 NAND3_X4 _57404_ (.A1(_10831_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3035]),
    .A3(_23123_),
    .ZN(_26165_));
 NAND4_X4 _57405_ (.A1(_26162_),
    .A2(_26163_),
    .A3(_26164_),
    .A4(_26165_),
    .ZN(_26166_));
 NAND3_X1 _57406_ (.A1(_22950_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2349]),
    .A3(_23006_),
    .ZN(_26167_));
 NAND3_X4 _57407_ (.A1(_23127_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [340]),
    .A3(_11176_),
    .ZN(_26168_));
 NAND3_X2 _57408_ (.A1(_24029_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2251]),
    .A3(_24046_),
    .ZN(_26169_));
 NAND3_X2 _57409_ (.A1(_23888_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2300]),
    .A3(_24052_),
    .ZN(_26170_));
 NAND4_X4 _57410_ (.A1(_26167_),
    .A2(_26168_),
    .A3(_26169_),
    .A4(_26170_),
    .ZN(_26171_));
 NAND3_X4 _57411_ (.A1(_23133_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2790]),
    .A3(_23033_),
    .ZN(_26172_));
 NAND3_X4 _57412_ (.A1(_22972_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3084]),
    .A3(_10790_),
    .ZN(_26173_));
 NAND3_X4 _57413_ (.A1(_23028_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1516]),
    .A3(_22981_),
    .ZN(_26174_));
 NAND3_X4 _57414_ (.A1(_23080_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1467]),
    .A3(_23205_),
    .ZN(_26175_));
 NAND4_X2 _57415_ (.A1(_26172_),
    .A2(_26173_),
    .A3(_26174_),
    .A4(_26175_),
    .ZN(_26176_));
 NAND3_X1 _57416_ (.A1(_23140_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2496]),
    .A3(_23023_),
    .ZN(_26177_));
 NAND3_X2 _57417_ (.A1(_23145_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [95]),
    .A3(_23196_),
    .ZN(_26178_));
 NAND3_X4 _57418_ (.A1(_23042_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1271]),
    .A3(_23205_),
    .ZN(_26179_));
 NAND3_X1 _57419_ (.A1(_23426_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2447]),
    .A3(_23422_),
    .ZN(_26180_));
 NAND4_X2 _57420_ (.A1(_26177_),
    .A2(_26178_),
    .A3(_26179_),
    .A4(_26180_),
    .ZN(_26181_));
 NOR4_X4 _57421_ (.A1(_26166_),
    .A2(_26171_),
    .A3(_26176_),
    .A4(_26181_),
    .ZN(_26182_));
 NAND4_X1 _57422_ (.A1(_26123_),
    .A2(_26142_),
    .A3(_26161_),
    .A4(_26182_),
    .ZN(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [46]));
 NAND3_X1 _57423_ (.A1(_23280_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1517]),
    .A3(_23931_),
    .ZN(_26183_));
 AOI22_X1 _57424_ (.A1(_23325_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1223]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1468]),
    .B2(_23326_),
    .ZN(_26184_));
 NAND3_X1 _57425_ (.A1(_24262_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1566]),
    .A3(_23412_),
    .ZN(_26185_));
 NAND3_X1 _57426_ (.A1(_23328_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1419]),
    .A3(_23412_),
    .ZN(_26186_));
 AND4_X2 _57427_ (.A1(_26183_),
    .A2(_26184_),
    .A3(_26185_),
    .A4(_26186_),
    .ZN(_26187_));
 NAND3_X1 _57428_ (.A1(_10868_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1272]),
    .A3(_23931_),
    .ZN(_26188_));
 AND3_X1 _57429_ (.A1(_10873_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [831]),
    .A3(_11089_),
    .ZN(_26189_));
 AOI221_X2 _57430_ (.A(_26189_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [929]),
    .B2(_11105_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [978]),
    .C2(_11099_),
    .ZN(_26190_));
 NAND3_X1 _57431_ (.A1(_10780_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1370]),
    .A3(_23693_),
    .ZN(_26191_));
 NAND3_X1 _57432_ (.A1(_22523_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1321]),
    .A3(_23693_),
    .ZN(_26192_));
 AND4_X2 _57433_ (.A1(_26188_),
    .A2(net57),
    .A3(_26191_),
    .A4(_26192_),
    .ZN(_26193_));
 AND3_X1 _57434_ (.A1(_23284_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1174]),
    .A3(_23494_),
    .ZN(_26194_));
 AOI221_X2 _57435_ (.A(_26194_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1125]),
    .B2(_22410_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1076]),
    .C2(_23632_),
    .ZN(_26195_));
 AOI22_X2 _57436_ (.A1(_22459_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1027]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [880]),
    .B2(_23268_),
    .ZN(_26196_));
 AND4_X4 _57437_ (.A1(_26187_),
    .A2(_26193_),
    .A3(_26195_),
    .A4(_26196_),
    .ZN(_26197_));
 NAND3_X1 _57438_ (.A1(_23421_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2938]),
    .A3(_23431_),
    .ZN(_26198_));
 AND3_X1 _57439_ (.A1(_10855_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2497]),
    .A3(_10890_),
    .ZN(_26199_));
 AOI221_X2 _57440_ (.A(_26199_),
    .B1(_10928_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2399]),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2546]),
    .C2(_10912_),
    .ZN(_26200_));
 NAND3_X1 _57441_ (.A1(_10868_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2840]),
    .A3(_23673_),
    .ZN(_26201_));
 NAND3_X2 _57442_ (.A1(_23982_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2889]),
    .A3(_23222_),
    .ZN(_26202_));
 AND4_X1 _57443_ (.A1(_26198_),
    .A2(_26200_),
    .A3(_26201_),
    .A4(_26202_),
    .ZN(_26203_));
 NAND3_X1 _57444_ (.A1(_23438_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3036]),
    .A3(_23431_),
    .ZN(_26204_));
 AOI22_X1 _57445_ (.A1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2791]),
    .A2(_23625_),
    .B1(_10839_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2987]),
    .ZN(_26205_));
 NAND3_X1 _57446_ (.A1(_24262_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3134]),
    .A3(_23222_),
    .ZN(_26206_));
 NAND3_X1 _57447_ (.A1(_24186_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3085]),
    .A3(_23222_),
    .ZN(_26207_));
 AND4_X2 _57448_ (.A1(_26204_),
    .A2(_26205_),
    .A3(_26206_),
    .A4(_26207_),
    .ZN(_26208_));
 NAND3_X1 _57449_ (.A1(_23438_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2644]),
    .A3(_23427_),
    .ZN(_26209_));
 AOI22_X4 _57450_ (.A1(_21654_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2595]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2448]),
    .B2(_10922_),
    .ZN(_26210_));
 NAND3_X1 _57451_ (.A1(_23245_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2742]),
    .A3(_23427_),
    .ZN(_26211_));
 NAND3_X1 _57452_ (.A1(_23240_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2693]),
    .A3(_23427_),
    .ZN(_26212_));
 AND4_X1 _57453_ (.A1(_26209_),
    .A2(_26210_),
    .A3(_26211_),
    .A4(_26212_),
    .ZN(_26213_));
 AND3_X4 _57454_ (.A1(_26203_),
    .A2(_26208_),
    .A3(_26213_),
    .ZN(_26214_));
 NAND3_X1 _57455_ (.A1(_24262_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [390]),
    .A3(_23709_),
    .ZN(_26215_));
 AOI22_X1 _57456_ (.A1(_23248_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [243]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [96]),
    .B2(_23714_),
    .ZN(_26216_));
 NAND3_X1 _57457_ (.A1(_22241_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [292]),
    .A3(_23451_),
    .ZN(_26217_));
 NAND3_X1 _57458_ (.A1(_23935_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [341]),
    .A3(_23451_),
    .ZN(_26218_));
 AND4_X1 _57459_ (.A1(_26215_),
    .A2(_26216_),
    .A3(_26217_),
    .A4(_26218_),
    .ZN(_26219_));
 NAND3_X2 _57460_ (.A1(_23158_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [586]),
    .A3(_23512_),
    .ZN(_26220_));
 NAND3_X2 _57461_ (.A1(_23173_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [537]),
    .A3(_23161_),
    .ZN(_26221_));
 NAND2_X4 _57462_ (.A1(_26220_),
    .A2(_26221_),
    .ZN(_26222_));
 AOI221_X4 _57463_ (.A(_26222_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [488]),
    .B2(_11158_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [439]),
    .C2(_22733_),
    .ZN(_26223_));
 NAND3_X1 _57464_ (.A1(_23242_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [635]),
    .A3(_23346_),
    .ZN(_26224_));
 NAND3_X1 _57465_ (.A1(_23390_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [782]),
    .A3(_23346_),
    .ZN(_26225_));
 NAND3_X1 _57466_ (.A1(_23757_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [684]),
    .A3(_23056_),
    .ZN(_26226_));
 NAND3_X1 _57467_ (.A1(_22943_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [733]),
    .A3(_23056_),
    .ZN(_26227_));
 AND4_X4 _57468_ (.A1(_26224_),
    .A2(_26225_),
    .A3(_26226_),
    .A4(_26227_),
    .ZN(_26228_));
 AND3_X1 _57469_ (.A1(_22521_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [145]),
    .A3(_22937_),
    .ZN(_26229_));
 AOI221_X4 _57470_ (.A(_26229_),
    .B1(_11205_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [47]),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [194]),
    .C2(_22806_),
    .ZN(_26230_));
 AND4_X4 _57471_ (.A1(_26219_),
    .A2(_26223_),
    .A3(_26228_),
    .A4(_26230_),
    .ZN(_26231_));
 NAND3_X1 _57472_ (.A1(_22954_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2154]),
    .A3(_22963_),
    .ZN(_26232_));
 OAI21_X2 _57473_ (.A(_26232_),
    .B1(_10969_),
    .B2(_21936_),
    .ZN(_26233_));
 NAND3_X4 _57474_ (.A1(_10878_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2007]),
    .A3(_10940_),
    .ZN(_26234_));
 OAI21_X1 _57475_ (.A(_26234_),
    .B1(_10973_),
    .B2(_21963_),
    .ZN(_26235_));
 NAND3_X1 _57476_ (.A1(_10779_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1762]),
    .A3(_22934_),
    .ZN(_26236_));
 NAND3_X2 _57477_ (.A1(_22522_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1713]),
    .A3(_22934_),
    .ZN(_26237_));
 NAND2_X4 _57478_ (.A1(_26236_),
    .A2(_26237_),
    .ZN(_26238_));
 AND3_X2 _57479_ (.A1(_10878_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1615]),
    .A3(_10988_),
    .ZN(_26239_));
 OR4_X2 _57480_ (.A1(_26233_),
    .A2(_26235_),
    .A3(_26238_),
    .A4(_26239_),
    .ZN(_26240_));
 NAND3_X4 _57481_ (.A1(_22933_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1811]),
    .A3(_22935_),
    .ZN(_26241_));
 OAI21_X4 _57482_ (.A(_26241_),
    .B1(_11020_),
    .B2(_22159_),
    .ZN(_26242_));
 NAND3_X1 _57483_ (.A1(_22958_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1860]),
    .A3(_23830_),
    .ZN(_26243_));
 NAND3_X1 _57484_ (.A1(_22961_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1909]),
    .A3(_23830_),
    .ZN(_26244_));
 OAI211_X2 _57485_ (.A(_26243_),
    .B(_26244_),
    .C1(_10984_),
    .C2(_22002_),
    .ZN(_26245_));
 NAND3_X1 _57486_ (.A1(_23236_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2350]),
    .A3(_22964_),
    .ZN(_26246_));
 NAND3_X2 _57487_ (.A1(_23028_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2301]),
    .A3(_23832_),
    .ZN(_26247_));
 NAND3_X2 _57488_ (.A1(_23839_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2203]),
    .A3(_23081_),
    .ZN(_26248_));
 NAND3_X2 _57489_ (.A1(_23438_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2252]),
    .A3(_23600_),
    .ZN(_26249_));
 NAND4_X4 _57490_ (.A1(_26246_),
    .A2(_26247_),
    .A3(_26248_),
    .A4(_26249_),
    .ZN(_26250_));
 NOR4_X4 _57491_ (.A1(_26240_),
    .A2(_26242_),
    .A3(_26245_),
    .A4(_26250_),
    .ZN(_26251_));
 NAND4_X2 _57492_ (.A1(_26197_),
    .A2(_26214_),
    .A3(_26231_),
    .A4(net6),
    .ZN(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [47]));
 AND3_X1 _57493_ (.A1(_23459_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1175]),
    .A3(_23804_),
    .ZN(_26252_));
 AOI221_X2 _57494_ (.A(_26252_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1126]),
    .B2(_22410_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1077]),
    .C2(_23632_),
    .ZN(_26253_));
 AOI22_X4 _57495_ (.A1(_22459_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1028]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [881]),
    .B2(_23268_),
    .ZN(_26254_));
 AND3_X1 _57496_ (.A1(_10816_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [342]),
    .A3(_22937_),
    .ZN(_26255_));
 AOI221_X2 _57497_ (.A(_26255_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [293]),
    .B2(_22777_),
    .C1(_11170_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [391]),
    .ZN(_26256_));
 AOI22_X4 _57498_ (.A1(_23248_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [244]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [97]),
    .B2(_23490_),
    .ZN(_26257_));
 NAND4_X2 _57499_ (.A1(net42),
    .A2(_26254_),
    .A3(_26256_),
    .A4(_26257_),
    .ZN(_26258_));
 AND3_X1 _57500_ (.A1(_10842_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1420]),
    .A3(_22979_),
    .ZN(_26259_));
 AOI221_X2 _57501_ (.A(_26259_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1518]),
    .B2(_11041_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1567]),
    .C2(_23179_),
    .ZN(_26260_));
 AND3_X1 _57502_ (.A1(_10877_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [832]),
    .A3(_11079_),
    .ZN(_26261_));
 AOI221_X2 _57503_ (.A(_26261_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [930]),
    .B2(_11106_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [979]),
    .C2(_11100_),
    .ZN(_26262_));
 NAND3_X2 _57504_ (.A1(_10831_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1469]),
    .A3(_22945_),
    .ZN(_26263_));
 NAND3_X1 _57505_ (.A1(_22954_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1371]),
    .A3(_22980_),
    .ZN(_26264_));
 NAND3_X1 _57506_ (.A1(_22522_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1322]),
    .A3(_22980_),
    .ZN(_26265_));
 NAND3_X1 _57507_ (.A1(_23041_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1273]),
    .A3(_22980_),
    .ZN(_26266_));
 NAND3_X1 _57508_ (.A1(_23084_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1224]),
    .A3(_22980_),
    .ZN(_26267_));
 AND4_X4 _57509_ (.A1(_26264_),
    .A2(_26265_),
    .A3(_26266_),
    .A4(_26267_),
    .ZN(_26268_));
 NAND4_X4 _57510_ (.A1(_26260_),
    .A2(net41),
    .A3(_26263_),
    .A4(_26268_),
    .ZN(_26269_));
 AND3_X1 _57511_ (.A1(_10877_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [48]),
    .A3(_22937_),
    .ZN(_26270_));
 AOI221_X2 _57512_ (.A(_26270_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [146]),
    .B2(_11200_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [195]),
    .C2(_11195_),
    .ZN(_26271_));
 NAND3_X2 _57513_ (.A1(_23008_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [440]),
    .A3(_23060_),
    .ZN(_26272_));
 NAND3_X2 _57514_ (.A1(_23062_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [489]),
    .A3(_23060_),
    .ZN(_26273_));
 AOI22_X4 _57515_ (.A1(_23622_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [587]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [538]),
    .B2(_11153_),
    .ZN(_26274_));
 NAND4_X4 _57516_ (.A1(_26271_),
    .A2(_26272_),
    .A3(_26273_),
    .A4(_26274_),
    .ZN(_26275_));
 AOI22_X4 _57517_ (.A1(_23638_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [783]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [734]),
    .B2(_23092_),
    .ZN(_26276_));
 NAND3_X2 _57518_ (.A1(_23192_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [636]),
    .A3(_23063_),
    .ZN(_26277_));
 OAI211_X4 _57519_ (.A(_26276_),
    .B(_26277_),
    .C1(_22663_),
    .C2(_11137_),
    .ZN(_26278_));
 NOR4_X4 _57520_ (.A1(_26258_),
    .A2(_26269_),
    .A3(_26275_),
    .A4(_26278_),
    .ZN(_26279_));
 OAI22_X1 _57521_ (.A1(_10875_),
    .A2(_21379_),
    .B1(_21572_),
    .B2(_10864_),
    .ZN(_26280_));
 AOI221_X4 _57522_ (.A(_26280_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2939]),
    .B2(_21466_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2890]),
    .C2(_21502_),
    .ZN(_26281_));
 NAND3_X1 _57523_ (.A1(_10845_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2988]),
    .A3(_23361_),
    .ZN(_26282_));
 AND3_X1 _57524_ (.A1(_22920_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3086]),
    .A3(_10788_),
    .ZN(_26283_));
 AOI221_X2 _57525_ (.A(_26283_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3037]),
    .B2(_10826_),
    .C1(_23224_),
    .C2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3135]),
    .ZN(_26284_));
 AND3_X1 _57526_ (.A1(_26281_),
    .A2(_26282_),
    .A3(_26284_),
    .ZN(_26285_));
 NAND3_X1 _57527_ (.A1(_23340_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2596]),
    .A3(_10893_),
    .ZN(_26286_));
 AND3_X1 _57528_ (.A1(_23810_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2743]),
    .A3(_23669_),
    .ZN(_26287_));
 AOI221_X2 _57529_ (.A(_26287_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2694]),
    .B2(_21601_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2645]),
    .C2(_23627_),
    .ZN(_26288_));
 AOI22_X2 _57530_ (.A1(_23587_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2547]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2498]),
    .B2(_21705_),
    .ZN(_26289_));
 AOI22_X2 _57531_ (.A1(_10929_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2400]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2449]),
    .B2(_10922_),
    .ZN(_26290_));
 AND4_X4 _57532_ (.A1(_26286_),
    .A2(_26288_),
    .A3(_26289_),
    .A4(_26290_),
    .ZN(_26291_));
 NAND3_X1 _57533_ (.A1(_10798_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2351]),
    .A3(_10939_),
    .ZN(_26292_));
 NAND3_X1 _57534_ (.A1(_23215_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2253]),
    .A3(_10939_),
    .ZN(_26293_));
 OAI211_X2 _57535_ (.A(_26292_),
    .B(_26293_),
    .C1(_10946_),
    .C2(_21845_),
    .ZN(_26294_));
 AOI221_X2 _57536_ (.A(_26294_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2204]),
    .B2(_10955_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2057]),
    .C2(_23156_),
    .ZN(_26295_));
 NAND3_X1 _57537_ (.A1(_23240_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1910]),
    .A3(_23393_),
    .ZN(_26296_));
 AOI22_X2 _57538_ (.A1(_11003_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1812]),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1665]),
    .B2(_23396_),
    .ZN(_26297_));
 NAND3_X1 _57539_ (.A1(_23390_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1959]),
    .A3(_23294_),
    .ZN(_26298_));
 NAND3_X1 _57540_ (.A1(_23757_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1861]),
    .A3(_23398_),
    .ZN(_26299_));
 AND4_X4 _57541_ (.A1(_26296_),
    .A2(_26297_),
    .A3(_26298_),
    .A4(_26299_),
    .ZN(_26300_));
 AND3_X1 _57542_ (.A1(_22521_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1714]),
    .A3(_23402_),
    .ZN(_26301_));
 AOI221_X4 _57543_ (.A(_26301_),
    .B1(_11025_),
    .B2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1616]),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1763]),
    .C2(_22078_),
    .ZN(_26302_));
 AND3_X1 _57544_ (.A1(_23083_),
    .A2(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2008]),
    .A3(_10939_),
    .ZN(_26303_));
 AOI221_X4 _57545_ (.A(_26303_),
    .B1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2106]),
    .B2(_10968_),
    .C1(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2155]),
    .C2(_23736_),
    .ZN(_26304_));
 AND4_X4 _57546_ (.A1(_26295_),
    .A2(_26300_),
    .A3(_26302_),
    .A4(_26304_),
    .ZN(_26305_));
 NAND4_X1 _57547_ (.A1(net5),
    .A2(_26285_),
    .A3(_26291_),
    .A4(_26305_),
    .ZN(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [48]));
 INV_X1 _57548_ (.A(_21259_),
    .ZN(_26306_));
 OR2_X1 _57549_ (.A1(_26306_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.w_addr_i ),
    .ZN(_26307_));
 BUF_X4 _57550_ (.A(_26307_),
    .Z(_26308_));
 BUF_X8 _57551_ (.A(_26308_),
    .Z(_26309_));
 MUX2_X1 _57552_ (.A(lce_cmd_i[0]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [0]),
    .S(_26309_),
    .Z(_05408_));
 MUX2_X1 _57553_ (.A(lce_cmd_i[1]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [1]),
    .S(_26309_),
    .Z(_05424_));
 MUX2_X1 _57554_ (.A(lce_cmd_i[2]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [2]),
    .S(_26309_),
    .Z(_05435_));
 MUX2_X1 _57555_ (.A(lce_cmd_i[3]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [3]),
    .S(_26309_),
    .Z(_05446_));
 MUX2_X1 _57556_ (.A(lce_cmd_i[4]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [4]),
    .S(_26309_),
    .Z(_05457_));
 MUX2_X1 _57557_ (.A(lce_cmd_i[5]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [5]),
    .S(_26309_),
    .Z(_05467_));
 MUX2_X1 _57558_ (.A(lce_cmd_i[6]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [6]),
    .S(_26309_),
    .Z(_05478_));
 MUX2_X1 _57559_ (.A(lce_cmd_i[7]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [7]),
    .S(_26309_),
    .Z(_05489_));
 MUX2_X1 _57560_ (.A(lce_cmd_i[8]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [8]),
    .S(_26309_),
    .Z(_05500_));
 MUX2_X1 _57561_ (.A(lce_cmd_i[9]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [9]),
    .S(_26309_),
    .Z(_05511_));
 BUF_X8 _57562_ (.A(_26308_),
    .Z(_26310_));
 MUX2_X1 _57563_ (.A(lce_cmd_i[10]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [10]),
    .S(_26310_),
    .Z(_05414_));
 MUX2_X1 _57564_ (.A(lce_cmd_i[11]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [11]),
    .S(_26310_),
    .Z(_05415_));
 MUX2_X1 _57565_ (.A(lce_cmd_i[12]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [12]),
    .S(_26310_),
    .Z(_05416_));
 MUX2_X1 _57566_ (.A(lce_cmd_i[13]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [13]),
    .S(_26310_),
    .Z(_05417_));
 MUX2_X1 _57567_ (.A(lce_cmd_i[14]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [14]),
    .S(_26310_),
    .Z(_05418_));
 MUX2_X1 _57568_ (.A(lce_cmd_i[15]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [15]),
    .S(_26310_),
    .Z(_05419_));
 MUX2_X1 _57569_ (.A(lce_cmd_i[16]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [16]),
    .S(_26310_),
    .Z(_05420_));
 MUX2_X1 _57570_ (.A(lce_cmd_i[17]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [17]),
    .S(_26310_),
    .Z(_05421_));
 MUX2_X1 _57571_ (.A(lce_cmd_i[18]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [18]),
    .S(_26310_),
    .Z(_05422_));
 MUX2_X1 _57572_ (.A(lce_cmd_i[19]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [19]),
    .S(_26310_),
    .Z(_05423_));
 BUF_X8 _57573_ (.A(_26308_),
    .Z(_26311_));
 MUX2_X1 _57574_ (.A(lce_cmd_i[20]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [20]),
    .S(_26311_),
    .Z(_05425_));
 MUX2_X1 _57575_ (.A(lce_cmd_i[21]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [21]),
    .S(_26311_),
    .Z(_05426_));
 MUX2_X1 _57576_ (.A(lce_cmd_i[22]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [22]),
    .S(_26311_),
    .Z(_05427_));
 MUX2_X1 _57577_ (.A(lce_cmd_i[23]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [23]),
    .S(_26311_),
    .Z(_05428_));
 MUX2_X1 _57578_ (.A(lce_cmd_i[24]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [24]),
    .S(_26311_),
    .Z(_05429_));
 MUX2_X1 _57579_ (.A(lce_cmd_i[25]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [25]),
    .S(_26311_),
    .Z(_05430_));
 MUX2_X1 _57580_ (.A(lce_cmd_i[26]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [26]),
    .S(_26311_),
    .Z(_05431_));
 MUX2_X1 _57581_ (.A(lce_cmd_i[27]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [27]),
    .S(_26311_),
    .Z(_05432_));
 MUX2_X1 _57582_ (.A(lce_cmd_i[28]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [28]),
    .S(_26311_),
    .Z(_05433_));
 MUX2_X1 _57583_ (.A(lce_cmd_i[29]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [29]),
    .S(_26311_),
    .Z(_05434_));
 BUF_X8 _57584_ (.A(_26308_),
    .Z(_26312_));
 MUX2_X1 _57585_ (.A(lce_cmd_i[30]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [30]),
    .S(_26312_),
    .Z(_05436_));
 MUX2_X1 _57586_ (.A(lce_cmd_i[31]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [31]),
    .S(_26312_),
    .Z(_05437_));
 MUX2_X1 _57587_ (.A(lce_cmd_i[32]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [32]),
    .S(_26312_),
    .Z(_05438_));
 MUX2_X1 _57588_ (.A(lce_cmd_i[33]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [33]),
    .S(_26312_),
    .Z(_05439_));
 MUX2_X1 _57589_ (.A(lce_cmd_i[34]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [34]),
    .S(_26312_),
    .Z(_05440_));
 MUX2_X1 _57590_ (.A(lce_cmd_i[35]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [35]),
    .S(_26312_),
    .Z(_05441_));
 MUX2_X1 _57591_ (.A(lce_cmd_i[36]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [36]),
    .S(_26312_),
    .Z(_05442_));
 MUX2_X1 _57592_ (.A(lce_cmd_i[37]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [37]),
    .S(_26312_),
    .Z(_05443_));
 MUX2_X1 _57593_ (.A(lce_cmd_i[38]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [38]),
    .S(_26312_),
    .Z(_05444_));
 MUX2_X1 _57594_ (.A(lce_cmd_i[39]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [39]),
    .S(_26312_),
    .Z(_05445_));
 BUF_X8 _57595_ (.A(_26308_),
    .Z(_26313_));
 MUX2_X1 _57596_ (.A(lce_cmd_i[40]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [40]),
    .S(_26313_),
    .Z(_05447_));
 MUX2_X1 _57597_ (.A(lce_cmd_i[41]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [41]),
    .S(_26313_),
    .Z(_05448_));
 MUX2_X1 _57598_ (.A(lce_cmd_i[42]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [42]),
    .S(_26313_),
    .Z(_05449_));
 MUX2_X1 _57599_ (.A(lce_cmd_i[43]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [43]),
    .S(_26313_),
    .Z(_05450_));
 MUX2_X1 _57600_ (.A(lce_cmd_i[44]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [44]),
    .S(_26313_),
    .Z(_05451_));
 MUX2_X1 _57601_ (.A(lce_cmd_i[45]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [45]),
    .S(_26313_),
    .Z(_05452_));
 MUX2_X1 _57602_ (.A(lce_cmd_i[46]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [46]),
    .S(_26313_),
    .Z(_05453_));
 MUX2_X1 _57603_ (.A(lce_cmd_i[47]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [47]),
    .S(_26313_),
    .Z(_05454_));
 MUX2_X1 _57604_ (.A(lce_cmd_i[48]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [48]),
    .S(_26313_),
    .Z(_05455_));
 MUX2_X1 _57605_ (.A(lce_cmd_i[49]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [49]),
    .S(_26313_),
    .Z(_05456_));
 MUX2_X1 _57606_ (.A(lce_cmd_i[50]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [50]),
    .S(_26308_),
    .Z(_05458_));
 MUX2_X1 _57607_ (.A(lce_cmd_i[51]),
    .B(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [51]),
    .S(_26308_),
    .Z(_05459_));
 MUX2_X1 _57608_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [53]),
    .B(lce_cmd_i[0]),
    .S(_21262_),
    .Z(_05460_));
 MUX2_X1 _57609_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [54]),
    .B(lce_cmd_i[1]),
    .S(_21262_),
    .Z(_05461_));
 MUX2_X1 _57610_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [55]),
    .B(lce_cmd_i[2]),
    .S(_21262_),
    .Z(_05462_));
 MUX2_X1 _57611_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [56]),
    .B(lce_cmd_i[3]),
    .S(_21262_),
    .Z(_05463_));
 MUX2_X1 _57612_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [57]),
    .B(lce_cmd_i[4]),
    .S(_21262_),
    .Z(_05464_));
 MUX2_X1 _57613_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [58]),
    .B(lce_cmd_i[5]),
    .S(_21262_),
    .Z(_05465_));
 MUX2_X1 _57614_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [59]),
    .B(lce_cmd_i[6]),
    .S(_21262_),
    .Z(_05466_));
 MUX2_X1 _57615_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [60]),
    .B(lce_cmd_i[7]),
    .S(_21262_),
    .Z(_05468_));
 MUX2_X1 _57616_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [61]),
    .B(lce_cmd_i[8]),
    .S(_21262_),
    .Z(_05469_));
 BUF_X8 _57617_ (.A(_21261_),
    .Z(_26314_));
 MUX2_X1 _57618_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [62]),
    .B(lce_cmd_i[9]),
    .S(_26314_),
    .Z(_05470_));
 MUX2_X1 _57619_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [63]),
    .B(lce_cmd_i[10]),
    .S(_26314_),
    .Z(_05471_));
 MUX2_X1 _57620_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [64]),
    .B(lce_cmd_i[11]),
    .S(_26314_),
    .Z(_05472_));
 MUX2_X1 _57621_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [65]),
    .B(lce_cmd_i[12]),
    .S(_26314_),
    .Z(_05473_));
 MUX2_X1 _57622_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [66]),
    .B(lce_cmd_i[13]),
    .S(_26314_),
    .Z(_05474_));
 MUX2_X1 _57623_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [67]),
    .B(lce_cmd_i[14]),
    .S(_26314_),
    .Z(_05475_));
 MUX2_X1 _57624_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [68]),
    .B(lce_cmd_i[15]),
    .S(_26314_),
    .Z(_05476_));
 MUX2_X1 _57625_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [69]),
    .B(lce_cmd_i[16]),
    .S(_26314_),
    .Z(_05477_));
 MUX2_X1 _57626_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [70]),
    .B(lce_cmd_i[17]),
    .S(_26314_),
    .Z(_05479_));
 MUX2_X1 _57627_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [71]),
    .B(lce_cmd_i[18]),
    .S(_26314_),
    .Z(_05480_));
 BUF_X4 _57628_ (.A(_21261_),
    .Z(_26315_));
 MUX2_X1 _57629_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [72]),
    .B(lce_cmd_i[19]),
    .S(_26315_),
    .Z(_05481_));
 MUX2_X1 _57630_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [73]),
    .B(lce_cmd_i[20]),
    .S(_26315_),
    .Z(_05482_));
 MUX2_X1 _57631_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [74]),
    .B(lce_cmd_i[21]),
    .S(_26315_),
    .Z(_05483_));
 MUX2_X1 _57632_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [75]),
    .B(lce_cmd_i[22]),
    .S(_26315_),
    .Z(_05484_));
 MUX2_X1 _57633_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [76]),
    .B(lce_cmd_i[23]),
    .S(_26315_),
    .Z(_05485_));
 MUX2_X1 _57634_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [77]),
    .B(lce_cmd_i[24]),
    .S(_26315_),
    .Z(_05486_));
 MUX2_X1 _57635_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [78]),
    .B(lce_cmd_i[25]),
    .S(_26315_),
    .Z(_05487_));
 MUX2_X1 _57636_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [79]),
    .B(lce_cmd_i[26]),
    .S(_26315_),
    .Z(_05488_));
 MUX2_X1 _57637_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [80]),
    .B(lce_cmd_i[27]),
    .S(_26315_),
    .Z(_05490_));
 MUX2_X1 _57638_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [81]),
    .B(lce_cmd_i[28]),
    .S(_26315_),
    .Z(_05491_));
 BUF_X8 _57639_ (.A(_21261_),
    .Z(_26316_));
 MUX2_X1 _57640_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [82]),
    .B(lce_cmd_i[29]),
    .S(_26316_),
    .Z(_05492_));
 MUX2_X1 _57641_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [83]),
    .B(lce_cmd_i[30]),
    .S(_26316_),
    .Z(_05493_));
 MUX2_X1 _57642_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [84]),
    .B(lce_cmd_i[31]),
    .S(_26316_),
    .Z(_05494_));
 MUX2_X1 _57643_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [85]),
    .B(lce_cmd_i[32]),
    .S(_26316_),
    .Z(_05495_));
 MUX2_X1 _57644_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [86]),
    .B(lce_cmd_i[33]),
    .S(_26316_),
    .Z(_05496_));
 MUX2_X1 _57645_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [87]),
    .B(lce_cmd_i[34]),
    .S(_26316_),
    .Z(_05497_));
 MUX2_X1 _57646_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [88]),
    .B(lce_cmd_i[35]),
    .S(_26316_),
    .Z(_05498_));
 MUX2_X1 _57647_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [89]),
    .B(lce_cmd_i[36]),
    .S(_26316_),
    .Z(_05499_));
 MUX2_X1 _57648_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [90]),
    .B(lce_cmd_i[37]),
    .S(_26316_),
    .Z(_05501_));
 MUX2_X1 _57649_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [91]),
    .B(lce_cmd_i[38]),
    .S(_26316_),
    .Z(_05502_));
 BUF_X8 _57650_ (.A(_21261_),
    .Z(_26317_));
 MUX2_X1 _57651_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [92]),
    .B(lce_cmd_i[39]),
    .S(_26317_),
    .Z(_05503_));
 MUX2_X1 _57652_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [93]),
    .B(lce_cmd_i[40]),
    .S(_26317_),
    .Z(_05504_));
 MUX2_X1 _57653_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [94]),
    .B(lce_cmd_i[41]),
    .S(_26317_),
    .Z(_05505_));
 MUX2_X1 _57654_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [95]),
    .B(lce_cmd_i[42]),
    .S(_26317_),
    .Z(_05506_));
 MUX2_X1 _57655_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [96]),
    .B(lce_cmd_i[43]),
    .S(_26317_),
    .Z(_05507_));
 MUX2_X1 _57656_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [97]),
    .B(lce_cmd_i[44]),
    .S(_26317_),
    .Z(_05508_));
 MUX2_X1 _57657_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [98]),
    .B(lce_cmd_i[45]),
    .S(_26317_),
    .Z(_05509_));
 MUX2_X1 _57658_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [99]),
    .B(lce_cmd_i[46]),
    .S(_26317_),
    .Z(_05510_));
 MUX2_X1 _57659_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [100]),
    .B(lce_cmd_i[47]),
    .S(_26317_),
    .Z(_05409_));
 MUX2_X1 _57660_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [101]),
    .B(lce_cmd_i[48]),
    .S(_26317_),
    .Z(_05410_));
 MUX2_X1 _57661_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [102]),
    .B(lce_cmd_i[49]),
    .S(_21261_),
    .Z(_05411_));
 MUX2_X1 _57662_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [103]),
    .B(lce_cmd_i[50]),
    .S(_21261_),
    .Z(_05412_));
 MUX2_X1 _57663_ (.A(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [104]),
    .B(lce_cmd_i[51]),
    .S(_21261_),
    .Z(_05413_));
 AND2_X2 _57664_ (.A1(_21282_),
    .A2(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.w_addr_i ),
    .ZN(_26318_));
 BUF_X16 _57665_ (.A(_26318_),
    .Z(_26319_));
 BUF_X16 _57666_ (.A(_26319_),
    .Z(_26320_));
 BUF_X16 _57667_ (.A(_26320_),
    .Z(_26321_));
 MUX2_X1 _57668_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [521]),
    .B(lce_data_cmd_i[3]),
    .S(_26321_),
    .Z(_06018_));
 MUX2_X1 _57669_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [541]),
    .B(lce_data_cmd_i[23]),
    .S(_26321_),
    .Z(_06039_));
 MUX2_X1 _57670_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [542]),
    .B(lce_data_cmd_i[24]),
    .S(_26321_),
    .Z(_06040_));
 MUX2_X1 _57671_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [543]),
    .B(lce_data_cmd_i[25]),
    .S(_26321_),
    .Z(_06041_));
 MUX2_X1 _57672_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [544]),
    .B(lce_data_cmd_i[26]),
    .S(_26321_),
    .Z(_06042_));
 MUX2_X1 _57673_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [545]),
    .B(lce_data_cmd_i[27]),
    .S(_26321_),
    .Z(_06043_));
 MUX2_X1 _57674_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [546]),
    .B(lce_data_cmd_i[28]),
    .S(_26321_),
    .Z(_06044_));
 MUX2_X1 _57675_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [547]),
    .B(lce_data_cmd_i[29]),
    .S(_26321_),
    .Z(_06045_));
 MUX2_X1 _57676_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [548]),
    .B(lce_data_cmd_i[30]),
    .S(_26321_),
    .Z(_06046_));
 MUX2_X1 _57677_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [549]),
    .B(lce_data_cmd_i[31]),
    .S(_26321_),
    .Z(_06047_));
 BUF_X16 _57678_ (.A(_26320_),
    .Z(_26322_));
 MUX2_X1 _57679_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [550]),
    .B(lce_data_cmd_i[32]),
    .S(_26322_),
    .Z(_06049_));
 MUX2_X1 _57680_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [551]),
    .B(lce_data_cmd_i[33]),
    .S(_26322_),
    .Z(_06050_));
 MUX2_X1 _57681_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [552]),
    .B(lce_data_cmd_i[34]),
    .S(_26322_),
    .Z(_06051_));
 MUX2_X1 _57682_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [553]),
    .B(lce_data_cmd_i[35]),
    .S(_26322_),
    .Z(_06052_));
 MUX2_X1 _57683_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [554]),
    .B(lce_data_cmd_i[36]),
    .S(_26322_),
    .Z(_06053_));
 MUX2_X1 _57684_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [555]),
    .B(lce_data_cmd_i[37]),
    .S(_26322_),
    .Z(_06054_));
 MUX2_X1 _57685_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [556]),
    .B(lce_data_cmd_i[38]),
    .S(_26322_),
    .Z(_06055_));
 MUX2_X1 _57686_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [557]),
    .B(lce_data_cmd_i[39]),
    .S(_26322_),
    .Z(_06056_));
 MUX2_X1 _57687_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [558]),
    .B(lce_data_cmd_i[40]),
    .S(_26322_),
    .Z(_06057_));
 MUX2_X1 _57688_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [559]),
    .B(lce_data_cmd_i[41]),
    .S(_26322_),
    .Z(_06058_));
 BUF_X8 _57689_ (.A(_26320_),
    .Z(_26323_));
 MUX2_X1 _57690_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [560]),
    .B(lce_data_cmd_i[42]),
    .S(_26323_),
    .Z(_06060_));
 MUX2_X1 _57691_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [561]),
    .B(lce_data_cmd_i[43]),
    .S(_26323_),
    .Z(_06061_));
 MUX2_X1 _57692_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [562]),
    .B(lce_data_cmd_i[44]),
    .S(_26323_),
    .Z(_06062_));
 MUX2_X1 _57693_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [563]),
    .B(lce_data_cmd_i[45]),
    .S(_26323_),
    .Z(_06063_));
 MUX2_X1 _57694_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [564]),
    .B(lce_data_cmd_i[46]),
    .S(_26323_),
    .Z(_06064_));
 MUX2_X1 _57695_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [565]),
    .B(lce_data_cmd_i[47]),
    .S(_26323_),
    .Z(_06065_));
 MUX2_X1 _57696_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [566]),
    .B(lce_data_cmd_i[48]),
    .S(_26323_),
    .Z(_06066_));
 MUX2_X1 _57697_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [567]),
    .B(lce_data_cmd_i[49]),
    .S(_26323_),
    .Z(_06067_));
 MUX2_X1 _57698_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [568]),
    .B(lce_data_cmd_i[50]),
    .S(_26323_),
    .Z(_06068_));
 MUX2_X1 _57699_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [569]),
    .B(lce_data_cmd_i[51]),
    .S(_26323_),
    .Z(_06069_));
 BUF_X32 _57700_ (.A(_26319_),
    .Z(_26324_));
 BUF_X32 _57701_ (.A(_26324_),
    .Z(_26325_));
 BUF_X8 _57702_ (.A(_26325_),
    .Z(_26326_));
 MUX2_X1 _57703_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [570]),
    .B(lce_data_cmd_i[52]),
    .S(_26326_),
    .Z(_06071_));
 MUX2_X1 _57704_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [571]),
    .B(lce_data_cmd_i[53]),
    .S(_26326_),
    .Z(_06072_));
 MUX2_X1 _57705_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [572]),
    .B(lce_data_cmd_i[54]),
    .S(_26326_),
    .Z(_06073_));
 MUX2_X1 _57706_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [573]),
    .B(lce_data_cmd_i[55]),
    .S(_26326_),
    .Z(_06074_));
 MUX2_X1 _57707_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [574]),
    .B(lce_data_cmd_i[56]),
    .S(_26326_),
    .Z(_06075_));
 MUX2_X1 _57708_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [575]),
    .B(lce_data_cmd_i[57]),
    .S(_26326_),
    .Z(_06076_));
 MUX2_X1 _57709_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [576]),
    .B(lce_data_cmd_i[58]),
    .S(_26326_),
    .Z(_06077_));
 MUX2_X1 _57710_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [577]),
    .B(lce_data_cmd_i[59]),
    .S(_26326_),
    .Z(_06078_));
 MUX2_X1 _57711_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [578]),
    .B(lce_data_cmd_i[60]),
    .S(_26326_),
    .Z(_06079_));
 MUX2_X1 _57712_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [579]),
    .B(lce_data_cmd_i[61]),
    .S(_26326_),
    .Z(_06080_));
 BUF_X32 _57713_ (.A(_26325_),
    .Z(_26327_));
 MUX2_X1 _57714_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [580]),
    .B(lce_data_cmd_i[62]),
    .S(_26327_),
    .Z(_06082_));
 MUX2_X1 _57715_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [581]),
    .B(lce_data_cmd_i[63]),
    .S(_26327_),
    .Z(_06083_));
 MUX2_X1 _57716_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [582]),
    .B(lce_data_cmd_i[64]),
    .S(_26327_),
    .Z(_06084_));
 MUX2_X1 _57717_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [583]),
    .B(lce_data_cmd_i[65]),
    .S(_26327_),
    .Z(_06085_));
 MUX2_X1 _57718_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [584]),
    .B(lce_data_cmd_i[66]),
    .S(_26327_),
    .Z(_06086_));
 MUX2_X1 _57719_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [585]),
    .B(lce_data_cmd_i[67]),
    .S(_26327_),
    .Z(_06087_));
 MUX2_X1 _57720_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [586]),
    .B(lce_data_cmd_i[68]),
    .S(_26327_),
    .Z(_06088_));
 MUX2_X1 _57721_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [587]),
    .B(lce_data_cmd_i[69]),
    .S(_26327_),
    .Z(_06089_));
 MUX2_X1 _57722_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [588]),
    .B(lce_data_cmd_i[70]),
    .S(_26327_),
    .Z(_06090_));
 MUX2_X1 _57723_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [589]),
    .B(lce_data_cmd_i[71]),
    .S(_26327_),
    .Z(_06091_));
 BUF_X16 _57724_ (.A(_26325_),
    .Z(_26328_));
 MUX2_X1 _57725_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [590]),
    .B(lce_data_cmd_i[72]),
    .S(_26328_),
    .Z(_06093_));
 MUX2_X1 _57726_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [591]),
    .B(lce_data_cmd_i[73]),
    .S(_26328_),
    .Z(_06094_));
 MUX2_X1 _57727_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [592]),
    .B(lce_data_cmd_i[74]),
    .S(_26328_),
    .Z(_06095_));
 MUX2_X1 _57728_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [593]),
    .B(lce_data_cmd_i[75]),
    .S(_26328_),
    .Z(_06096_));
 MUX2_X1 _57729_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [594]),
    .B(lce_data_cmd_i[76]),
    .S(_26328_),
    .Z(_06097_));
 MUX2_X1 _57730_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [595]),
    .B(lce_data_cmd_i[77]),
    .S(_26328_),
    .Z(_06098_));
 MUX2_X1 _57731_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [596]),
    .B(lce_data_cmd_i[78]),
    .S(_26328_),
    .Z(_06099_));
 MUX2_X1 _57732_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [597]),
    .B(lce_data_cmd_i[79]),
    .S(_26328_),
    .Z(_06100_));
 MUX2_X1 _57733_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [598]),
    .B(lce_data_cmd_i[80]),
    .S(_26328_),
    .Z(_06101_));
 MUX2_X1 _57734_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [599]),
    .B(lce_data_cmd_i[81]),
    .S(_26328_),
    .Z(_06102_));
 BUF_X8 _57735_ (.A(_26325_),
    .Z(_26329_));
 MUX2_X1 _57736_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [600]),
    .B(lce_data_cmd_i[82]),
    .S(_26329_),
    .Z(_06104_));
 MUX2_X1 _57737_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [601]),
    .B(lce_data_cmd_i[83]),
    .S(_26329_),
    .Z(_06105_));
 MUX2_X1 _57738_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [602]),
    .B(lce_data_cmd_i[84]),
    .S(_26329_),
    .Z(_06106_));
 MUX2_X1 _57739_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [603]),
    .B(lce_data_cmd_i[85]),
    .S(_26329_),
    .Z(_06107_));
 MUX2_X1 _57740_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [604]),
    .B(lce_data_cmd_i[86]),
    .S(_26329_),
    .Z(_06108_));
 MUX2_X1 _57741_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [605]),
    .B(lce_data_cmd_i[87]),
    .S(_26329_),
    .Z(_06109_));
 MUX2_X1 _57742_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [606]),
    .B(lce_data_cmd_i[88]),
    .S(_26329_),
    .Z(_06110_));
 MUX2_X1 _57743_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [607]),
    .B(lce_data_cmd_i[89]),
    .S(_26329_),
    .Z(_06111_));
 MUX2_X1 _57744_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [608]),
    .B(lce_data_cmd_i[90]),
    .S(_26329_),
    .Z(_06112_));
 MUX2_X1 _57745_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [609]),
    .B(lce_data_cmd_i[91]),
    .S(_26329_),
    .Z(_06113_));
 BUF_X8 _57746_ (.A(_26325_),
    .Z(_26330_));
 MUX2_X1 _57747_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [610]),
    .B(lce_data_cmd_i[92]),
    .S(_26330_),
    .Z(_06115_));
 MUX2_X1 _57748_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [611]),
    .B(lce_data_cmd_i[93]),
    .S(_26330_),
    .Z(_06116_));
 MUX2_X1 _57749_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [612]),
    .B(lce_data_cmd_i[94]),
    .S(_26330_),
    .Z(_06117_));
 MUX2_X1 _57750_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [613]),
    .B(lce_data_cmd_i[95]),
    .S(_26330_),
    .Z(_06118_));
 MUX2_X1 _57751_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [614]),
    .B(lce_data_cmd_i[96]),
    .S(_26330_),
    .Z(_06119_));
 MUX2_X1 _57752_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [615]),
    .B(lce_data_cmd_i[97]),
    .S(_26330_),
    .Z(_06120_));
 MUX2_X1 _57753_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [616]),
    .B(lce_data_cmd_i[98]),
    .S(_26330_),
    .Z(_06121_));
 MUX2_X1 _57754_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [617]),
    .B(lce_data_cmd_i[99]),
    .S(_26330_),
    .Z(_06122_));
 MUX2_X1 _57755_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [618]),
    .B(lce_data_cmd_i[100]),
    .S(_26330_),
    .Z(_06123_));
 MUX2_X1 _57756_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [619]),
    .B(lce_data_cmd_i[101]),
    .S(_26330_),
    .Z(_06124_));
 BUF_X8 _57757_ (.A(_26325_),
    .Z(_26331_));
 MUX2_X1 _57758_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [620]),
    .B(lce_data_cmd_i[102]),
    .S(_26331_),
    .Z(_06126_));
 MUX2_X1 _57759_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [621]),
    .B(lce_data_cmd_i[103]),
    .S(_26331_),
    .Z(_06127_));
 MUX2_X1 _57760_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [622]),
    .B(lce_data_cmd_i[104]),
    .S(_26331_),
    .Z(_06128_));
 MUX2_X1 _57761_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [623]),
    .B(lce_data_cmd_i[105]),
    .S(_26331_),
    .Z(_06129_));
 MUX2_X1 _57762_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [624]),
    .B(lce_data_cmd_i[106]),
    .S(_26331_),
    .Z(_06130_));
 MUX2_X1 _57763_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [625]),
    .B(lce_data_cmd_i[107]),
    .S(_26331_),
    .Z(_06131_));
 MUX2_X1 _57764_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [626]),
    .B(lce_data_cmd_i[108]),
    .S(_26331_),
    .Z(_06132_));
 MUX2_X1 _57765_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [627]),
    .B(lce_data_cmd_i[109]),
    .S(_26331_),
    .Z(_06133_));
 MUX2_X1 _57766_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [628]),
    .B(lce_data_cmd_i[110]),
    .S(_26331_),
    .Z(_06134_));
 MUX2_X1 _57767_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [629]),
    .B(lce_data_cmd_i[111]),
    .S(_26331_),
    .Z(_06135_));
 BUF_X8 _57768_ (.A(_26325_),
    .Z(_26332_));
 MUX2_X1 _57769_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [630]),
    .B(lce_data_cmd_i[112]),
    .S(_26332_),
    .Z(_06137_));
 MUX2_X1 _57770_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [631]),
    .B(lce_data_cmd_i[113]),
    .S(_26332_),
    .Z(_06138_));
 MUX2_X1 _57771_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [632]),
    .B(lce_data_cmd_i[114]),
    .S(_26332_),
    .Z(_06139_));
 MUX2_X1 _57772_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [633]),
    .B(lce_data_cmd_i[115]),
    .S(_26332_),
    .Z(_06140_));
 MUX2_X1 _57773_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [634]),
    .B(lce_data_cmd_i[116]),
    .S(_26332_),
    .Z(_06141_));
 MUX2_X1 _57774_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [635]),
    .B(lce_data_cmd_i[117]),
    .S(_26332_),
    .Z(_06142_));
 MUX2_X1 _57775_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [636]),
    .B(lce_data_cmd_i[118]),
    .S(_26332_),
    .Z(_06143_));
 MUX2_X1 _57776_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [637]),
    .B(lce_data_cmd_i[119]),
    .S(_26332_),
    .Z(_06144_));
 MUX2_X1 _57777_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [638]),
    .B(lce_data_cmd_i[120]),
    .S(_26332_),
    .Z(_06145_));
 MUX2_X1 _57778_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [639]),
    .B(lce_data_cmd_i[121]),
    .S(_26332_),
    .Z(_06146_));
 BUF_X8 _57779_ (.A(_26325_),
    .Z(_26333_));
 MUX2_X1 _57780_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [518]),
    .B(lce_data_cmd_i[0]),
    .S(_26333_),
    .Z(_06014_));
 MUX2_X1 _57781_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [937]),
    .B(lce_data_cmd_i[419]),
    .S(_26333_),
    .Z(_06477_));
 MUX2_X1 _57782_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [938]),
    .B(lce_data_cmd_i[420]),
    .S(_26333_),
    .Z(_06478_));
 MUX2_X1 _57783_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [939]),
    .B(lce_data_cmd_i[421]),
    .S(_26333_),
    .Z(_06479_));
 MUX2_X1 _57784_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [940]),
    .B(lce_data_cmd_i[422]),
    .S(_26333_),
    .Z(_06481_));
 MUX2_X1 _57785_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [941]),
    .B(lce_data_cmd_i[423]),
    .S(_26333_),
    .Z(_06482_));
 MUX2_X1 _57786_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [942]),
    .B(lce_data_cmd_i[424]),
    .S(_26333_),
    .Z(_06483_));
 MUX2_X1 _57787_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [943]),
    .B(lce_data_cmd_i[425]),
    .S(_26333_),
    .Z(_06484_));
 MUX2_X1 _57788_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [944]),
    .B(lce_data_cmd_i[426]),
    .S(_26333_),
    .Z(_06485_));
 MUX2_X1 _57789_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [945]),
    .B(lce_data_cmd_i[427]),
    .S(_26333_),
    .Z(_06486_));
 BUF_X8 _57790_ (.A(_26325_),
    .Z(_26334_));
 MUX2_X1 _57791_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [946]),
    .B(lce_data_cmd_i[428]),
    .S(_26334_),
    .Z(_06487_));
 MUX2_X1 _57792_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [947]),
    .B(lce_data_cmd_i[429]),
    .S(_26334_),
    .Z(_06488_));
 MUX2_X1 _57793_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [948]),
    .B(lce_data_cmd_i[430]),
    .S(_26334_),
    .Z(_06489_));
 MUX2_X1 _57794_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [949]),
    .B(lce_data_cmd_i[431]),
    .S(_26334_),
    .Z(_06490_));
 MUX2_X1 _57795_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [950]),
    .B(lce_data_cmd_i[432]),
    .S(_26334_),
    .Z(_06492_));
 MUX2_X1 _57796_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [951]),
    .B(lce_data_cmd_i[433]),
    .S(_26334_),
    .Z(_06493_));
 MUX2_X1 _57797_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [952]),
    .B(lce_data_cmd_i[434]),
    .S(_26334_),
    .Z(_06494_));
 MUX2_X1 _57798_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [953]),
    .B(lce_data_cmd_i[435]),
    .S(_26334_),
    .Z(_06495_));
 MUX2_X1 _57799_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [954]),
    .B(lce_data_cmd_i[436]),
    .S(_26334_),
    .Z(_06496_));
 MUX2_X1 _57800_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [955]),
    .B(lce_data_cmd_i[437]),
    .S(_26334_),
    .Z(_06497_));
 BUF_X8 _57801_ (.A(_26325_),
    .Z(_26335_));
 MUX2_X1 _57802_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [956]),
    .B(lce_data_cmd_i[438]),
    .S(_26335_),
    .Z(_06498_));
 MUX2_X1 _57803_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [957]),
    .B(lce_data_cmd_i[439]),
    .S(_26335_),
    .Z(_06499_));
 MUX2_X1 _57804_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [958]),
    .B(lce_data_cmd_i[440]),
    .S(_26335_),
    .Z(_06500_));
 MUX2_X1 _57805_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [959]),
    .B(lce_data_cmd_i[441]),
    .S(_26335_),
    .Z(_06501_));
 MUX2_X1 _57806_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [960]),
    .B(lce_data_cmd_i[442]),
    .S(_26335_),
    .Z(_06503_));
 MUX2_X1 _57807_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [961]),
    .B(lce_data_cmd_i[443]),
    .S(_26335_),
    .Z(_06504_));
 MUX2_X1 _57808_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [962]),
    .B(lce_data_cmd_i[444]),
    .S(_26335_),
    .Z(_06505_));
 MUX2_X1 _57809_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [963]),
    .B(lce_data_cmd_i[445]),
    .S(_26335_),
    .Z(_06506_));
 MUX2_X1 _57810_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [964]),
    .B(lce_data_cmd_i[446]),
    .S(_26335_),
    .Z(_06507_));
 MUX2_X1 _57811_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [965]),
    .B(lce_data_cmd_i[447]),
    .S(_26335_),
    .Z(_06508_));
 BUF_X32 _57812_ (.A(_26324_),
    .Z(_26336_));
 BUF_X8 _57813_ (.A(_26336_),
    .Z(_26337_));
 MUX2_X1 _57814_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [966]),
    .B(lce_data_cmd_i[448]),
    .S(_26337_),
    .Z(_06509_));
 MUX2_X1 _57815_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [967]),
    .B(lce_data_cmd_i[449]),
    .S(_26337_),
    .Z(_06510_));
 MUX2_X1 _57816_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [968]),
    .B(lce_data_cmd_i[450]),
    .S(_26337_),
    .Z(_06511_));
 MUX2_X1 _57817_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [969]),
    .B(lce_data_cmd_i[451]),
    .S(_26337_),
    .Z(_06512_));
 MUX2_X1 _57818_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [970]),
    .B(lce_data_cmd_i[452]),
    .S(_26337_),
    .Z(_06514_));
 MUX2_X1 _57819_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [971]),
    .B(lce_data_cmd_i[453]),
    .S(_26337_),
    .Z(_06515_));
 MUX2_X1 _57820_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [972]),
    .B(lce_data_cmd_i[454]),
    .S(_26337_),
    .Z(_06516_));
 MUX2_X1 _57821_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [973]),
    .B(lce_data_cmd_i[455]),
    .S(_26337_),
    .Z(_06517_));
 MUX2_X1 _57822_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [974]),
    .B(lce_data_cmd_i[456]),
    .S(_26337_),
    .Z(_06518_));
 MUX2_X1 _57823_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [975]),
    .B(lce_data_cmd_i[457]),
    .S(_26337_),
    .Z(_06519_));
 BUF_X8 _57824_ (.A(_26336_),
    .Z(_26338_));
 MUX2_X1 _57825_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [976]),
    .B(lce_data_cmd_i[458]),
    .S(_26338_),
    .Z(_06520_));
 MUX2_X1 _57826_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [977]),
    .B(lce_data_cmd_i[459]),
    .S(_26338_),
    .Z(_06521_));
 MUX2_X1 _57827_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [978]),
    .B(lce_data_cmd_i[460]),
    .S(_26338_),
    .Z(_06522_));
 MUX2_X1 _57828_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [979]),
    .B(lce_data_cmd_i[461]),
    .S(_26338_),
    .Z(_06523_));
 MUX2_X1 _57829_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [980]),
    .B(lce_data_cmd_i[462]),
    .S(_26338_),
    .Z(_06525_));
 MUX2_X1 _57830_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [981]),
    .B(lce_data_cmd_i[463]),
    .S(_26338_),
    .Z(_06526_));
 MUX2_X1 _57831_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [982]),
    .B(lce_data_cmd_i[464]),
    .S(_26338_),
    .Z(_06527_));
 MUX2_X1 _57832_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [983]),
    .B(lce_data_cmd_i[465]),
    .S(_26338_),
    .Z(_06528_));
 MUX2_X1 _57833_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [984]),
    .B(lce_data_cmd_i[466]),
    .S(_26338_),
    .Z(_06529_));
 MUX2_X1 _57834_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [985]),
    .B(lce_data_cmd_i[467]),
    .S(_26338_),
    .Z(_06530_));
 BUF_X4 _57835_ (.A(_26336_),
    .Z(_26339_));
 MUX2_X1 _57836_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [986]),
    .B(lce_data_cmd_i[468]),
    .S(_26339_),
    .Z(_06531_));
 MUX2_X1 _57837_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [987]),
    .B(lce_data_cmd_i[469]),
    .S(_26339_),
    .Z(_06532_));
 MUX2_X1 _57838_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [988]),
    .B(lce_data_cmd_i[470]),
    .S(_26339_),
    .Z(_06533_));
 MUX2_X1 _57839_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [989]),
    .B(lce_data_cmd_i[471]),
    .S(_26339_),
    .Z(_06534_));
 MUX2_X1 _57840_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [990]),
    .B(lce_data_cmd_i[472]),
    .S(_26339_),
    .Z(_06536_));
 MUX2_X1 _57841_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [991]),
    .B(lce_data_cmd_i[473]),
    .S(_26339_),
    .Z(_06537_));
 MUX2_X1 _57842_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [992]),
    .B(lce_data_cmd_i[474]),
    .S(_26339_),
    .Z(_06538_));
 MUX2_X1 _57843_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [993]),
    .B(lce_data_cmd_i[475]),
    .S(_26339_),
    .Z(_06539_));
 MUX2_X1 _57844_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [994]),
    .B(lce_data_cmd_i[476]),
    .S(_26339_),
    .Z(_06540_));
 MUX2_X1 _57845_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [995]),
    .B(lce_data_cmd_i[477]),
    .S(_26339_),
    .Z(_06541_));
 BUF_X8 _57846_ (.A(_26336_),
    .Z(_26340_));
 MUX2_X1 _57847_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [996]),
    .B(lce_data_cmd_i[478]),
    .S(_26340_),
    .Z(_06542_));
 MUX2_X1 _57848_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [997]),
    .B(lce_data_cmd_i[479]),
    .S(_26340_),
    .Z(_06543_));
 MUX2_X1 _57849_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [998]),
    .B(lce_data_cmd_i[480]),
    .S(_26340_),
    .Z(_06544_));
 MUX2_X1 _57850_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [999]),
    .B(lce_data_cmd_i[481]),
    .S(_26340_),
    .Z(_06545_));
 MUX2_X1 _57851_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1000]),
    .B(lce_data_cmd_i[482]),
    .S(_26340_),
    .Z(_05515_));
 MUX2_X1 _57852_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1001]),
    .B(lce_data_cmd_i[483]),
    .S(_26340_),
    .Z(_05516_));
 MUX2_X1 _57853_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1002]),
    .B(lce_data_cmd_i[484]),
    .S(_26340_),
    .Z(_05517_));
 MUX2_X1 _57854_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1003]),
    .B(lce_data_cmd_i[485]),
    .S(_26340_),
    .Z(_05518_));
 MUX2_X1 _57855_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1004]),
    .B(lce_data_cmd_i[486]),
    .S(_26340_),
    .Z(_05519_));
 MUX2_X1 _57856_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1005]),
    .B(lce_data_cmd_i[487]),
    .S(_26340_),
    .Z(_05520_));
 BUF_X8 _57857_ (.A(_26336_),
    .Z(_26341_));
 MUX2_X1 _57858_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1006]),
    .B(lce_data_cmd_i[488]),
    .S(_26341_),
    .Z(_05521_));
 MUX2_X1 _57859_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1007]),
    .B(lce_data_cmd_i[489]),
    .S(_26341_),
    .Z(_05522_));
 MUX2_X1 _57860_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1008]),
    .B(lce_data_cmd_i[490]),
    .S(_26341_),
    .Z(_05523_));
 MUX2_X1 _57861_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1009]),
    .B(lce_data_cmd_i[491]),
    .S(_26341_),
    .Z(_05524_));
 MUX2_X1 _57862_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1010]),
    .B(lce_data_cmd_i[492]),
    .S(_26341_),
    .Z(_05526_));
 MUX2_X1 _57863_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1011]),
    .B(lce_data_cmd_i[493]),
    .S(_26341_),
    .Z(_05527_));
 MUX2_X1 _57864_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1012]),
    .B(lce_data_cmd_i[494]),
    .S(_26341_),
    .Z(_05528_));
 MUX2_X1 _57865_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1013]),
    .B(lce_data_cmd_i[495]),
    .S(_26341_),
    .Z(_05529_));
 MUX2_X1 _57866_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1014]),
    .B(lce_data_cmd_i[496]),
    .S(_26341_),
    .Z(_05530_));
 MUX2_X1 _57867_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1015]),
    .B(lce_data_cmd_i[497]),
    .S(_26341_),
    .Z(_05531_));
 BUF_X8 _57868_ (.A(_26336_),
    .Z(_26342_));
 MUX2_X1 _57869_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1016]),
    .B(lce_data_cmd_i[498]),
    .S(_26342_),
    .Z(_05532_));
 MUX2_X1 _57870_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1017]),
    .B(lce_data_cmd_i[499]),
    .S(_26342_),
    .Z(_05533_));
 MUX2_X1 _57871_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1018]),
    .B(lce_data_cmd_i[500]),
    .S(_26342_),
    .Z(_05534_));
 MUX2_X1 _57872_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1019]),
    .B(lce_data_cmd_i[501]),
    .S(_26342_),
    .Z(_05535_));
 MUX2_X1 _57873_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1020]),
    .B(lce_data_cmd_i[502]),
    .S(_26342_),
    .Z(_05537_));
 MUX2_X1 _57874_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1021]),
    .B(lce_data_cmd_i[503]),
    .S(_26342_),
    .Z(_05538_));
 MUX2_X1 _57875_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1022]),
    .B(lce_data_cmd_i[504]),
    .S(_26342_),
    .Z(_05539_));
 MUX2_X1 _57876_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1023]),
    .B(lce_data_cmd_i[505]),
    .S(_26342_),
    .Z(_05540_));
 MUX2_X1 _57877_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1024]),
    .B(lce_data_cmd_i[506]),
    .S(_26342_),
    .Z(_05541_));
 MUX2_X1 _57878_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1025]),
    .B(lce_data_cmd_i[507]),
    .S(_26342_),
    .Z(_05542_));
 BUF_X8 _57879_ (.A(_26336_),
    .Z(_26343_));
 MUX2_X1 _57880_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1026]),
    .B(lce_data_cmd_i[508]),
    .S(_26343_),
    .Z(_05543_));
 MUX2_X1 _57881_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1027]),
    .B(lce_data_cmd_i[509]),
    .S(_26343_),
    .Z(_05544_));
 MUX2_X1 _57882_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1028]),
    .B(lce_data_cmd_i[510]),
    .S(_26343_),
    .Z(_05545_));
 MUX2_X1 _57883_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1029]),
    .B(lce_data_cmd_i[511]),
    .S(_26343_),
    .Z(_05546_));
 MUX2_X1 _57884_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1030]),
    .B(lce_data_cmd_i[512]),
    .S(_26343_),
    .Z(_05548_));
 MUX2_X1 _57885_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1031]),
    .B(lce_data_cmd_i[513]),
    .S(_26343_),
    .Z(_05549_));
 MUX2_X1 _57886_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1032]),
    .B(lce_data_cmd_i[514]),
    .S(_26343_),
    .Z(_05550_));
 MUX2_X1 _57887_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1033]),
    .B(lce_data_cmd_i[515]),
    .S(_26343_),
    .Z(_05551_));
 MUX2_X1 _57888_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1034]),
    .B(lce_data_cmd_i[516]),
    .S(_26343_),
    .Z(_05552_));
 MUX2_X1 _57889_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1035]),
    .B(lce_data_cmd_i[517]),
    .S(_26343_),
    .Z(_05553_));
 BUF_X8 _57890_ (.A(_26336_),
    .Z(_26344_));
 MUX2_X1 _57891_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [519]),
    .B(lce_data_cmd_i[1]),
    .S(_26344_),
    .Z(_06015_));
 MUX2_X1 _57892_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [838]),
    .B(lce_data_cmd_i[320]),
    .S(_26344_),
    .Z(_06367_));
 MUX2_X1 _57893_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [839]),
    .B(lce_data_cmd_i[321]),
    .S(_26344_),
    .Z(_06368_));
 MUX2_X1 _57894_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [840]),
    .B(lce_data_cmd_i[322]),
    .S(_26344_),
    .Z(_06370_));
 MUX2_X1 _57895_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [841]),
    .B(lce_data_cmd_i[323]),
    .S(_26344_),
    .Z(_06371_));
 MUX2_X1 _57896_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [842]),
    .B(lce_data_cmd_i[324]),
    .S(_26344_),
    .Z(_06372_));
 MUX2_X1 _57897_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [843]),
    .B(lce_data_cmd_i[325]),
    .S(_26344_),
    .Z(_06373_));
 MUX2_X1 _57898_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [844]),
    .B(lce_data_cmd_i[326]),
    .S(_26344_),
    .Z(_06374_));
 MUX2_X1 _57899_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [845]),
    .B(lce_data_cmd_i[327]),
    .S(_26344_),
    .Z(_06375_));
 MUX2_X1 _57900_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [846]),
    .B(lce_data_cmd_i[328]),
    .S(_26344_),
    .Z(_06376_));
 BUF_X8 _57901_ (.A(_26336_),
    .Z(_26345_));
 MUX2_X1 _57902_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [847]),
    .B(lce_data_cmd_i[329]),
    .S(_26345_),
    .Z(_06377_));
 MUX2_X1 _57903_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [848]),
    .B(lce_data_cmd_i[330]),
    .S(_26345_),
    .Z(_06378_));
 MUX2_X1 _57904_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [849]),
    .B(lce_data_cmd_i[331]),
    .S(_26345_),
    .Z(_06379_));
 MUX2_X1 _57905_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [850]),
    .B(lce_data_cmd_i[332]),
    .S(_26345_),
    .Z(_06381_));
 MUX2_X1 _57906_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [851]),
    .B(lce_data_cmd_i[333]),
    .S(_26345_),
    .Z(_06382_));
 MUX2_X1 _57907_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [852]),
    .B(lce_data_cmd_i[334]),
    .S(_26345_),
    .Z(_06383_));
 MUX2_X1 _57908_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [853]),
    .B(lce_data_cmd_i[335]),
    .S(_26345_),
    .Z(_06384_));
 MUX2_X1 _57909_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [854]),
    .B(lce_data_cmd_i[336]),
    .S(_26345_),
    .Z(_06385_));
 MUX2_X1 _57910_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [855]),
    .B(lce_data_cmd_i[337]),
    .S(_26345_),
    .Z(_06386_));
 MUX2_X1 _57911_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [856]),
    .B(lce_data_cmd_i[338]),
    .S(_26345_),
    .Z(_06387_));
 BUF_X8 _57912_ (.A(_26336_),
    .Z(_26346_));
 MUX2_X1 _57913_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [857]),
    .B(lce_data_cmd_i[339]),
    .S(_26346_),
    .Z(_06388_));
 MUX2_X1 _57914_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [858]),
    .B(lce_data_cmd_i[340]),
    .S(_26346_),
    .Z(_06389_));
 MUX2_X1 _57915_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [859]),
    .B(lce_data_cmd_i[341]),
    .S(_26346_),
    .Z(_06390_));
 MUX2_X1 _57916_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [860]),
    .B(lce_data_cmd_i[342]),
    .S(_26346_),
    .Z(_06392_));
 MUX2_X1 _57917_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [861]),
    .B(lce_data_cmd_i[343]),
    .S(_26346_),
    .Z(_06393_));
 MUX2_X1 _57918_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [862]),
    .B(lce_data_cmd_i[344]),
    .S(_26346_),
    .Z(_06394_));
 MUX2_X1 _57919_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [863]),
    .B(lce_data_cmd_i[345]),
    .S(_26346_),
    .Z(_06395_));
 MUX2_X1 _57920_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [864]),
    .B(lce_data_cmd_i[346]),
    .S(_26346_),
    .Z(_06396_));
 MUX2_X1 _57921_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [865]),
    .B(lce_data_cmd_i[347]),
    .S(_26346_),
    .Z(_06397_));
 MUX2_X1 _57922_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [866]),
    .B(lce_data_cmd_i[348]),
    .S(_26346_),
    .Z(_06398_));
 BUF_X32 _57923_ (.A(_26319_),
    .Z(_26347_));
 BUF_X8 _57924_ (.A(_26347_),
    .Z(_26348_));
 MUX2_X1 _57925_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [867]),
    .B(lce_data_cmd_i[349]),
    .S(_26348_),
    .Z(_06399_));
 MUX2_X1 _57926_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [868]),
    .B(lce_data_cmd_i[350]),
    .S(_26348_),
    .Z(_06400_));
 MUX2_X1 _57927_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [869]),
    .B(lce_data_cmd_i[351]),
    .S(_26348_),
    .Z(_06401_));
 MUX2_X1 _57928_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [870]),
    .B(lce_data_cmd_i[352]),
    .S(_26348_),
    .Z(_06403_));
 MUX2_X1 _57929_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [871]),
    .B(lce_data_cmd_i[353]),
    .S(_26348_),
    .Z(_06404_));
 MUX2_X1 _57930_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [872]),
    .B(lce_data_cmd_i[354]),
    .S(_26348_),
    .Z(_06405_));
 MUX2_X1 _57931_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [873]),
    .B(lce_data_cmd_i[355]),
    .S(_26348_),
    .Z(_06406_));
 MUX2_X1 _57932_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [874]),
    .B(lce_data_cmd_i[356]),
    .S(_26348_),
    .Z(_06407_));
 MUX2_X1 _57933_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [875]),
    .B(lce_data_cmd_i[357]),
    .S(_26348_),
    .Z(_06408_));
 MUX2_X1 _57934_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [876]),
    .B(lce_data_cmd_i[358]),
    .S(_26348_),
    .Z(_06409_));
 BUF_X8 _57935_ (.A(_26347_),
    .Z(_26349_));
 MUX2_X1 _57936_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [877]),
    .B(lce_data_cmd_i[359]),
    .S(_26349_),
    .Z(_06410_));
 MUX2_X1 _57937_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [878]),
    .B(lce_data_cmd_i[360]),
    .S(_26349_),
    .Z(_06411_));
 MUX2_X1 _57938_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [879]),
    .B(lce_data_cmd_i[361]),
    .S(_26349_),
    .Z(_06412_));
 MUX2_X1 _57939_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [880]),
    .B(lce_data_cmd_i[362]),
    .S(_26349_),
    .Z(_06414_));
 MUX2_X1 _57940_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [881]),
    .B(lce_data_cmd_i[363]),
    .S(_26349_),
    .Z(_06415_));
 MUX2_X1 _57941_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [882]),
    .B(lce_data_cmd_i[364]),
    .S(_26349_),
    .Z(_06416_));
 MUX2_X1 _57942_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [883]),
    .B(lce_data_cmd_i[365]),
    .S(_26349_),
    .Z(_06417_));
 MUX2_X1 _57943_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [884]),
    .B(lce_data_cmd_i[366]),
    .S(_26349_),
    .Z(_06418_));
 MUX2_X1 _57944_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [885]),
    .B(lce_data_cmd_i[367]),
    .S(_26349_),
    .Z(_06419_));
 MUX2_X1 _57945_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [886]),
    .B(lce_data_cmd_i[368]),
    .S(_26349_),
    .Z(_06420_));
 BUF_X8 _57946_ (.A(_26347_),
    .Z(_26350_));
 MUX2_X1 _57947_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [887]),
    .B(lce_data_cmd_i[369]),
    .S(_26350_),
    .Z(_06421_));
 MUX2_X1 _57948_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [888]),
    .B(lce_data_cmd_i[370]),
    .S(_26350_),
    .Z(_06422_));
 MUX2_X1 _57949_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [889]),
    .B(lce_data_cmd_i[371]),
    .S(_26350_),
    .Z(_06423_));
 MUX2_X1 _57950_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [890]),
    .B(lce_data_cmd_i[372]),
    .S(_26350_),
    .Z(_06425_));
 MUX2_X1 _57951_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [891]),
    .B(lce_data_cmd_i[373]),
    .S(_26350_),
    .Z(_06426_));
 MUX2_X1 _57952_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [892]),
    .B(lce_data_cmd_i[374]),
    .S(_26350_),
    .Z(_06427_));
 MUX2_X1 _57953_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [893]),
    .B(lce_data_cmd_i[375]),
    .S(_26350_),
    .Z(_06428_));
 MUX2_X1 _57954_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [894]),
    .B(lce_data_cmd_i[376]),
    .S(_26350_),
    .Z(_06429_));
 MUX2_X1 _57955_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [895]),
    .B(lce_data_cmd_i[377]),
    .S(_26350_),
    .Z(_06430_));
 MUX2_X1 _57956_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [896]),
    .B(lce_data_cmd_i[378]),
    .S(_26350_),
    .Z(_06431_));
 BUF_X8 _57957_ (.A(_26347_),
    .Z(_26351_));
 MUX2_X1 _57958_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [897]),
    .B(lce_data_cmd_i[379]),
    .S(_26351_),
    .Z(_06432_));
 MUX2_X1 _57959_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [898]),
    .B(lce_data_cmd_i[380]),
    .S(_26351_),
    .Z(_06433_));
 MUX2_X1 _57960_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [899]),
    .B(lce_data_cmd_i[381]),
    .S(_26351_),
    .Z(_06434_));
 MUX2_X1 _57961_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [900]),
    .B(lce_data_cmd_i[382]),
    .S(_26351_),
    .Z(_06437_));
 MUX2_X1 _57962_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [901]),
    .B(lce_data_cmd_i[383]),
    .S(_26351_),
    .Z(_06438_));
 MUX2_X1 _57963_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [902]),
    .B(lce_data_cmd_i[384]),
    .S(_26351_),
    .Z(_06439_));
 MUX2_X1 _57964_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [903]),
    .B(lce_data_cmd_i[385]),
    .S(_26351_),
    .Z(_06440_));
 MUX2_X1 _57965_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [904]),
    .B(lce_data_cmd_i[386]),
    .S(_26351_),
    .Z(_06441_));
 MUX2_X1 _57966_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [905]),
    .B(lce_data_cmd_i[387]),
    .S(_26351_),
    .Z(_06442_));
 MUX2_X1 _57967_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [906]),
    .B(lce_data_cmd_i[388]),
    .S(_26351_),
    .Z(_06443_));
 BUF_X16 _57968_ (.A(_26347_),
    .Z(_26352_));
 MUX2_X1 _57969_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [907]),
    .B(lce_data_cmd_i[389]),
    .S(_26352_),
    .Z(_06444_));
 MUX2_X1 _57970_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [908]),
    .B(lce_data_cmd_i[390]),
    .S(_26352_),
    .Z(_06445_));
 MUX2_X1 _57971_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [909]),
    .B(lce_data_cmd_i[391]),
    .S(_26352_),
    .Z(_06446_));
 MUX2_X1 _57972_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [910]),
    .B(lce_data_cmd_i[392]),
    .S(_26352_),
    .Z(_06448_));
 MUX2_X1 _57973_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [911]),
    .B(lce_data_cmd_i[393]),
    .S(_26352_),
    .Z(_06449_));
 MUX2_X1 _57974_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [912]),
    .B(lce_data_cmd_i[394]),
    .S(_26352_),
    .Z(_06450_));
 MUX2_X1 _57975_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [913]),
    .B(lce_data_cmd_i[395]),
    .S(_26352_),
    .Z(_06451_));
 MUX2_X1 _57976_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [914]),
    .B(lce_data_cmd_i[396]),
    .S(_26352_),
    .Z(_06452_));
 MUX2_X1 _57977_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [915]),
    .B(lce_data_cmd_i[397]),
    .S(_26352_),
    .Z(_06453_));
 MUX2_X1 _57978_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [916]),
    .B(lce_data_cmd_i[398]),
    .S(_26352_),
    .Z(_06454_));
 BUF_X8 _57979_ (.A(_26347_),
    .Z(_26353_));
 MUX2_X1 _57980_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [917]),
    .B(lce_data_cmd_i[399]),
    .S(_26353_),
    .Z(_06455_));
 MUX2_X1 _57981_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [918]),
    .B(lce_data_cmd_i[400]),
    .S(_26353_),
    .Z(_06456_));
 MUX2_X1 _57982_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [919]),
    .B(lce_data_cmd_i[401]),
    .S(_26353_),
    .Z(_06457_));
 MUX2_X1 _57983_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [920]),
    .B(lce_data_cmd_i[402]),
    .S(_26353_),
    .Z(_06459_));
 MUX2_X1 _57984_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [921]),
    .B(lce_data_cmd_i[403]),
    .S(_26353_),
    .Z(_06460_));
 MUX2_X1 _57985_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [922]),
    .B(lce_data_cmd_i[404]),
    .S(_26353_),
    .Z(_06461_));
 MUX2_X1 _57986_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [923]),
    .B(lce_data_cmd_i[405]),
    .S(_26353_),
    .Z(_06462_));
 MUX2_X1 _57987_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [924]),
    .B(lce_data_cmd_i[406]),
    .S(_26353_),
    .Z(_06463_));
 MUX2_X1 _57988_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [925]),
    .B(lce_data_cmd_i[407]),
    .S(_26353_),
    .Z(_06464_));
 MUX2_X1 _57989_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [926]),
    .B(lce_data_cmd_i[408]),
    .S(_26353_),
    .Z(_06465_));
 BUF_X4 _57990_ (.A(_26347_),
    .Z(_26354_));
 MUX2_X1 _57991_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [927]),
    .B(lce_data_cmd_i[409]),
    .S(_26354_),
    .Z(_06466_));
 MUX2_X1 _57992_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [928]),
    .B(lce_data_cmd_i[410]),
    .S(_26354_),
    .Z(_06467_));
 MUX2_X1 _57993_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [929]),
    .B(lce_data_cmd_i[411]),
    .S(_26354_),
    .Z(_06468_));
 MUX2_X1 _57994_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [930]),
    .B(lce_data_cmd_i[412]),
    .S(_26354_),
    .Z(_06470_));
 MUX2_X1 _57995_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [931]),
    .B(lce_data_cmd_i[413]),
    .S(_26354_),
    .Z(_06471_));
 MUX2_X1 _57996_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [932]),
    .B(lce_data_cmd_i[414]),
    .S(_26354_),
    .Z(_06472_));
 MUX2_X1 _57997_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [933]),
    .B(lce_data_cmd_i[415]),
    .S(_26354_),
    .Z(_06473_));
 MUX2_X1 _57998_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [934]),
    .B(lce_data_cmd_i[416]),
    .S(_26354_),
    .Z(_06474_));
 MUX2_X1 _57999_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [935]),
    .B(lce_data_cmd_i[417]),
    .S(_26354_),
    .Z(_06475_));
 MUX2_X1 _58000_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [936]),
    .B(lce_data_cmd_i[418]),
    .S(_26354_),
    .Z(_06476_));
 BUF_X8 _58001_ (.A(_26347_),
    .Z(_26355_));
 MUX2_X1 _58002_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [520]),
    .B(lce_data_cmd_i[2]),
    .S(_26355_),
    .Z(_06017_));
 MUX2_X1 _58003_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [739]),
    .B(lce_data_cmd_i[221]),
    .S(_26355_),
    .Z(_06257_));
 MUX2_X1 _58004_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [740]),
    .B(lce_data_cmd_i[222]),
    .S(_26355_),
    .Z(_06259_));
 MUX2_X1 _58005_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [741]),
    .B(lce_data_cmd_i[223]),
    .S(_26355_),
    .Z(_06260_));
 MUX2_X1 _58006_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [742]),
    .B(lce_data_cmd_i[224]),
    .S(_26355_),
    .Z(_06261_));
 MUX2_X1 _58007_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [743]),
    .B(lce_data_cmd_i[225]),
    .S(_26355_),
    .Z(_06262_));
 MUX2_X1 _58008_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [744]),
    .B(lce_data_cmd_i[226]),
    .S(_26355_),
    .Z(_06263_));
 MUX2_X1 _58009_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [745]),
    .B(lce_data_cmd_i[227]),
    .S(_26355_),
    .Z(_06264_));
 MUX2_X1 _58010_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [746]),
    .B(lce_data_cmd_i[228]),
    .S(_26355_),
    .Z(_06265_));
 MUX2_X1 _58011_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [747]),
    .B(lce_data_cmd_i[229]),
    .S(_26355_),
    .Z(_06266_));
 BUF_X8 _58012_ (.A(_26347_),
    .Z(_26356_));
 MUX2_X1 _58013_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [748]),
    .B(lce_data_cmd_i[230]),
    .S(_26356_),
    .Z(_06267_));
 MUX2_X1 _58014_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [749]),
    .B(lce_data_cmd_i[231]),
    .S(_26356_),
    .Z(_06268_));
 MUX2_X1 _58015_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [750]),
    .B(lce_data_cmd_i[232]),
    .S(_26356_),
    .Z(_06270_));
 MUX2_X1 _58016_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [751]),
    .B(lce_data_cmd_i[233]),
    .S(_26356_),
    .Z(_06271_));
 MUX2_X1 _58017_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [752]),
    .B(lce_data_cmd_i[234]),
    .S(_26356_),
    .Z(_06272_));
 MUX2_X1 _58018_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [753]),
    .B(lce_data_cmd_i[235]),
    .S(_26356_),
    .Z(_06273_));
 MUX2_X1 _58019_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [754]),
    .B(lce_data_cmd_i[236]),
    .S(_26356_),
    .Z(_06274_));
 MUX2_X1 _58020_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [755]),
    .B(lce_data_cmd_i[237]),
    .S(_26356_),
    .Z(_06275_));
 MUX2_X1 _58021_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [756]),
    .B(lce_data_cmd_i[238]),
    .S(_26356_),
    .Z(_06276_));
 MUX2_X1 _58022_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [757]),
    .B(lce_data_cmd_i[239]),
    .S(_26356_),
    .Z(_06277_));
 BUF_X8 _58023_ (.A(_26347_),
    .Z(_26357_));
 MUX2_X1 _58024_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [758]),
    .B(lce_data_cmd_i[240]),
    .S(_26357_),
    .Z(_06278_));
 MUX2_X1 _58025_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [759]),
    .B(lce_data_cmd_i[241]),
    .S(_26357_),
    .Z(_06279_));
 MUX2_X1 _58026_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [760]),
    .B(lce_data_cmd_i[242]),
    .S(_26357_),
    .Z(_06281_));
 MUX2_X1 _58027_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [761]),
    .B(lce_data_cmd_i[243]),
    .S(_26357_),
    .Z(_06282_));
 MUX2_X1 _58028_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [762]),
    .B(lce_data_cmd_i[244]),
    .S(_26357_),
    .Z(_06283_));
 MUX2_X1 _58029_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [763]),
    .B(lce_data_cmd_i[245]),
    .S(_26357_),
    .Z(_06284_));
 MUX2_X1 _58030_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [764]),
    .B(lce_data_cmd_i[246]),
    .S(_26357_),
    .Z(_06285_));
 MUX2_X1 _58031_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [765]),
    .B(lce_data_cmd_i[247]),
    .S(_26357_),
    .Z(_06286_));
 MUX2_X1 _58032_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [766]),
    .B(lce_data_cmd_i[248]),
    .S(_26357_),
    .Z(_06287_));
 MUX2_X1 _58033_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [767]),
    .B(lce_data_cmd_i[249]),
    .S(_26357_),
    .Z(_06288_));
 BUF_X32 _58034_ (.A(_26319_),
    .Z(_26358_));
 BUF_X8 _58035_ (.A(_26358_),
    .Z(_26359_));
 MUX2_X1 _58036_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [768]),
    .B(lce_data_cmd_i[250]),
    .S(_26359_),
    .Z(_06289_));
 MUX2_X1 _58037_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [769]),
    .B(lce_data_cmd_i[251]),
    .S(_26359_),
    .Z(_06290_));
 MUX2_X1 _58038_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [770]),
    .B(lce_data_cmd_i[252]),
    .S(_26359_),
    .Z(_06292_));
 MUX2_X1 _58039_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [771]),
    .B(lce_data_cmd_i[253]),
    .S(_26359_),
    .Z(_06293_));
 MUX2_X1 _58040_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [772]),
    .B(lce_data_cmd_i[254]),
    .S(_26359_),
    .Z(_06294_));
 MUX2_X1 _58041_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [773]),
    .B(lce_data_cmd_i[255]),
    .S(_26359_),
    .Z(_06295_));
 MUX2_X1 _58042_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [774]),
    .B(lce_data_cmd_i[256]),
    .S(_26359_),
    .Z(_06296_));
 MUX2_X1 _58043_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [775]),
    .B(lce_data_cmd_i[257]),
    .S(_26359_),
    .Z(_06297_));
 MUX2_X1 _58044_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [776]),
    .B(lce_data_cmd_i[258]),
    .S(_26359_),
    .Z(_06298_));
 MUX2_X1 _58045_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [777]),
    .B(lce_data_cmd_i[259]),
    .S(_26359_),
    .Z(_06299_));
 BUF_X16 _58046_ (.A(_26358_),
    .Z(_26360_));
 MUX2_X1 _58047_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [778]),
    .B(lce_data_cmd_i[260]),
    .S(_26360_),
    .Z(_06300_));
 MUX2_X1 _58048_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [779]),
    .B(lce_data_cmd_i[261]),
    .S(_26360_),
    .Z(_06301_));
 MUX2_X1 _58049_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [780]),
    .B(lce_data_cmd_i[262]),
    .S(_26360_),
    .Z(_06303_));
 MUX2_X1 _58050_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [781]),
    .B(lce_data_cmd_i[263]),
    .S(_26360_),
    .Z(_06304_));
 MUX2_X1 _58051_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [782]),
    .B(lce_data_cmd_i[264]),
    .S(_26360_),
    .Z(_06305_));
 MUX2_X1 _58052_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [783]),
    .B(lce_data_cmd_i[265]),
    .S(_26360_),
    .Z(_06306_));
 MUX2_X1 _58053_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [784]),
    .B(lce_data_cmd_i[266]),
    .S(_26360_),
    .Z(_06307_));
 MUX2_X1 _58054_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [785]),
    .B(lce_data_cmd_i[267]),
    .S(_26360_),
    .Z(_06308_));
 MUX2_X1 _58055_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [786]),
    .B(lce_data_cmd_i[268]),
    .S(_26360_),
    .Z(_06309_));
 MUX2_X1 _58056_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [787]),
    .B(lce_data_cmd_i[269]),
    .S(_26360_),
    .Z(_06310_));
 BUF_X8 _58057_ (.A(_26358_),
    .Z(_26361_));
 MUX2_X1 _58058_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [788]),
    .B(lce_data_cmd_i[270]),
    .S(_26361_),
    .Z(_06311_));
 MUX2_X1 _58059_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [789]),
    .B(lce_data_cmd_i[271]),
    .S(_26361_),
    .Z(_06312_));
 MUX2_X1 _58060_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [790]),
    .B(lce_data_cmd_i[272]),
    .S(_26361_),
    .Z(_06314_));
 MUX2_X1 _58061_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [791]),
    .B(lce_data_cmd_i[273]),
    .S(_26361_),
    .Z(_06315_));
 MUX2_X1 _58062_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [792]),
    .B(lce_data_cmd_i[274]),
    .S(_26361_),
    .Z(_06316_));
 MUX2_X1 _58063_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [793]),
    .B(lce_data_cmd_i[275]),
    .S(_26361_),
    .Z(_06317_));
 MUX2_X1 _58064_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [794]),
    .B(lce_data_cmd_i[276]),
    .S(_26361_),
    .Z(_06318_));
 MUX2_X1 _58065_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [795]),
    .B(lce_data_cmd_i[277]),
    .S(_26361_),
    .Z(_06319_));
 MUX2_X1 _58066_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [796]),
    .B(lce_data_cmd_i[278]),
    .S(_26361_),
    .Z(_06320_));
 MUX2_X1 _58067_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [797]),
    .B(lce_data_cmd_i[279]),
    .S(_26361_),
    .Z(_06321_));
 BUF_X8 _58068_ (.A(_26358_),
    .Z(_26362_));
 MUX2_X1 _58069_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [798]),
    .B(lce_data_cmd_i[280]),
    .S(_26362_),
    .Z(_06322_));
 MUX2_X1 _58070_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [799]),
    .B(lce_data_cmd_i[281]),
    .S(_26362_),
    .Z(_06323_));
 MUX2_X1 _58071_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [800]),
    .B(lce_data_cmd_i[282]),
    .S(_26362_),
    .Z(_06326_));
 MUX2_X1 _58072_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [801]),
    .B(lce_data_cmd_i[283]),
    .S(_26362_),
    .Z(_06327_));
 MUX2_X1 _58073_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [802]),
    .B(lce_data_cmd_i[284]),
    .S(_26362_),
    .Z(_06328_));
 MUX2_X1 _58074_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [803]),
    .B(lce_data_cmd_i[285]),
    .S(_26362_),
    .Z(_06329_));
 MUX2_X1 _58075_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [804]),
    .B(lce_data_cmd_i[286]),
    .S(_26362_),
    .Z(_06330_));
 MUX2_X1 _58076_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [805]),
    .B(lce_data_cmd_i[287]),
    .S(_26362_),
    .Z(_06331_));
 MUX2_X1 _58077_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [806]),
    .B(lce_data_cmd_i[288]),
    .S(_26362_),
    .Z(_06332_));
 MUX2_X1 _58078_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [807]),
    .B(lce_data_cmd_i[289]),
    .S(_26362_),
    .Z(_06333_));
 BUF_X8 _58079_ (.A(_26358_),
    .Z(_26363_));
 MUX2_X1 _58080_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [808]),
    .B(lce_data_cmd_i[290]),
    .S(_26363_),
    .Z(_06334_));
 MUX2_X1 _58081_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [809]),
    .B(lce_data_cmd_i[291]),
    .S(_26363_),
    .Z(_06335_));
 MUX2_X1 _58082_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [810]),
    .B(lce_data_cmd_i[292]),
    .S(_26363_),
    .Z(_06337_));
 MUX2_X1 _58083_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [811]),
    .B(lce_data_cmd_i[293]),
    .S(_26363_),
    .Z(_06338_));
 MUX2_X1 _58084_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [812]),
    .B(lce_data_cmd_i[294]),
    .S(_26363_),
    .Z(_06339_));
 MUX2_X1 _58085_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [813]),
    .B(lce_data_cmd_i[295]),
    .S(_26363_),
    .Z(_06340_));
 MUX2_X1 _58086_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [814]),
    .B(lce_data_cmd_i[296]),
    .S(_26363_),
    .Z(_06341_));
 MUX2_X1 _58087_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [815]),
    .B(lce_data_cmd_i[297]),
    .S(_26363_),
    .Z(_06342_));
 MUX2_X1 _58088_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [816]),
    .B(lce_data_cmd_i[298]),
    .S(_26363_),
    .Z(_06343_));
 MUX2_X1 _58089_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [817]),
    .B(lce_data_cmd_i[299]),
    .S(_26363_),
    .Z(_06344_));
 BUF_X4 _58090_ (.A(_26358_),
    .Z(_26364_));
 MUX2_X1 _58091_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [818]),
    .B(lce_data_cmd_i[300]),
    .S(_26364_),
    .Z(_06345_));
 MUX2_X1 _58092_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [819]),
    .B(lce_data_cmd_i[301]),
    .S(_26364_),
    .Z(_06346_));
 MUX2_X1 _58093_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [820]),
    .B(lce_data_cmd_i[302]),
    .S(_26364_),
    .Z(_06348_));
 MUX2_X1 _58094_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [821]),
    .B(lce_data_cmd_i[303]),
    .S(_26364_),
    .Z(_06349_));
 MUX2_X1 _58095_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [822]),
    .B(lce_data_cmd_i[304]),
    .S(_26364_),
    .Z(_06350_));
 MUX2_X1 _58096_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [823]),
    .B(lce_data_cmd_i[305]),
    .S(_26364_),
    .Z(_06351_));
 MUX2_X1 _58097_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [824]),
    .B(lce_data_cmd_i[306]),
    .S(_26364_),
    .Z(_06352_));
 MUX2_X1 _58098_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [825]),
    .B(lce_data_cmd_i[307]),
    .S(_26364_),
    .Z(_06353_));
 MUX2_X1 _58099_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [826]),
    .B(lce_data_cmd_i[308]),
    .S(_26364_),
    .Z(_06354_));
 MUX2_X1 _58100_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [827]),
    .B(lce_data_cmd_i[309]),
    .S(_26364_),
    .Z(_06355_));
 BUF_X16 _58101_ (.A(_26358_),
    .Z(_26365_));
 MUX2_X1 _58102_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [828]),
    .B(lce_data_cmd_i[310]),
    .S(_26365_),
    .Z(_06356_));
 MUX2_X1 _58103_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [829]),
    .B(lce_data_cmd_i[311]),
    .S(_26365_),
    .Z(_06357_));
 MUX2_X1 _58104_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [830]),
    .B(lce_data_cmd_i[312]),
    .S(_26365_),
    .Z(_06359_));
 MUX2_X1 _58105_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [831]),
    .B(lce_data_cmd_i[313]),
    .S(_26365_),
    .Z(_06360_));
 MUX2_X1 _58106_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [832]),
    .B(lce_data_cmd_i[314]),
    .S(_26365_),
    .Z(_06361_));
 MUX2_X1 _58107_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [833]),
    .B(lce_data_cmd_i[315]),
    .S(_26365_),
    .Z(_06362_));
 MUX2_X1 _58108_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [834]),
    .B(lce_data_cmd_i[316]),
    .S(_26365_),
    .Z(_06363_));
 MUX2_X1 _58109_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [835]),
    .B(lce_data_cmd_i[317]),
    .S(_26365_),
    .Z(_06364_));
 MUX2_X1 _58110_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [836]),
    .B(lce_data_cmd_i[318]),
    .S(_26365_),
    .Z(_06365_));
 MUX2_X1 _58111_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [837]),
    .B(lce_data_cmd_i[319]),
    .S(_26365_),
    .Z(_06366_));
 BUF_X8 _58112_ (.A(_26358_),
    .Z(_26366_));
 MUX2_X1 _58113_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [640]),
    .B(lce_data_cmd_i[122]),
    .S(_26366_),
    .Z(_06148_));
 MUX2_X1 _58114_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [641]),
    .B(lce_data_cmd_i[123]),
    .S(_26366_),
    .Z(_06149_));
 MUX2_X1 _58115_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [642]),
    .B(lce_data_cmd_i[124]),
    .S(_26366_),
    .Z(_06150_));
 MUX2_X1 _58116_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [643]),
    .B(lce_data_cmd_i[125]),
    .S(_26366_),
    .Z(_06151_));
 MUX2_X1 _58117_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [644]),
    .B(lce_data_cmd_i[126]),
    .S(_26366_),
    .Z(_06152_));
 MUX2_X1 _58118_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [645]),
    .B(lce_data_cmd_i[127]),
    .S(_26366_),
    .Z(_06153_));
 MUX2_X1 _58119_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [646]),
    .B(lce_data_cmd_i[128]),
    .S(_26366_),
    .Z(_06154_));
 MUX2_X1 _58120_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [647]),
    .B(lce_data_cmd_i[129]),
    .S(_26366_),
    .Z(_06155_));
 MUX2_X1 _58121_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [648]),
    .B(lce_data_cmd_i[130]),
    .S(_26366_),
    .Z(_06156_));
 MUX2_X1 _58122_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [649]),
    .B(lce_data_cmd_i[131]),
    .S(_26366_),
    .Z(_06157_));
 BUF_X8 _58123_ (.A(_26358_),
    .Z(_26367_));
 MUX2_X1 _58124_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [650]),
    .B(lce_data_cmd_i[132]),
    .S(_26367_),
    .Z(_06159_));
 MUX2_X1 _58125_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [651]),
    .B(lce_data_cmd_i[133]),
    .S(_26367_),
    .Z(_06160_));
 MUX2_X1 _58126_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [652]),
    .B(lce_data_cmd_i[134]),
    .S(_26367_),
    .Z(_06161_));
 MUX2_X1 _58127_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [653]),
    .B(lce_data_cmd_i[135]),
    .S(_26367_),
    .Z(_06162_));
 MUX2_X1 _58128_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [654]),
    .B(lce_data_cmd_i[136]),
    .S(_26367_),
    .Z(_06163_));
 MUX2_X1 _58129_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [655]),
    .B(lce_data_cmd_i[137]),
    .S(_26367_),
    .Z(_06164_));
 MUX2_X1 _58130_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [656]),
    .B(lce_data_cmd_i[138]),
    .S(_26367_),
    .Z(_06165_));
 MUX2_X1 _58131_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [657]),
    .B(lce_data_cmd_i[139]),
    .S(_26367_),
    .Z(_06166_));
 MUX2_X1 _58132_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [658]),
    .B(lce_data_cmd_i[140]),
    .S(_26367_),
    .Z(_06167_));
 MUX2_X1 _58133_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [659]),
    .B(lce_data_cmd_i[141]),
    .S(_26367_),
    .Z(_06168_));
 BUF_X8 _58134_ (.A(_26358_),
    .Z(_26368_));
 MUX2_X1 _58135_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [660]),
    .B(lce_data_cmd_i[142]),
    .S(_26368_),
    .Z(_06170_));
 MUX2_X1 _58136_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [661]),
    .B(lce_data_cmd_i[143]),
    .S(_26368_),
    .Z(_06171_));
 MUX2_X1 _58137_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [662]),
    .B(lce_data_cmd_i[144]),
    .S(_26368_),
    .Z(_06172_));
 MUX2_X1 _58138_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [663]),
    .B(lce_data_cmd_i[145]),
    .S(_26368_),
    .Z(_06173_));
 MUX2_X1 _58139_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [664]),
    .B(lce_data_cmd_i[146]),
    .S(_26368_),
    .Z(_06174_));
 MUX2_X1 _58140_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [665]),
    .B(lce_data_cmd_i[147]),
    .S(_26368_),
    .Z(_06175_));
 MUX2_X1 _58141_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [666]),
    .B(lce_data_cmd_i[148]),
    .S(_26368_),
    .Z(_06176_));
 MUX2_X1 _58142_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [667]),
    .B(lce_data_cmd_i[149]),
    .S(_26368_),
    .Z(_06177_));
 MUX2_X1 _58143_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [668]),
    .B(lce_data_cmd_i[150]),
    .S(_26368_),
    .Z(_06178_));
 MUX2_X1 _58144_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [669]),
    .B(lce_data_cmd_i[151]),
    .S(_26368_),
    .Z(_06179_));
 BUF_X8 _58145_ (.A(_26324_),
    .Z(_26369_));
 MUX2_X1 _58146_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [670]),
    .B(lce_data_cmd_i[152]),
    .S(_26369_),
    .Z(_06181_));
 MUX2_X1 _58147_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [671]),
    .B(lce_data_cmd_i[153]),
    .S(_26369_),
    .Z(_06182_));
 MUX2_X1 _58148_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [672]),
    .B(lce_data_cmd_i[154]),
    .S(_26369_),
    .Z(_06183_));
 MUX2_X1 _58149_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [673]),
    .B(lce_data_cmd_i[155]),
    .S(_26369_),
    .Z(_06184_));
 MUX2_X1 _58150_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [674]),
    .B(lce_data_cmd_i[156]),
    .S(_26369_),
    .Z(_06185_));
 MUX2_X1 _58151_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [675]),
    .B(lce_data_cmd_i[157]),
    .S(_26369_),
    .Z(_06186_));
 MUX2_X1 _58152_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [676]),
    .B(lce_data_cmd_i[158]),
    .S(_26369_),
    .Z(_06187_));
 MUX2_X1 _58153_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [677]),
    .B(lce_data_cmd_i[159]),
    .S(_26369_),
    .Z(_06188_));
 MUX2_X1 _58154_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [678]),
    .B(lce_data_cmd_i[160]),
    .S(_26369_),
    .Z(_06189_));
 MUX2_X1 _58155_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [679]),
    .B(lce_data_cmd_i[161]),
    .S(_26369_),
    .Z(_06190_));
 BUF_X8 _58156_ (.A(_26324_),
    .Z(_26370_));
 MUX2_X1 _58157_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [680]),
    .B(lce_data_cmd_i[162]),
    .S(_26370_),
    .Z(_06192_));
 MUX2_X1 _58158_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [681]),
    .B(lce_data_cmd_i[163]),
    .S(_26370_),
    .Z(_06193_));
 MUX2_X1 _58159_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [682]),
    .B(lce_data_cmd_i[164]),
    .S(_26370_),
    .Z(_06194_));
 MUX2_X1 _58160_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [683]),
    .B(lce_data_cmd_i[165]),
    .S(_26370_),
    .Z(_06195_));
 MUX2_X1 _58161_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [684]),
    .B(lce_data_cmd_i[166]),
    .S(_26370_),
    .Z(_06196_));
 MUX2_X1 _58162_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [685]),
    .B(lce_data_cmd_i[167]),
    .S(_26370_),
    .Z(_06197_));
 MUX2_X1 _58163_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [686]),
    .B(lce_data_cmd_i[168]),
    .S(_26370_),
    .Z(_06198_));
 MUX2_X1 _58164_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [687]),
    .B(lce_data_cmd_i[169]),
    .S(_26370_),
    .Z(_06199_));
 MUX2_X1 _58165_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [688]),
    .B(lce_data_cmd_i[170]),
    .S(_26370_),
    .Z(_06200_));
 MUX2_X1 _58166_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [689]),
    .B(lce_data_cmd_i[171]),
    .S(_26370_),
    .Z(_06201_));
 BUF_X8 _58167_ (.A(_26324_),
    .Z(_26371_));
 MUX2_X1 _58168_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [690]),
    .B(lce_data_cmd_i[172]),
    .S(_26371_),
    .Z(_06203_));
 MUX2_X1 _58169_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [691]),
    .B(lce_data_cmd_i[173]),
    .S(_26371_),
    .Z(_06204_));
 MUX2_X1 _58170_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [692]),
    .B(lce_data_cmd_i[174]),
    .S(_26371_),
    .Z(_06205_));
 MUX2_X1 _58171_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [693]),
    .B(lce_data_cmd_i[175]),
    .S(_26371_),
    .Z(_06206_));
 MUX2_X1 _58172_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [694]),
    .B(lce_data_cmd_i[176]),
    .S(_26371_),
    .Z(_06207_));
 MUX2_X1 _58173_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [695]),
    .B(lce_data_cmd_i[177]),
    .S(_26371_),
    .Z(_06208_));
 MUX2_X1 _58174_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [696]),
    .B(lce_data_cmd_i[178]),
    .S(_26371_),
    .Z(_06209_));
 MUX2_X1 _58175_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [697]),
    .B(lce_data_cmd_i[179]),
    .S(_26371_),
    .Z(_06210_));
 MUX2_X1 _58176_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [698]),
    .B(lce_data_cmd_i[180]),
    .S(_26371_),
    .Z(_06211_));
 MUX2_X1 _58177_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [699]),
    .B(lce_data_cmd_i[181]),
    .S(_26371_),
    .Z(_06212_));
 BUF_X8 _58178_ (.A(_26324_),
    .Z(_26372_));
 MUX2_X1 _58179_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [700]),
    .B(lce_data_cmd_i[182]),
    .S(_26372_),
    .Z(_06215_));
 MUX2_X1 _58180_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [701]),
    .B(lce_data_cmd_i[183]),
    .S(_26372_),
    .Z(_06216_));
 MUX2_X1 _58181_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [702]),
    .B(lce_data_cmd_i[184]),
    .S(_26372_),
    .Z(_06217_));
 MUX2_X1 _58182_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [703]),
    .B(lce_data_cmd_i[185]),
    .S(_26372_),
    .Z(_06218_));
 MUX2_X1 _58183_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [704]),
    .B(lce_data_cmd_i[186]),
    .S(_26372_),
    .Z(_06219_));
 MUX2_X1 _58184_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [705]),
    .B(lce_data_cmd_i[187]),
    .S(_26372_),
    .Z(_06220_));
 MUX2_X1 _58185_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [706]),
    .B(lce_data_cmd_i[188]),
    .S(_26372_),
    .Z(_06221_));
 MUX2_X1 _58186_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [707]),
    .B(lce_data_cmd_i[189]),
    .S(_26372_),
    .Z(_06222_));
 MUX2_X1 _58187_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [708]),
    .B(lce_data_cmd_i[190]),
    .S(_26372_),
    .Z(_06223_));
 MUX2_X1 _58188_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [709]),
    .B(lce_data_cmd_i[191]),
    .S(_26372_),
    .Z(_06224_));
 BUF_X16 _58189_ (.A(_26324_),
    .Z(_26373_));
 MUX2_X1 _58190_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [710]),
    .B(lce_data_cmd_i[192]),
    .S(_26373_),
    .Z(_06226_));
 MUX2_X1 _58191_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [711]),
    .B(lce_data_cmd_i[193]),
    .S(_26373_),
    .Z(_06227_));
 MUX2_X1 _58192_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [712]),
    .B(lce_data_cmd_i[194]),
    .S(_26373_),
    .Z(_06228_));
 MUX2_X1 _58193_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [713]),
    .B(lce_data_cmd_i[195]),
    .S(_26373_),
    .Z(_06229_));
 MUX2_X1 _58194_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [714]),
    .B(lce_data_cmd_i[196]),
    .S(_26373_),
    .Z(_06230_));
 MUX2_X1 _58195_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [715]),
    .B(lce_data_cmd_i[197]),
    .S(_26373_),
    .Z(_06231_));
 MUX2_X1 _58196_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [716]),
    .B(lce_data_cmd_i[198]),
    .S(_26373_),
    .Z(_06232_));
 MUX2_X1 _58197_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [717]),
    .B(lce_data_cmd_i[199]),
    .S(_26373_),
    .Z(_06233_));
 MUX2_X1 _58198_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [718]),
    .B(lce_data_cmd_i[200]),
    .S(_26373_),
    .Z(_06234_));
 MUX2_X1 _58199_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [719]),
    .B(lce_data_cmd_i[201]),
    .S(_26373_),
    .Z(_06235_));
 BUF_X16 _58200_ (.A(_26324_),
    .Z(_26374_));
 MUX2_X1 _58201_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [720]),
    .B(lce_data_cmd_i[202]),
    .S(_26374_),
    .Z(_06237_));
 MUX2_X1 _58202_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [721]),
    .B(lce_data_cmd_i[203]),
    .S(_26374_),
    .Z(_06238_));
 MUX2_X1 _58203_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [722]),
    .B(lce_data_cmd_i[204]),
    .S(_26374_),
    .Z(_06239_));
 MUX2_X1 _58204_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [723]),
    .B(lce_data_cmd_i[205]),
    .S(_26374_),
    .Z(_06240_));
 MUX2_X1 _58205_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [724]),
    .B(lce_data_cmd_i[206]),
    .S(_26374_),
    .Z(_06241_));
 MUX2_X1 _58206_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [725]),
    .B(lce_data_cmd_i[207]),
    .S(_26374_),
    .Z(_06242_));
 MUX2_X1 _58207_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [726]),
    .B(lce_data_cmd_i[208]),
    .S(_26374_),
    .Z(_06243_));
 MUX2_X1 _58208_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [727]),
    .B(lce_data_cmd_i[209]),
    .S(_26374_),
    .Z(_06244_));
 MUX2_X1 _58209_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [728]),
    .B(lce_data_cmd_i[210]),
    .S(_26374_),
    .Z(_06245_));
 MUX2_X1 _58210_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [729]),
    .B(lce_data_cmd_i[211]),
    .S(_26374_),
    .Z(_06246_));
 BUF_X16 _58211_ (.A(_26324_),
    .Z(_26375_));
 MUX2_X1 _58212_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [730]),
    .B(lce_data_cmd_i[212]),
    .S(_26375_),
    .Z(_06248_));
 MUX2_X1 _58213_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [731]),
    .B(lce_data_cmd_i[213]),
    .S(_26375_),
    .Z(_06249_));
 MUX2_X1 _58214_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [732]),
    .B(lce_data_cmd_i[214]),
    .S(_26375_),
    .Z(_06250_));
 MUX2_X1 _58215_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [733]),
    .B(lce_data_cmd_i[215]),
    .S(_26375_),
    .Z(_06251_));
 MUX2_X1 _58216_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [734]),
    .B(lce_data_cmd_i[216]),
    .S(_26375_),
    .Z(_06252_));
 MUX2_X1 _58217_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [735]),
    .B(lce_data_cmd_i[217]),
    .S(_26375_),
    .Z(_06253_));
 MUX2_X1 _58218_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [736]),
    .B(lce_data_cmd_i[218]),
    .S(_26375_),
    .Z(_06254_));
 MUX2_X1 _58219_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [737]),
    .B(lce_data_cmd_i[219]),
    .S(_26375_),
    .Z(_06255_));
 MUX2_X1 _58220_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [738]),
    .B(lce_data_cmd_i[220]),
    .S(_26375_),
    .Z(_06256_));
 MUX2_X1 _58221_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [522]),
    .B(lce_data_cmd_i[4]),
    .S(_26375_),
    .Z(_06019_));
 BUF_X16 _58222_ (.A(_26324_),
    .Z(_26376_));
 MUX2_X1 _58223_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [524]),
    .B(lce_data_cmd_i[6]),
    .S(_26376_),
    .Z(_06020_));
 MUX2_X1 _58224_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [525]),
    .B(lce_data_cmd_i[7]),
    .S(_26376_),
    .Z(_06021_));
 MUX2_X1 _58225_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [526]),
    .B(lce_data_cmd_i[8]),
    .S(_26376_),
    .Z(_06022_));
 MUX2_X1 _58226_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [527]),
    .B(lce_data_cmd_i[9]),
    .S(_26376_),
    .Z(_06023_));
 MUX2_X1 _58227_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [528]),
    .B(lce_data_cmd_i[10]),
    .S(_26376_),
    .Z(_06024_));
 MUX2_X1 _58228_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [529]),
    .B(lce_data_cmd_i[11]),
    .S(_26376_),
    .Z(_06025_));
 MUX2_X1 _58229_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [530]),
    .B(lce_data_cmd_i[12]),
    .S(_26376_),
    .Z(_06027_));
 MUX2_X1 _58230_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [531]),
    .B(lce_data_cmd_i[13]),
    .S(_26376_),
    .Z(_06028_));
 MUX2_X1 _58231_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [532]),
    .B(lce_data_cmd_i[14]),
    .S(_26376_),
    .Z(_06029_));
 MUX2_X1 _58232_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [533]),
    .B(lce_data_cmd_i[15]),
    .S(_26376_),
    .Z(_06030_));
 MUX2_X1 _58233_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [534]),
    .B(lce_data_cmd_i[16]),
    .S(_26320_),
    .Z(_06031_));
 MUX2_X1 _58234_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [535]),
    .B(lce_data_cmd_i[17]),
    .S(_26320_),
    .Z(_06032_));
 MUX2_X1 _58235_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [536]),
    .B(lce_data_cmd_i[18]),
    .S(_26320_),
    .Z(_06033_));
 MUX2_X1 _58236_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [537]),
    .B(lce_data_cmd_i[19]),
    .S(_26320_),
    .Z(_06034_));
 MUX2_X1 _58237_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [538]),
    .B(lce_data_cmd_i[20]),
    .S(_26320_),
    .Z(_06035_));
 MUX2_X1 _58238_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [539]),
    .B(lce_data_cmd_i[21]),
    .S(_26320_),
    .Z(_06036_));
 MUX2_X1 _58239_ (.A(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [540]),
    .B(lce_data_cmd_i[22]),
    .S(_26320_),
    .Z(_06038_));
 NAND2_X4 _58240_ (.A1(_21282_),
    .A2(_21283_),
    .ZN(_26377_));
 BUF_X16 _58241_ (.A(_26377_),
    .Z(_26378_));
 BUF_X8 _58242_ (.A(_26378_),
    .Z(_26379_));
 MUX2_X1 _58243_ (.A(lce_data_cmd_i[0]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [0]),
    .S(_26379_),
    .Z(_05514_));
 MUX2_X1 _58244_ (.A(lce_data_cmd_i[419]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [419]),
    .S(_26379_),
    .Z(_05904_));
 MUX2_X1 _58245_ (.A(lce_data_cmd_i[420]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [420]),
    .S(_26379_),
    .Z(_05906_));
 MUX2_X1 _58246_ (.A(lce_data_cmd_i[421]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [421]),
    .S(_26379_),
    .Z(_05907_));
 MUX2_X1 _58247_ (.A(lce_data_cmd_i[422]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [422]),
    .S(_26379_),
    .Z(_05908_));
 MUX2_X1 _58248_ (.A(lce_data_cmd_i[423]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [423]),
    .S(_26379_),
    .Z(_05909_));
 MUX2_X1 _58249_ (.A(lce_data_cmd_i[424]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [424]),
    .S(_26379_),
    .Z(_05910_));
 MUX2_X1 _58250_ (.A(lce_data_cmd_i[425]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [425]),
    .S(_26379_),
    .Z(_05911_));
 MUX2_X1 _58251_ (.A(lce_data_cmd_i[426]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [426]),
    .S(_26379_),
    .Z(_05912_));
 MUX2_X1 _58252_ (.A(lce_data_cmd_i[427]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [427]),
    .S(_26379_),
    .Z(_05913_));
 BUF_X8 _58253_ (.A(_26378_),
    .Z(_26380_));
 MUX2_X1 _58254_ (.A(lce_data_cmd_i[428]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [428]),
    .S(_26380_),
    .Z(_05914_));
 MUX2_X1 _58255_ (.A(lce_data_cmd_i[429]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [429]),
    .S(_26380_),
    .Z(_05915_));
 MUX2_X1 _58256_ (.A(lce_data_cmd_i[430]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [430]),
    .S(_26380_),
    .Z(_05917_));
 MUX2_X1 _58257_ (.A(lce_data_cmd_i[431]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [431]),
    .S(_26380_),
    .Z(_05918_));
 MUX2_X1 _58258_ (.A(lce_data_cmd_i[432]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [432]),
    .S(_26380_),
    .Z(_05919_));
 MUX2_X1 _58259_ (.A(lce_data_cmd_i[433]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [433]),
    .S(_26380_),
    .Z(_05920_));
 MUX2_X1 _58260_ (.A(lce_data_cmd_i[434]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [434]),
    .S(_26380_),
    .Z(_05921_));
 MUX2_X1 _58261_ (.A(lce_data_cmd_i[435]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [435]),
    .S(_26380_),
    .Z(_05922_));
 MUX2_X1 _58262_ (.A(lce_data_cmd_i[436]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [436]),
    .S(_26380_),
    .Z(_05923_));
 MUX2_X1 _58263_ (.A(lce_data_cmd_i[437]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [437]),
    .S(_26380_),
    .Z(_05924_));
 BUF_X8 _58264_ (.A(_26378_),
    .Z(_26381_));
 MUX2_X1 _58265_ (.A(lce_data_cmd_i[438]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [438]),
    .S(_26381_),
    .Z(_05925_));
 MUX2_X1 _58266_ (.A(lce_data_cmd_i[439]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [439]),
    .S(_26381_),
    .Z(_05926_));
 MUX2_X1 _58267_ (.A(lce_data_cmd_i[440]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [440]),
    .S(_26381_),
    .Z(_05928_));
 MUX2_X1 _58268_ (.A(lce_data_cmd_i[441]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [441]),
    .S(_26381_),
    .Z(_05929_));
 MUX2_X1 _58269_ (.A(lce_data_cmd_i[442]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [442]),
    .S(_26381_),
    .Z(_05930_));
 MUX2_X1 _58270_ (.A(lce_data_cmd_i[443]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [443]),
    .S(_26381_),
    .Z(_05931_));
 MUX2_X1 _58271_ (.A(lce_data_cmd_i[444]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [444]),
    .S(_26381_),
    .Z(_05932_));
 MUX2_X1 _58272_ (.A(lce_data_cmd_i[445]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [445]),
    .S(_26381_),
    .Z(_05933_));
 MUX2_X1 _58273_ (.A(lce_data_cmd_i[446]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [446]),
    .S(_26381_),
    .Z(_05934_));
 MUX2_X1 _58274_ (.A(lce_data_cmd_i[447]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [447]),
    .S(_26381_),
    .Z(_05935_));
 BUF_X32 _58275_ (.A(_26377_),
    .Z(_26382_));
 BUF_X32 _58276_ (.A(_26382_),
    .Z(_26383_));
 BUF_X8 _58277_ (.A(_26383_),
    .Z(_26384_));
 MUX2_X1 _58278_ (.A(lce_data_cmd_i[448]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [448]),
    .S(_26384_),
    .Z(_05936_));
 MUX2_X1 _58279_ (.A(lce_data_cmd_i[449]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [449]),
    .S(_26384_),
    .Z(_05937_));
 MUX2_X1 _58280_ (.A(lce_data_cmd_i[450]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [450]),
    .S(_26384_),
    .Z(_05939_));
 MUX2_X1 _58281_ (.A(lce_data_cmd_i[451]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [451]),
    .S(_26384_),
    .Z(_05940_));
 MUX2_X1 _58282_ (.A(lce_data_cmd_i[452]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [452]),
    .S(_26384_),
    .Z(_05941_));
 MUX2_X1 _58283_ (.A(lce_data_cmd_i[453]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [453]),
    .S(_26384_),
    .Z(_05942_));
 MUX2_X1 _58284_ (.A(lce_data_cmd_i[454]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [454]),
    .S(_26384_),
    .Z(_05943_));
 MUX2_X1 _58285_ (.A(lce_data_cmd_i[455]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [455]),
    .S(_26384_),
    .Z(_05944_));
 MUX2_X1 _58286_ (.A(lce_data_cmd_i[456]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [456]),
    .S(_26384_),
    .Z(_05945_));
 MUX2_X1 _58287_ (.A(lce_data_cmd_i[457]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [457]),
    .S(_26384_),
    .Z(_05946_));
 BUF_X8 _58288_ (.A(_26383_),
    .Z(_26385_));
 MUX2_X1 _58289_ (.A(lce_data_cmd_i[458]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [458]),
    .S(_26385_),
    .Z(_05947_));
 MUX2_X1 _58290_ (.A(lce_data_cmd_i[459]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [459]),
    .S(_26385_),
    .Z(_05948_));
 MUX2_X1 _58291_ (.A(lce_data_cmd_i[460]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [460]),
    .S(_26385_),
    .Z(_05950_));
 MUX2_X1 _58292_ (.A(lce_data_cmd_i[461]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [461]),
    .S(_26385_),
    .Z(_05951_));
 MUX2_X1 _58293_ (.A(lce_data_cmd_i[462]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [462]),
    .S(_26385_),
    .Z(_05952_));
 MUX2_X1 _58294_ (.A(lce_data_cmd_i[463]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [463]),
    .S(_26385_),
    .Z(_05953_));
 MUX2_X1 _58295_ (.A(lce_data_cmd_i[464]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [464]),
    .S(_26385_),
    .Z(_05954_));
 MUX2_X1 _58296_ (.A(lce_data_cmd_i[465]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [465]),
    .S(_26385_),
    .Z(_05955_));
 MUX2_X1 _58297_ (.A(lce_data_cmd_i[466]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [466]),
    .S(_26385_),
    .Z(_05956_));
 MUX2_X1 _58298_ (.A(lce_data_cmd_i[467]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [467]),
    .S(_26385_),
    .Z(_05957_));
 BUF_X4 _58299_ (.A(_26383_),
    .Z(_26386_));
 MUX2_X1 _58300_ (.A(lce_data_cmd_i[468]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [468]),
    .S(_26386_),
    .Z(_05958_));
 MUX2_X1 _58301_ (.A(lce_data_cmd_i[469]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [469]),
    .S(_26386_),
    .Z(_05959_));
 MUX2_X1 _58302_ (.A(lce_data_cmd_i[470]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [470]),
    .S(_26386_),
    .Z(_05961_));
 MUX2_X1 _58303_ (.A(lce_data_cmd_i[471]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [471]),
    .S(_26386_),
    .Z(_05962_));
 MUX2_X1 _58304_ (.A(lce_data_cmd_i[472]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [472]),
    .S(_26386_),
    .Z(_05963_));
 MUX2_X1 _58305_ (.A(lce_data_cmd_i[473]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [473]),
    .S(_26386_),
    .Z(_05964_));
 MUX2_X1 _58306_ (.A(lce_data_cmd_i[474]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [474]),
    .S(_26386_),
    .Z(_05965_));
 MUX2_X1 _58307_ (.A(lce_data_cmd_i[475]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [475]),
    .S(_26386_),
    .Z(_05966_));
 MUX2_X1 _58308_ (.A(lce_data_cmd_i[476]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [476]),
    .S(_26386_),
    .Z(_05967_));
 MUX2_X1 _58309_ (.A(lce_data_cmd_i[477]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [477]),
    .S(_26386_),
    .Z(_05968_));
 BUF_X8 _58310_ (.A(_26383_),
    .Z(_26387_));
 MUX2_X1 _58311_ (.A(lce_data_cmd_i[478]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [478]),
    .S(_26387_),
    .Z(_05969_));
 MUX2_X1 _58312_ (.A(lce_data_cmd_i[479]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [479]),
    .S(_26387_),
    .Z(_05970_));
 MUX2_X1 _58313_ (.A(lce_data_cmd_i[480]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [480]),
    .S(_26387_),
    .Z(_05972_));
 MUX2_X1 _58314_ (.A(lce_data_cmd_i[481]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [481]),
    .S(_26387_),
    .Z(_05973_));
 MUX2_X1 _58315_ (.A(lce_data_cmd_i[482]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [482]),
    .S(_26387_),
    .Z(_05974_));
 MUX2_X1 _58316_ (.A(lce_data_cmd_i[483]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [483]),
    .S(_26387_),
    .Z(_05975_));
 MUX2_X1 _58317_ (.A(lce_data_cmd_i[484]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [484]),
    .S(_26387_),
    .Z(_05976_));
 MUX2_X1 _58318_ (.A(lce_data_cmd_i[485]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [485]),
    .S(_26387_),
    .Z(_05977_));
 MUX2_X1 _58319_ (.A(lce_data_cmd_i[486]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [486]),
    .S(_26387_),
    .Z(_05978_));
 MUX2_X1 _58320_ (.A(lce_data_cmd_i[487]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [487]),
    .S(_26387_),
    .Z(_05979_));
 BUF_X8 _58321_ (.A(_26383_),
    .Z(_26388_));
 MUX2_X1 _58322_ (.A(lce_data_cmd_i[488]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [488]),
    .S(_26388_),
    .Z(_05980_));
 MUX2_X1 _58323_ (.A(lce_data_cmd_i[489]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [489]),
    .S(_26388_),
    .Z(_05981_));
 MUX2_X1 _58324_ (.A(lce_data_cmd_i[490]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [490]),
    .S(_26388_),
    .Z(_05983_));
 MUX2_X1 _58325_ (.A(lce_data_cmd_i[491]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [491]),
    .S(_26388_),
    .Z(_05984_));
 MUX2_X1 _58326_ (.A(lce_data_cmd_i[492]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [492]),
    .S(_26388_),
    .Z(_05985_));
 MUX2_X1 _58327_ (.A(lce_data_cmd_i[493]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [493]),
    .S(_26388_),
    .Z(_05986_));
 MUX2_X1 _58328_ (.A(lce_data_cmd_i[494]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [494]),
    .S(_26388_),
    .Z(_05987_));
 MUX2_X1 _58329_ (.A(lce_data_cmd_i[495]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [495]),
    .S(_26388_),
    .Z(_05988_));
 MUX2_X1 _58330_ (.A(lce_data_cmd_i[496]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [496]),
    .S(_26388_),
    .Z(_05989_));
 MUX2_X1 _58331_ (.A(lce_data_cmd_i[497]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [497]),
    .S(_26388_),
    .Z(_05990_));
 BUF_X8 _58332_ (.A(_26383_),
    .Z(_26389_));
 MUX2_X1 _58333_ (.A(lce_data_cmd_i[498]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [498]),
    .S(_26389_),
    .Z(_05991_));
 MUX2_X1 _58334_ (.A(lce_data_cmd_i[499]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [499]),
    .S(_26389_),
    .Z(_05992_));
 MUX2_X1 _58335_ (.A(lce_data_cmd_i[500]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [500]),
    .S(_26389_),
    .Z(_05995_));
 MUX2_X1 _58336_ (.A(lce_data_cmd_i[501]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [501]),
    .S(_26389_),
    .Z(_05996_));
 MUX2_X1 _58337_ (.A(lce_data_cmd_i[502]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [502]),
    .S(_26389_),
    .Z(_05997_));
 MUX2_X1 _58338_ (.A(lce_data_cmd_i[503]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [503]),
    .S(_26389_),
    .Z(_05998_));
 MUX2_X1 _58339_ (.A(lce_data_cmd_i[504]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [504]),
    .S(_26389_),
    .Z(_05999_));
 MUX2_X1 _58340_ (.A(lce_data_cmd_i[505]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [505]),
    .S(_26389_),
    .Z(_06000_));
 MUX2_X1 _58341_ (.A(lce_data_cmd_i[506]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [506]),
    .S(_26389_),
    .Z(_06001_));
 MUX2_X1 _58342_ (.A(lce_data_cmd_i[507]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [507]),
    .S(_26389_),
    .Z(_06002_));
 BUF_X8 _58343_ (.A(_26383_),
    .Z(_26390_));
 MUX2_X1 _58344_ (.A(lce_data_cmd_i[508]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [508]),
    .S(_26390_),
    .Z(_06003_));
 MUX2_X1 _58345_ (.A(lce_data_cmd_i[509]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [509]),
    .S(_26390_),
    .Z(_06004_));
 MUX2_X1 _58346_ (.A(lce_data_cmd_i[510]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [510]),
    .S(_26390_),
    .Z(_06006_));
 MUX2_X1 _58347_ (.A(lce_data_cmd_i[511]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [511]),
    .S(_26390_),
    .Z(_06007_));
 MUX2_X1 _58348_ (.A(lce_data_cmd_i[512]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [512]),
    .S(_26390_),
    .Z(_06008_));
 MUX2_X1 _58349_ (.A(lce_data_cmd_i[513]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [513]),
    .S(_26390_),
    .Z(_06009_));
 MUX2_X1 _58350_ (.A(lce_data_cmd_i[514]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [514]),
    .S(_26390_),
    .Z(_06010_));
 MUX2_X1 _58351_ (.A(lce_data_cmd_i[515]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [515]),
    .S(_26390_),
    .Z(_06011_));
 MUX2_X1 _58352_ (.A(lce_data_cmd_i[516]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [516]),
    .S(_26390_),
    .Z(_06012_));
 MUX2_X1 _58353_ (.A(lce_data_cmd_i[517]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [517]),
    .S(_26390_),
    .Z(_06013_));
 BUF_X8 _58354_ (.A(_26383_),
    .Z(_26391_));
 MUX2_X1 _58355_ (.A(lce_data_cmd_i[1]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1]),
    .S(_26391_),
    .Z(_05661_));
 MUX2_X1 _58356_ (.A(lce_data_cmd_i[320]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [320]),
    .S(_26391_),
    .Z(_05795_));
 MUX2_X1 _58357_ (.A(lce_data_cmd_i[321]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [321]),
    .S(_26391_),
    .Z(_05796_));
 MUX2_X1 _58358_ (.A(lce_data_cmd_i[322]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [322]),
    .S(_26391_),
    .Z(_05797_));
 MUX2_X1 _58359_ (.A(lce_data_cmd_i[323]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [323]),
    .S(_26391_),
    .Z(_05798_));
 MUX2_X1 _58360_ (.A(lce_data_cmd_i[324]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [324]),
    .S(_26391_),
    .Z(_05799_));
 MUX2_X1 _58361_ (.A(lce_data_cmd_i[325]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [325]),
    .S(_26391_),
    .Z(_05800_));
 MUX2_X1 _58362_ (.A(lce_data_cmd_i[326]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [326]),
    .S(_26391_),
    .Z(_05801_));
 MUX2_X1 _58363_ (.A(lce_data_cmd_i[327]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [327]),
    .S(_26391_),
    .Z(_05802_));
 MUX2_X1 _58364_ (.A(lce_data_cmd_i[328]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [328]),
    .S(_26391_),
    .Z(_05803_));
 BUF_X8 _58365_ (.A(_26383_),
    .Z(_26392_));
 MUX2_X1 _58366_ (.A(lce_data_cmd_i[329]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [329]),
    .S(_26392_),
    .Z(_05804_));
 MUX2_X1 _58367_ (.A(lce_data_cmd_i[330]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [330]),
    .S(_26392_),
    .Z(_05806_));
 MUX2_X1 _58368_ (.A(lce_data_cmd_i[331]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [331]),
    .S(_26392_),
    .Z(_05807_));
 MUX2_X1 _58369_ (.A(lce_data_cmd_i[332]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [332]),
    .S(_26392_),
    .Z(_05808_));
 MUX2_X1 _58370_ (.A(lce_data_cmd_i[333]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [333]),
    .S(_26392_),
    .Z(_05809_));
 MUX2_X1 _58371_ (.A(lce_data_cmd_i[334]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [334]),
    .S(_26392_),
    .Z(_05810_));
 MUX2_X1 _58372_ (.A(lce_data_cmd_i[335]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [335]),
    .S(_26392_),
    .Z(_05811_));
 MUX2_X1 _58373_ (.A(lce_data_cmd_i[336]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [336]),
    .S(_26392_),
    .Z(_05812_));
 MUX2_X1 _58374_ (.A(lce_data_cmd_i[337]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [337]),
    .S(_26392_),
    .Z(_05813_));
 MUX2_X1 _58375_ (.A(lce_data_cmd_i[338]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [338]),
    .S(_26392_),
    .Z(_05814_));
 BUF_X8 _58376_ (.A(_26383_),
    .Z(_26393_));
 MUX2_X1 _58377_ (.A(lce_data_cmd_i[339]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [339]),
    .S(_26393_),
    .Z(_05815_));
 MUX2_X1 _58378_ (.A(lce_data_cmd_i[340]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [340]),
    .S(_26393_),
    .Z(_05817_));
 MUX2_X1 _58379_ (.A(lce_data_cmd_i[341]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [341]),
    .S(_26393_),
    .Z(_05818_));
 MUX2_X1 _58380_ (.A(lce_data_cmd_i[342]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [342]),
    .S(_26393_),
    .Z(_05819_));
 MUX2_X1 _58381_ (.A(lce_data_cmd_i[343]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [343]),
    .S(_26393_),
    .Z(_05820_));
 MUX2_X1 _58382_ (.A(lce_data_cmd_i[344]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [344]),
    .S(_26393_),
    .Z(_05821_));
 MUX2_X1 _58383_ (.A(lce_data_cmd_i[345]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [345]),
    .S(_26393_),
    .Z(_05822_));
 MUX2_X1 _58384_ (.A(lce_data_cmd_i[346]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [346]),
    .S(_26393_),
    .Z(_05823_));
 MUX2_X1 _58385_ (.A(lce_data_cmd_i[347]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [347]),
    .S(_26393_),
    .Z(_05824_));
 MUX2_X1 _58386_ (.A(lce_data_cmd_i[348]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [348]),
    .S(_26393_),
    .Z(_05825_));
 BUF_X32 _58387_ (.A(_26382_),
    .Z(_26394_));
 BUF_X8 _58388_ (.A(_26394_),
    .Z(_26395_));
 MUX2_X1 _58389_ (.A(lce_data_cmd_i[349]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [349]),
    .S(_26395_),
    .Z(_05826_));
 MUX2_X1 _58390_ (.A(lce_data_cmd_i[350]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [350]),
    .S(_26395_),
    .Z(_05828_));
 MUX2_X1 _58391_ (.A(lce_data_cmd_i[351]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [351]),
    .S(_26395_),
    .Z(_05829_));
 MUX2_X1 _58392_ (.A(lce_data_cmd_i[352]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [352]),
    .S(_26395_),
    .Z(_05830_));
 MUX2_X1 _58393_ (.A(lce_data_cmd_i[353]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [353]),
    .S(_26395_),
    .Z(_05831_));
 MUX2_X1 _58394_ (.A(lce_data_cmd_i[354]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [354]),
    .S(_26395_),
    .Z(_05832_));
 MUX2_X1 _58395_ (.A(lce_data_cmd_i[355]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [355]),
    .S(_26395_),
    .Z(_05833_));
 MUX2_X1 _58396_ (.A(lce_data_cmd_i[356]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [356]),
    .S(_26395_),
    .Z(_05834_));
 MUX2_X1 _58397_ (.A(lce_data_cmd_i[357]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [357]),
    .S(_26395_),
    .Z(_05835_));
 MUX2_X1 _58398_ (.A(lce_data_cmd_i[358]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [358]),
    .S(_26395_),
    .Z(_05836_));
 BUF_X8 _58399_ (.A(_26394_),
    .Z(_26396_));
 MUX2_X1 _58400_ (.A(lce_data_cmd_i[359]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [359]),
    .S(_26396_),
    .Z(_05837_));
 MUX2_X1 _58401_ (.A(lce_data_cmd_i[360]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [360]),
    .S(_26396_),
    .Z(_05839_));
 MUX2_X1 _58402_ (.A(lce_data_cmd_i[361]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [361]),
    .S(_26396_),
    .Z(_05840_));
 MUX2_X1 _58403_ (.A(lce_data_cmd_i[362]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [362]),
    .S(_26396_),
    .Z(_05841_));
 MUX2_X1 _58404_ (.A(lce_data_cmd_i[363]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [363]),
    .S(_26396_),
    .Z(_05842_));
 MUX2_X1 _58405_ (.A(lce_data_cmd_i[364]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [364]),
    .S(_26396_),
    .Z(_05843_));
 MUX2_X1 _58406_ (.A(lce_data_cmd_i[365]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [365]),
    .S(_26396_),
    .Z(_05844_));
 MUX2_X1 _58407_ (.A(lce_data_cmd_i[366]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [366]),
    .S(_26396_),
    .Z(_05845_));
 MUX2_X1 _58408_ (.A(lce_data_cmd_i[367]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [367]),
    .S(_26396_),
    .Z(_05846_));
 MUX2_X1 _58409_ (.A(lce_data_cmd_i[368]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [368]),
    .S(_26396_),
    .Z(_05847_));
 BUF_X8 _58410_ (.A(_26394_),
    .Z(_26397_));
 MUX2_X1 _58411_ (.A(lce_data_cmd_i[369]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [369]),
    .S(_26397_),
    .Z(_05848_));
 MUX2_X1 _58412_ (.A(lce_data_cmd_i[370]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [370]),
    .S(_26397_),
    .Z(_05850_));
 MUX2_X1 _58413_ (.A(lce_data_cmd_i[371]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [371]),
    .S(_26397_),
    .Z(_05851_));
 MUX2_X1 _58414_ (.A(lce_data_cmd_i[372]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [372]),
    .S(_26397_),
    .Z(_05852_));
 MUX2_X1 _58415_ (.A(lce_data_cmd_i[373]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [373]),
    .S(_26397_),
    .Z(_05853_));
 MUX2_X1 _58416_ (.A(lce_data_cmd_i[374]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [374]),
    .S(_26397_),
    .Z(_05854_));
 MUX2_X1 _58417_ (.A(lce_data_cmd_i[375]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [375]),
    .S(_26397_),
    .Z(_05855_));
 MUX2_X1 _58418_ (.A(lce_data_cmd_i[376]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [376]),
    .S(_26397_),
    .Z(_05856_));
 MUX2_X1 _58419_ (.A(lce_data_cmd_i[377]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [377]),
    .S(_26397_),
    .Z(_05857_));
 MUX2_X1 _58420_ (.A(lce_data_cmd_i[378]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [378]),
    .S(_26397_),
    .Z(_05858_));
 BUF_X8 _58421_ (.A(_26394_),
    .Z(_26398_));
 MUX2_X1 _58422_ (.A(lce_data_cmd_i[379]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [379]),
    .S(_26398_),
    .Z(_05859_));
 MUX2_X1 _58423_ (.A(lce_data_cmd_i[380]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [380]),
    .S(_26398_),
    .Z(_05861_));
 MUX2_X1 _58424_ (.A(lce_data_cmd_i[381]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [381]),
    .S(_26398_),
    .Z(_05862_));
 MUX2_X1 _58425_ (.A(lce_data_cmd_i[382]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [382]),
    .S(_26398_),
    .Z(_05863_));
 MUX2_X1 _58426_ (.A(lce_data_cmd_i[383]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [383]),
    .S(_26398_),
    .Z(_05864_));
 MUX2_X1 _58427_ (.A(lce_data_cmd_i[384]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [384]),
    .S(_26398_),
    .Z(_05865_));
 MUX2_X1 _58428_ (.A(lce_data_cmd_i[385]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [385]),
    .S(_26398_),
    .Z(_05866_));
 MUX2_X1 _58429_ (.A(lce_data_cmd_i[386]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [386]),
    .S(_26398_),
    .Z(_05867_));
 MUX2_X1 _58430_ (.A(lce_data_cmd_i[387]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [387]),
    .S(_26398_),
    .Z(_05868_));
 MUX2_X1 _58431_ (.A(lce_data_cmd_i[388]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [388]),
    .S(_26398_),
    .Z(_05869_));
 BUF_X16 _58432_ (.A(_26394_),
    .Z(_26399_));
 MUX2_X1 _58433_ (.A(lce_data_cmd_i[389]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [389]),
    .S(_26399_),
    .Z(_05870_));
 MUX2_X1 _58434_ (.A(lce_data_cmd_i[390]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [390]),
    .S(_26399_),
    .Z(_05872_));
 MUX2_X1 _58435_ (.A(lce_data_cmd_i[391]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [391]),
    .S(_26399_),
    .Z(_05873_));
 MUX2_X1 _58436_ (.A(lce_data_cmd_i[392]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [392]),
    .S(_26399_),
    .Z(_05874_));
 MUX2_X1 _58437_ (.A(lce_data_cmd_i[393]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [393]),
    .S(_26399_),
    .Z(_05875_));
 MUX2_X1 _58438_ (.A(lce_data_cmd_i[394]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [394]),
    .S(_26399_),
    .Z(_05876_));
 MUX2_X1 _58439_ (.A(lce_data_cmd_i[395]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [395]),
    .S(_26399_),
    .Z(_05877_));
 MUX2_X1 _58440_ (.A(lce_data_cmd_i[396]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [396]),
    .S(_26399_),
    .Z(_05878_));
 MUX2_X1 _58441_ (.A(lce_data_cmd_i[397]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [397]),
    .S(_26399_),
    .Z(_05879_));
 MUX2_X1 _58442_ (.A(lce_data_cmd_i[398]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [398]),
    .S(_26399_),
    .Z(_05880_));
 BUF_X8 _58443_ (.A(_26394_),
    .Z(_26400_));
 MUX2_X1 _58444_ (.A(lce_data_cmd_i[399]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [399]),
    .S(_26400_),
    .Z(_05881_));
 MUX2_X1 _58445_ (.A(lce_data_cmd_i[400]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [400]),
    .S(_26400_),
    .Z(_05884_));
 MUX2_X1 _58446_ (.A(lce_data_cmd_i[401]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [401]),
    .S(_26400_),
    .Z(_05885_));
 MUX2_X1 _58447_ (.A(lce_data_cmd_i[402]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [402]),
    .S(_26400_),
    .Z(_05886_));
 MUX2_X1 _58448_ (.A(lce_data_cmd_i[403]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [403]),
    .S(_26400_),
    .Z(_05887_));
 MUX2_X1 _58449_ (.A(lce_data_cmd_i[404]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [404]),
    .S(_26400_),
    .Z(_05888_));
 MUX2_X1 _58450_ (.A(lce_data_cmd_i[405]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [405]),
    .S(_26400_),
    .Z(_05889_));
 MUX2_X1 _58451_ (.A(lce_data_cmd_i[406]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [406]),
    .S(_26400_),
    .Z(_05890_));
 MUX2_X1 _58452_ (.A(lce_data_cmd_i[407]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [407]),
    .S(_26400_),
    .Z(_05891_));
 MUX2_X1 _58453_ (.A(lce_data_cmd_i[408]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [408]),
    .S(_26400_),
    .Z(_05892_));
 BUF_X4 _58454_ (.A(_26394_),
    .Z(_26401_));
 MUX2_X1 _58455_ (.A(lce_data_cmd_i[409]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [409]),
    .S(_26401_),
    .Z(_05893_));
 MUX2_X1 _58456_ (.A(lce_data_cmd_i[410]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [410]),
    .S(_26401_),
    .Z(_05895_));
 MUX2_X1 _58457_ (.A(lce_data_cmd_i[411]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [411]),
    .S(_26401_),
    .Z(_05896_));
 MUX2_X1 _58458_ (.A(lce_data_cmd_i[412]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [412]),
    .S(_26401_),
    .Z(_05897_));
 MUX2_X1 _58459_ (.A(lce_data_cmd_i[413]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [413]),
    .S(_26401_),
    .Z(_05898_));
 MUX2_X1 _58460_ (.A(lce_data_cmd_i[414]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [414]),
    .S(_26401_),
    .Z(_05899_));
 MUX2_X1 _58461_ (.A(lce_data_cmd_i[415]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [415]),
    .S(_26401_),
    .Z(_05900_));
 MUX2_X1 _58462_ (.A(lce_data_cmd_i[416]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [416]),
    .S(_26401_),
    .Z(_05901_));
 MUX2_X1 _58463_ (.A(lce_data_cmd_i[417]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [417]),
    .S(_26401_),
    .Z(_05902_));
 MUX2_X1 _58464_ (.A(lce_data_cmd_i[418]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [418]),
    .S(_26401_),
    .Z(_05903_));
 BUF_X8 _58465_ (.A(_26394_),
    .Z(_26402_));
 MUX2_X1 _58466_ (.A(lce_data_cmd_i[2]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [2]),
    .S(_26402_),
    .Z(_05772_));
 MUX2_X1 _58467_ (.A(lce_data_cmd_i[221]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [221]),
    .S(_26402_),
    .Z(_05685_));
 MUX2_X1 _58468_ (.A(lce_data_cmd_i[222]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [222]),
    .S(_26402_),
    .Z(_05686_));
 MUX2_X1 _58469_ (.A(lce_data_cmd_i[223]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [223]),
    .S(_26402_),
    .Z(_05687_));
 MUX2_X1 _58470_ (.A(lce_data_cmd_i[224]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [224]),
    .S(_26402_),
    .Z(_05688_));
 MUX2_X1 _58471_ (.A(lce_data_cmd_i[225]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [225]),
    .S(_26402_),
    .Z(_05689_));
 MUX2_X1 _58472_ (.A(lce_data_cmd_i[226]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [226]),
    .S(_26402_),
    .Z(_05690_));
 MUX2_X1 _58473_ (.A(lce_data_cmd_i[227]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [227]),
    .S(_26402_),
    .Z(_05691_));
 MUX2_X1 _58474_ (.A(lce_data_cmd_i[228]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [228]),
    .S(_26402_),
    .Z(_05692_));
 MUX2_X1 _58475_ (.A(lce_data_cmd_i[229]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [229]),
    .S(_26402_),
    .Z(_05693_));
 BUF_X8 _58476_ (.A(_26394_),
    .Z(_26403_));
 MUX2_X1 _58477_ (.A(lce_data_cmd_i[230]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [230]),
    .S(_26403_),
    .Z(_05695_));
 MUX2_X1 _58478_ (.A(lce_data_cmd_i[231]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [231]),
    .S(_26403_),
    .Z(_05696_));
 MUX2_X1 _58479_ (.A(lce_data_cmd_i[232]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [232]),
    .S(_26403_),
    .Z(_05697_));
 MUX2_X1 _58480_ (.A(lce_data_cmd_i[233]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [233]),
    .S(_26403_),
    .Z(_05698_));
 MUX2_X1 _58481_ (.A(lce_data_cmd_i[234]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [234]),
    .S(_26403_),
    .Z(_05699_));
 MUX2_X1 _58482_ (.A(lce_data_cmd_i[235]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [235]),
    .S(_26403_),
    .Z(_05700_));
 MUX2_X1 _58483_ (.A(lce_data_cmd_i[236]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [236]),
    .S(_26403_),
    .Z(_05701_));
 MUX2_X1 _58484_ (.A(lce_data_cmd_i[237]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [237]),
    .S(_26403_),
    .Z(_05702_));
 MUX2_X1 _58485_ (.A(lce_data_cmd_i[238]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [238]),
    .S(_26403_),
    .Z(_05703_));
 MUX2_X1 _58486_ (.A(lce_data_cmd_i[239]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [239]),
    .S(_26403_),
    .Z(_05704_));
 BUF_X8 _58487_ (.A(_26394_),
    .Z(_26404_));
 MUX2_X1 _58488_ (.A(lce_data_cmd_i[240]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [240]),
    .S(_26404_),
    .Z(_05706_));
 MUX2_X1 _58489_ (.A(lce_data_cmd_i[241]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [241]),
    .S(_26404_),
    .Z(_05707_));
 MUX2_X1 _58490_ (.A(lce_data_cmd_i[242]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [242]),
    .S(_26404_),
    .Z(_05708_));
 MUX2_X1 _58491_ (.A(lce_data_cmd_i[243]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [243]),
    .S(_26404_),
    .Z(_05709_));
 MUX2_X1 _58492_ (.A(lce_data_cmd_i[244]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [244]),
    .S(_26404_),
    .Z(_05710_));
 MUX2_X1 _58493_ (.A(lce_data_cmd_i[245]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [245]),
    .S(_26404_),
    .Z(_05711_));
 MUX2_X1 _58494_ (.A(lce_data_cmd_i[246]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [246]),
    .S(_26404_),
    .Z(_05712_));
 MUX2_X1 _58495_ (.A(lce_data_cmd_i[247]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [247]),
    .S(_26404_),
    .Z(_05713_));
 MUX2_X1 _58496_ (.A(lce_data_cmd_i[248]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [248]),
    .S(_26404_),
    .Z(_05714_));
 MUX2_X1 _58497_ (.A(lce_data_cmd_i[249]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [249]),
    .S(_26404_),
    .Z(_05715_));
 BUF_X32 _58498_ (.A(_26377_),
    .Z(_26405_));
 BUF_X8 _58499_ (.A(_26405_),
    .Z(_26406_));
 MUX2_X1 _58500_ (.A(lce_data_cmd_i[250]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [250]),
    .S(_26406_),
    .Z(_05717_));
 MUX2_X1 _58501_ (.A(lce_data_cmd_i[251]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [251]),
    .S(_26406_),
    .Z(_05718_));
 MUX2_X1 _58502_ (.A(lce_data_cmd_i[252]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [252]),
    .S(_26406_),
    .Z(_05719_));
 MUX2_X1 _58503_ (.A(lce_data_cmd_i[253]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [253]),
    .S(_26406_),
    .Z(_05720_));
 MUX2_X1 _58504_ (.A(lce_data_cmd_i[254]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [254]),
    .S(_26406_),
    .Z(_05721_));
 MUX2_X1 _58505_ (.A(lce_data_cmd_i[255]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [255]),
    .S(_26406_),
    .Z(_05722_));
 MUX2_X1 _58506_ (.A(lce_data_cmd_i[256]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [256]),
    .S(_26406_),
    .Z(_05723_));
 MUX2_X1 _58507_ (.A(lce_data_cmd_i[257]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [257]),
    .S(_26406_),
    .Z(_05724_));
 MUX2_X1 _58508_ (.A(lce_data_cmd_i[258]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [258]),
    .S(_26406_),
    .Z(_05725_));
 MUX2_X1 _58509_ (.A(lce_data_cmd_i[259]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [259]),
    .S(_26406_),
    .Z(_05726_));
 BUF_X16 _58510_ (.A(_26405_),
    .Z(_26407_));
 MUX2_X1 _58511_ (.A(lce_data_cmd_i[260]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [260]),
    .S(_26407_),
    .Z(_05728_));
 MUX2_X1 _58512_ (.A(lce_data_cmd_i[261]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [261]),
    .S(_26407_),
    .Z(_05729_));
 MUX2_X1 _58513_ (.A(lce_data_cmd_i[262]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [262]),
    .S(_26407_),
    .Z(_05730_));
 MUX2_X1 _58514_ (.A(lce_data_cmd_i[263]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [263]),
    .S(_26407_),
    .Z(_05731_));
 MUX2_X1 _58515_ (.A(lce_data_cmd_i[264]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [264]),
    .S(_26407_),
    .Z(_05732_));
 MUX2_X1 _58516_ (.A(lce_data_cmd_i[265]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [265]),
    .S(_26407_),
    .Z(_05733_));
 MUX2_X1 _58517_ (.A(lce_data_cmd_i[266]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [266]),
    .S(_26407_),
    .Z(_05734_));
 MUX2_X1 _58518_ (.A(lce_data_cmd_i[267]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [267]),
    .S(_26407_),
    .Z(_05735_));
 MUX2_X1 _58519_ (.A(lce_data_cmd_i[268]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [268]),
    .S(_26407_),
    .Z(_05736_));
 MUX2_X1 _58520_ (.A(lce_data_cmd_i[269]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [269]),
    .S(_26407_),
    .Z(_05737_));
 BUF_X8 _58521_ (.A(_26405_),
    .Z(_26408_));
 MUX2_X1 _58522_ (.A(lce_data_cmd_i[270]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [270]),
    .S(_26408_),
    .Z(_05739_));
 MUX2_X1 _58523_ (.A(lce_data_cmd_i[271]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [271]),
    .S(_26408_),
    .Z(_05740_));
 MUX2_X1 _58524_ (.A(lce_data_cmd_i[272]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [272]),
    .S(_26408_),
    .Z(_05741_));
 MUX2_X1 _58525_ (.A(lce_data_cmd_i[273]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [273]),
    .S(_26408_),
    .Z(_05742_));
 MUX2_X1 _58526_ (.A(lce_data_cmd_i[274]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [274]),
    .S(_26408_),
    .Z(_05743_));
 MUX2_X1 _58527_ (.A(lce_data_cmd_i[275]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [275]),
    .S(_26408_),
    .Z(_05744_));
 MUX2_X1 _58528_ (.A(lce_data_cmd_i[276]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [276]),
    .S(_26408_),
    .Z(_05745_));
 MUX2_X1 _58529_ (.A(lce_data_cmd_i[277]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [277]),
    .S(_26408_),
    .Z(_05746_));
 MUX2_X1 _58530_ (.A(lce_data_cmd_i[278]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [278]),
    .S(_26408_),
    .Z(_05747_));
 MUX2_X1 _58531_ (.A(lce_data_cmd_i[279]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [279]),
    .S(_26408_),
    .Z(_05748_));
 BUF_X4 _58532_ (.A(_26405_),
    .Z(_26409_));
 MUX2_X1 _58533_ (.A(lce_data_cmd_i[280]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [280]),
    .S(_26409_),
    .Z(_05750_));
 MUX2_X1 _58534_ (.A(lce_data_cmd_i[281]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [281]),
    .S(_26409_),
    .Z(_05751_));
 MUX2_X1 _58535_ (.A(lce_data_cmd_i[282]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [282]),
    .S(_26409_),
    .Z(_05752_));
 MUX2_X1 _58536_ (.A(lce_data_cmd_i[283]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [283]),
    .S(_26409_),
    .Z(_05753_));
 MUX2_X1 _58537_ (.A(lce_data_cmd_i[284]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [284]),
    .S(_26409_),
    .Z(_05754_));
 MUX2_X1 _58538_ (.A(lce_data_cmd_i[285]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [285]),
    .S(_26409_),
    .Z(_05755_));
 MUX2_X1 _58539_ (.A(lce_data_cmd_i[286]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [286]),
    .S(_26409_),
    .Z(_05756_));
 MUX2_X1 _58540_ (.A(lce_data_cmd_i[287]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [287]),
    .S(_26409_),
    .Z(_05757_));
 MUX2_X1 _58541_ (.A(lce_data_cmd_i[288]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [288]),
    .S(_26409_),
    .Z(_05758_));
 MUX2_X1 _58542_ (.A(lce_data_cmd_i[289]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [289]),
    .S(_26409_),
    .Z(_05759_));
 BUF_X8 _58543_ (.A(_26405_),
    .Z(_26410_));
 MUX2_X1 _58544_ (.A(lce_data_cmd_i[290]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [290]),
    .S(_26410_),
    .Z(_05761_));
 MUX2_X1 _58545_ (.A(lce_data_cmd_i[291]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [291]),
    .S(_26410_),
    .Z(_05762_));
 MUX2_X1 _58546_ (.A(lce_data_cmd_i[292]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [292]),
    .S(_26410_),
    .Z(_05763_));
 MUX2_X1 _58547_ (.A(lce_data_cmd_i[293]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [293]),
    .S(_26410_),
    .Z(_05764_));
 MUX2_X1 _58548_ (.A(lce_data_cmd_i[294]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [294]),
    .S(_26410_),
    .Z(_05765_));
 MUX2_X1 _58549_ (.A(lce_data_cmd_i[295]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [295]),
    .S(_26410_),
    .Z(_05766_));
 MUX2_X1 _58550_ (.A(lce_data_cmd_i[296]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [296]),
    .S(_26410_),
    .Z(_05767_));
 MUX2_X1 _58551_ (.A(lce_data_cmd_i[297]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [297]),
    .S(_26410_),
    .Z(_05768_));
 MUX2_X1 _58552_ (.A(lce_data_cmd_i[298]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [298]),
    .S(_26410_),
    .Z(_05769_));
 MUX2_X1 _58553_ (.A(lce_data_cmd_i[299]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [299]),
    .S(_26410_),
    .Z(_05770_));
 BUF_X8 _58554_ (.A(_26405_),
    .Z(_26411_));
 MUX2_X1 _58555_ (.A(lce_data_cmd_i[300]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [300]),
    .S(_26411_),
    .Z(_05773_));
 MUX2_X1 _58556_ (.A(lce_data_cmd_i[301]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [301]),
    .S(_26411_),
    .Z(_05774_));
 MUX2_X1 _58557_ (.A(lce_data_cmd_i[302]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [302]),
    .S(_26411_),
    .Z(_05775_));
 MUX2_X1 _58558_ (.A(lce_data_cmd_i[303]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [303]),
    .S(_26411_),
    .Z(_05776_));
 MUX2_X1 _58559_ (.A(lce_data_cmd_i[304]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [304]),
    .S(_26411_),
    .Z(_05777_));
 MUX2_X1 _58560_ (.A(lce_data_cmd_i[305]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [305]),
    .S(_26411_),
    .Z(_05778_));
 MUX2_X1 _58561_ (.A(lce_data_cmd_i[306]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [306]),
    .S(_26411_),
    .Z(_05779_));
 MUX2_X1 _58562_ (.A(lce_data_cmd_i[307]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [307]),
    .S(_26411_),
    .Z(_05780_));
 MUX2_X1 _58563_ (.A(lce_data_cmd_i[308]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [308]),
    .S(_26411_),
    .Z(_05781_));
 MUX2_X1 _58564_ (.A(lce_data_cmd_i[309]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [309]),
    .S(_26411_),
    .Z(_05782_));
 BUF_X16 _58565_ (.A(_26405_),
    .Z(_26412_));
 MUX2_X1 _58566_ (.A(lce_data_cmd_i[310]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [310]),
    .S(_26412_),
    .Z(_05784_));
 MUX2_X1 _58567_ (.A(lce_data_cmd_i[311]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [311]),
    .S(_26412_),
    .Z(_05785_));
 MUX2_X1 _58568_ (.A(lce_data_cmd_i[312]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [312]),
    .S(_26412_),
    .Z(_05786_));
 MUX2_X1 _58569_ (.A(lce_data_cmd_i[313]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [313]),
    .S(_26412_),
    .Z(_05787_));
 MUX2_X1 _58570_ (.A(lce_data_cmd_i[314]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [314]),
    .S(_26412_),
    .Z(_05788_));
 MUX2_X1 _58571_ (.A(lce_data_cmd_i[315]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [315]),
    .S(_26412_),
    .Z(_05789_));
 MUX2_X1 _58572_ (.A(lce_data_cmd_i[316]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [316]),
    .S(_26412_),
    .Z(_05790_));
 MUX2_X1 _58573_ (.A(lce_data_cmd_i[317]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [317]),
    .S(_26412_),
    .Z(_05791_));
 MUX2_X1 _58574_ (.A(lce_data_cmd_i[318]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [318]),
    .S(_26412_),
    .Z(_05792_));
 MUX2_X1 _58575_ (.A(lce_data_cmd_i[319]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [319]),
    .S(_26412_),
    .Z(_05793_));
 BUF_X8 _58576_ (.A(_26405_),
    .Z(_26413_));
 MUX2_X1 _58577_ (.A(lce_data_cmd_i[3]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [3]),
    .S(_26413_),
    .Z(_05883_));
 MUX2_X1 _58578_ (.A(lce_data_cmd_i[122]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [122]),
    .S(_26413_),
    .Z(_05575_));
 MUX2_X1 _58579_ (.A(lce_data_cmd_i[123]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [123]),
    .S(_26413_),
    .Z(_05576_));
 MUX2_X1 _58580_ (.A(lce_data_cmd_i[124]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [124]),
    .S(_26413_),
    .Z(_05577_));
 MUX2_X1 _58581_ (.A(lce_data_cmd_i[125]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [125]),
    .S(_26413_),
    .Z(_05578_));
 MUX2_X1 _58582_ (.A(lce_data_cmd_i[126]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [126]),
    .S(_26413_),
    .Z(_05579_));
 MUX2_X1 _58583_ (.A(lce_data_cmd_i[127]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [127]),
    .S(_26413_),
    .Z(_05580_));
 MUX2_X1 _58584_ (.A(lce_data_cmd_i[128]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [128]),
    .S(_26413_),
    .Z(_05581_));
 MUX2_X1 _58585_ (.A(lce_data_cmd_i[129]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [129]),
    .S(_26413_),
    .Z(_05582_));
 MUX2_X1 _58586_ (.A(lce_data_cmd_i[130]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [130]),
    .S(_26413_),
    .Z(_05584_));
 BUF_X8 _58587_ (.A(_26405_),
    .Z(_26414_));
 MUX2_X1 _58588_ (.A(lce_data_cmd_i[131]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [131]),
    .S(_26414_),
    .Z(_05585_));
 MUX2_X1 _58589_ (.A(lce_data_cmd_i[132]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [132]),
    .S(_26414_),
    .Z(_05586_));
 MUX2_X1 _58590_ (.A(lce_data_cmd_i[133]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [133]),
    .S(_26414_),
    .Z(_05587_));
 MUX2_X1 _58591_ (.A(lce_data_cmd_i[134]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [134]),
    .S(_26414_),
    .Z(_05588_));
 MUX2_X1 _58592_ (.A(lce_data_cmd_i[135]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [135]),
    .S(_26414_),
    .Z(_05589_));
 MUX2_X1 _58593_ (.A(lce_data_cmd_i[136]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [136]),
    .S(_26414_),
    .Z(_05590_));
 MUX2_X1 _58594_ (.A(lce_data_cmd_i[137]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [137]),
    .S(_26414_),
    .Z(_05591_));
 MUX2_X1 _58595_ (.A(lce_data_cmd_i[138]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [138]),
    .S(_26414_),
    .Z(_05592_));
 MUX2_X1 _58596_ (.A(lce_data_cmd_i[139]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [139]),
    .S(_26414_),
    .Z(_05593_));
 MUX2_X1 _58597_ (.A(lce_data_cmd_i[140]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [140]),
    .S(_26414_),
    .Z(_05595_));
 BUF_X8 _58598_ (.A(_26405_),
    .Z(_26415_));
 MUX2_X1 _58599_ (.A(lce_data_cmd_i[141]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [141]),
    .S(_26415_),
    .Z(_05596_));
 MUX2_X1 _58600_ (.A(lce_data_cmd_i[142]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [142]),
    .S(_26415_),
    .Z(_05597_));
 MUX2_X1 _58601_ (.A(lce_data_cmd_i[143]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [143]),
    .S(_26415_),
    .Z(_05598_));
 MUX2_X1 _58602_ (.A(lce_data_cmd_i[144]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [144]),
    .S(_26415_),
    .Z(_05599_));
 MUX2_X1 _58603_ (.A(lce_data_cmd_i[145]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [145]),
    .S(_26415_),
    .Z(_05600_));
 MUX2_X1 _58604_ (.A(lce_data_cmd_i[146]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [146]),
    .S(_26415_),
    .Z(_05601_));
 MUX2_X1 _58605_ (.A(lce_data_cmd_i[147]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [147]),
    .S(_26415_),
    .Z(_05602_));
 MUX2_X1 _58606_ (.A(lce_data_cmd_i[148]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [148]),
    .S(_26415_),
    .Z(_05603_));
 MUX2_X1 _58607_ (.A(lce_data_cmd_i[149]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [149]),
    .S(_26415_),
    .Z(_05604_));
 MUX2_X1 _58608_ (.A(lce_data_cmd_i[150]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [150]),
    .S(_26415_),
    .Z(_05606_));
 BUF_X32 _58609_ (.A(_26377_),
    .Z(_26416_));
 BUF_X8 _58610_ (.A(_26416_),
    .Z(_26417_));
 MUX2_X1 _58611_ (.A(lce_data_cmd_i[151]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [151]),
    .S(_26417_),
    .Z(_05607_));
 MUX2_X1 _58612_ (.A(lce_data_cmd_i[152]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [152]),
    .S(_26417_),
    .Z(_05608_));
 MUX2_X1 _58613_ (.A(lce_data_cmd_i[153]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [153]),
    .S(_26417_),
    .Z(_05609_));
 MUX2_X1 _58614_ (.A(lce_data_cmd_i[154]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [154]),
    .S(_26417_),
    .Z(_05610_));
 MUX2_X1 _58615_ (.A(lce_data_cmd_i[155]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [155]),
    .S(_26417_),
    .Z(_05611_));
 MUX2_X1 _58616_ (.A(lce_data_cmd_i[156]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [156]),
    .S(_26417_),
    .Z(_05612_));
 MUX2_X1 _58617_ (.A(lce_data_cmd_i[157]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [157]),
    .S(_26417_),
    .Z(_05613_));
 MUX2_X1 _58618_ (.A(lce_data_cmd_i[158]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [158]),
    .S(_26417_),
    .Z(_05614_));
 MUX2_X1 _58619_ (.A(lce_data_cmd_i[159]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [159]),
    .S(_26417_),
    .Z(_05615_));
 MUX2_X1 _58620_ (.A(lce_data_cmd_i[160]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [160]),
    .S(_26417_),
    .Z(_05617_));
 BUF_X8 _58621_ (.A(_26416_),
    .Z(_26418_));
 MUX2_X1 _58622_ (.A(lce_data_cmd_i[161]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [161]),
    .S(_26418_),
    .Z(_05618_));
 MUX2_X1 _58623_ (.A(lce_data_cmd_i[162]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [162]),
    .S(_26418_),
    .Z(_05619_));
 MUX2_X1 _58624_ (.A(lce_data_cmd_i[163]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [163]),
    .S(_26418_),
    .Z(_05620_));
 MUX2_X1 _58625_ (.A(lce_data_cmd_i[164]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [164]),
    .S(_26418_),
    .Z(_05621_));
 MUX2_X1 _58626_ (.A(lce_data_cmd_i[165]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [165]),
    .S(_26418_),
    .Z(_05622_));
 MUX2_X1 _58627_ (.A(lce_data_cmd_i[166]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [166]),
    .S(_26418_),
    .Z(_05623_));
 MUX2_X1 _58628_ (.A(lce_data_cmd_i[167]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [167]),
    .S(_26418_),
    .Z(_05624_));
 MUX2_X1 _58629_ (.A(lce_data_cmd_i[168]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [168]),
    .S(_26418_),
    .Z(_05625_));
 MUX2_X1 _58630_ (.A(lce_data_cmd_i[169]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [169]),
    .S(_26418_),
    .Z(_05626_));
 MUX2_X1 _58631_ (.A(lce_data_cmd_i[170]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [170]),
    .S(_26418_),
    .Z(_05628_));
 BUF_X4 _58632_ (.A(_26416_),
    .Z(_26419_));
 MUX2_X1 _58633_ (.A(lce_data_cmd_i[171]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [171]),
    .S(_26419_),
    .Z(_05629_));
 MUX2_X1 _58634_ (.A(lce_data_cmd_i[172]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [172]),
    .S(_26419_),
    .Z(_05630_));
 MUX2_X1 _58635_ (.A(lce_data_cmd_i[173]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [173]),
    .S(_26419_),
    .Z(_05631_));
 MUX2_X1 _58636_ (.A(lce_data_cmd_i[174]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [174]),
    .S(_26419_),
    .Z(_05632_));
 MUX2_X1 _58637_ (.A(lce_data_cmd_i[175]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [175]),
    .S(_26419_),
    .Z(_05633_));
 MUX2_X1 _58638_ (.A(lce_data_cmd_i[176]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [176]),
    .S(_26419_),
    .Z(_05634_));
 MUX2_X1 _58639_ (.A(lce_data_cmd_i[177]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [177]),
    .S(_26419_),
    .Z(_05635_));
 MUX2_X1 _58640_ (.A(lce_data_cmd_i[178]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [178]),
    .S(_26419_),
    .Z(_05636_));
 MUX2_X1 _58641_ (.A(lce_data_cmd_i[179]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [179]),
    .S(_26419_),
    .Z(_05637_));
 MUX2_X1 _58642_ (.A(lce_data_cmd_i[180]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [180]),
    .S(_26419_),
    .Z(_05639_));
 BUF_X8 _58643_ (.A(_26416_),
    .Z(_26420_));
 MUX2_X1 _58644_ (.A(lce_data_cmd_i[181]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [181]),
    .S(_26420_),
    .Z(_05640_));
 MUX2_X1 _58645_ (.A(lce_data_cmd_i[182]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [182]),
    .S(_26420_),
    .Z(_05641_));
 MUX2_X1 _58646_ (.A(lce_data_cmd_i[183]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [183]),
    .S(_26420_),
    .Z(_05642_));
 MUX2_X1 _58647_ (.A(lce_data_cmd_i[184]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [184]),
    .S(_26420_),
    .Z(_05643_));
 MUX2_X1 _58648_ (.A(lce_data_cmd_i[185]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [185]),
    .S(_26420_),
    .Z(_05644_));
 MUX2_X1 _58649_ (.A(lce_data_cmd_i[186]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [186]),
    .S(_26420_),
    .Z(_05645_));
 MUX2_X1 _58650_ (.A(lce_data_cmd_i[187]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [187]),
    .S(_26420_),
    .Z(_05646_));
 MUX2_X1 _58651_ (.A(lce_data_cmd_i[188]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [188]),
    .S(_26420_),
    .Z(_05647_));
 MUX2_X1 _58652_ (.A(lce_data_cmd_i[189]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [189]),
    .S(_26420_),
    .Z(_05648_));
 MUX2_X1 _58653_ (.A(lce_data_cmd_i[190]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [190]),
    .S(_26420_),
    .Z(_05650_));
 BUF_X8 _58654_ (.A(_26416_),
    .Z(_26421_));
 MUX2_X1 _58655_ (.A(lce_data_cmd_i[191]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [191]),
    .S(_26421_),
    .Z(_05651_));
 MUX2_X1 _58656_ (.A(lce_data_cmd_i[192]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [192]),
    .S(_26421_),
    .Z(_05652_));
 MUX2_X1 _58657_ (.A(lce_data_cmd_i[193]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [193]),
    .S(_26421_),
    .Z(_05653_));
 MUX2_X1 _58658_ (.A(lce_data_cmd_i[194]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [194]),
    .S(_26421_),
    .Z(_05654_));
 MUX2_X1 _58659_ (.A(lce_data_cmd_i[195]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [195]),
    .S(_26421_),
    .Z(_05655_));
 MUX2_X1 _58660_ (.A(lce_data_cmd_i[196]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [196]),
    .S(_26421_),
    .Z(_05656_));
 MUX2_X1 _58661_ (.A(lce_data_cmd_i[197]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [197]),
    .S(_26421_),
    .Z(_05657_));
 MUX2_X1 _58662_ (.A(lce_data_cmd_i[198]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [198]),
    .S(_26421_),
    .Z(_05658_));
 MUX2_X1 _58663_ (.A(lce_data_cmd_i[199]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [199]),
    .S(_26421_),
    .Z(_05659_));
 MUX2_X1 _58664_ (.A(lce_data_cmd_i[200]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [200]),
    .S(_26421_),
    .Z(_05662_));
 BUF_X16 _58665_ (.A(_26416_),
    .Z(_26422_));
 MUX2_X1 _58666_ (.A(lce_data_cmd_i[201]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [201]),
    .S(_26422_),
    .Z(_05663_));
 MUX2_X1 _58667_ (.A(lce_data_cmd_i[202]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [202]),
    .S(_26422_),
    .Z(_05664_));
 MUX2_X1 _58668_ (.A(lce_data_cmd_i[203]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [203]),
    .S(_26422_),
    .Z(_05665_));
 MUX2_X1 _58669_ (.A(lce_data_cmd_i[204]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [204]),
    .S(_26422_),
    .Z(_05666_));
 MUX2_X1 _58670_ (.A(lce_data_cmd_i[205]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [205]),
    .S(_26422_),
    .Z(_05667_));
 MUX2_X1 _58671_ (.A(lce_data_cmd_i[206]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [206]),
    .S(_26422_),
    .Z(_05668_));
 MUX2_X1 _58672_ (.A(lce_data_cmd_i[207]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [207]),
    .S(_26422_),
    .Z(_05669_));
 MUX2_X1 _58673_ (.A(lce_data_cmd_i[208]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [208]),
    .S(_26422_),
    .Z(_05670_));
 MUX2_X1 _58674_ (.A(lce_data_cmd_i[209]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [209]),
    .S(_26422_),
    .Z(_05671_));
 MUX2_X1 _58675_ (.A(lce_data_cmd_i[210]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [210]),
    .S(_26422_),
    .Z(_05673_));
 BUF_X8 _58676_ (.A(_26416_),
    .Z(_26423_));
 MUX2_X1 _58677_ (.A(lce_data_cmd_i[211]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [211]),
    .S(_26423_),
    .Z(_05674_));
 MUX2_X1 _58678_ (.A(lce_data_cmd_i[212]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [212]),
    .S(_26423_),
    .Z(_05675_));
 MUX2_X1 _58679_ (.A(lce_data_cmd_i[213]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [213]),
    .S(_26423_),
    .Z(_05676_));
 MUX2_X1 _58680_ (.A(lce_data_cmd_i[214]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [214]),
    .S(_26423_),
    .Z(_05677_));
 MUX2_X1 _58681_ (.A(lce_data_cmd_i[215]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [215]),
    .S(_26423_),
    .Z(_05678_));
 MUX2_X1 _58682_ (.A(lce_data_cmd_i[216]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [216]),
    .S(_26423_),
    .Z(_05679_));
 MUX2_X1 _58683_ (.A(lce_data_cmd_i[217]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [217]),
    .S(_26423_),
    .Z(_05680_));
 MUX2_X1 _58684_ (.A(lce_data_cmd_i[218]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [218]),
    .S(_26423_),
    .Z(_05681_));
 MUX2_X1 _58685_ (.A(lce_data_cmd_i[219]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [219]),
    .S(_26423_),
    .Z(_05682_));
 MUX2_X1 _58686_ (.A(lce_data_cmd_i[220]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [220]),
    .S(_26423_),
    .Z(_05684_));
 BUF_X16 _58687_ (.A(_26416_),
    .Z(_26424_));
 MUX2_X1 _58688_ (.A(lce_data_cmd_i[4]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [4]),
    .S(_26424_),
    .Z(_05994_));
 MUX2_X1 _58689_ (.A(lce_data_cmd_i[6]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [6]),
    .S(_26424_),
    .Z(_06214_));
 MUX2_X1 _58690_ (.A(lce_data_cmd_i[7]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [7]),
    .S(_26424_),
    .Z(_06325_));
 MUX2_X1 _58691_ (.A(lce_data_cmd_i[8]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [8]),
    .S(_26424_),
    .Z(_06436_));
 MUX2_X1 _58692_ (.A(lce_data_cmd_i[9]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [9]),
    .S(_26424_),
    .Z(_06547_));
 MUX2_X1 _58693_ (.A(lce_data_cmd_i[10]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [10]),
    .S(_26424_),
    .Z(_05561_));
 MUX2_X1 _58694_ (.A(lce_data_cmd_i[11]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [11]),
    .S(_26424_),
    .Z(_05572_));
 MUX2_X1 _58695_ (.A(lce_data_cmd_i[12]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [12]),
    .S(_26424_),
    .Z(_05583_));
 MUX2_X1 _58696_ (.A(lce_data_cmd_i[13]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [13]),
    .S(_26424_),
    .Z(_05594_));
 MUX2_X1 _58697_ (.A(lce_data_cmd_i[14]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [14]),
    .S(_26424_),
    .Z(_05605_));
 BUF_X8 _58698_ (.A(_26416_),
    .Z(_26425_));
 MUX2_X1 _58699_ (.A(lce_data_cmd_i[15]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [15]),
    .S(_26425_),
    .Z(_05616_));
 MUX2_X1 _58700_ (.A(lce_data_cmd_i[16]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [16]),
    .S(_26425_),
    .Z(_05627_));
 MUX2_X1 _58701_ (.A(lce_data_cmd_i[17]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [17]),
    .S(_26425_),
    .Z(_05638_));
 MUX2_X1 _58702_ (.A(lce_data_cmd_i[18]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [18]),
    .S(_26425_),
    .Z(_05649_));
 MUX2_X1 _58703_ (.A(lce_data_cmd_i[19]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [19]),
    .S(_26425_),
    .Z(_05660_));
 MUX2_X1 _58704_ (.A(lce_data_cmd_i[20]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [20]),
    .S(_26425_),
    .Z(_05672_));
 MUX2_X1 _58705_ (.A(lce_data_cmd_i[21]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [21]),
    .S(_26425_),
    .Z(_05683_));
 MUX2_X1 _58706_ (.A(lce_data_cmd_i[22]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [22]),
    .S(_26425_),
    .Z(_05694_));
 MUX2_X1 _58707_ (.A(lce_data_cmd_i[23]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [23]),
    .S(_26425_),
    .Z(_05705_));
 MUX2_X1 _58708_ (.A(lce_data_cmd_i[24]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [24]),
    .S(_26425_),
    .Z(_05716_));
 BUF_X16 _58709_ (.A(_26416_),
    .Z(_26426_));
 MUX2_X1 _58710_ (.A(lce_data_cmd_i[25]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [25]),
    .S(_26426_),
    .Z(_05727_));
 MUX2_X1 _58711_ (.A(lce_data_cmd_i[26]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [26]),
    .S(_26426_),
    .Z(_05738_));
 MUX2_X1 _58712_ (.A(lce_data_cmd_i[27]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [27]),
    .S(_26426_),
    .Z(_05749_));
 MUX2_X1 _58713_ (.A(lce_data_cmd_i[28]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [28]),
    .S(_26426_),
    .Z(_05760_));
 MUX2_X1 _58714_ (.A(lce_data_cmd_i[29]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [29]),
    .S(_26426_),
    .Z(_05771_));
 MUX2_X1 _58715_ (.A(lce_data_cmd_i[30]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [30]),
    .S(_26426_),
    .Z(_05783_));
 MUX2_X1 _58716_ (.A(lce_data_cmd_i[31]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [31]),
    .S(_26426_),
    .Z(_05794_));
 MUX2_X1 _58717_ (.A(lce_data_cmd_i[32]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [32]),
    .S(_26426_),
    .Z(_05805_));
 MUX2_X1 _58718_ (.A(lce_data_cmd_i[33]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [33]),
    .S(_26426_),
    .Z(_05816_));
 MUX2_X1 _58719_ (.A(lce_data_cmd_i[34]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [34]),
    .S(_26426_),
    .Z(_05827_));
 BUF_X16 _58720_ (.A(_26382_),
    .Z(_26427_));
 MUX2_X1 _58721_ (.A(lce_data_cmd_i[35]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [35]),
    .S(_26427_),
    .Z(_05838_));
 MUX2_X1 _58722_ (.A(lce_data_cmd_i[36]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [36]),
    .S(_26427_),
    .Z(_05849_));
 MUX2_X1 _58723_ (.A(lce_data_cmd_i[37]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [37]),
    .S(_26427_),
    .Z(_05860_));
 MUX2_X1 _58724_ (.A(lce_data_cmd_i[38]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [38]),
    .S(_26427_),
    .Z(_05871_));
 MUX2_X1 _58725_ (.A(lce_data_cmd_i[39]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [39]),
    .S(_26427_),
    .Z(_05882_));
 MUX2_X1 _58726_ (.A(lce_data_cmd_i[40]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [40]),
    .S(_26427_),
    .Z(_05894_));
 MUX2_X1 _58727_ (.A(lce_data_cmd_i[41]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [41]),
    .S(_26427_),
    .Z(_05905_));
 MUX2_X1 _58728_ (.A(lce_data_cmd_i[42]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [42]),
    .S(_26427_),
    .Z(_05916_));
 MUX2_X1 _58729_ (.A(lce_data_cmd_i[43]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [43]),
    .S(_26427_),
    .Z(_05927_));
 MUX2_X1 _58730_ (.A(lce_data_cmd_i[44]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [44]),
    .S(_26427_),
    .Z(_05938_));
 BUF_X8 _58731_ (.A(_26382_),
    .Z(_26428_));
 MUX2_X1 _58732_ (.A(lce_data_cmd_i[45]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [45]),
    .S(_26428_),
    .Z(_05949_));
 MUX2_X1 _58733_ (.A(lce_data_cmd_i[46]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [46]),
    .S(_26428_),
    .Z(_05960_));
 MUX2_X1 _58734_ (.A(lce_data_cmd_i[47]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [47]),
    .S(_26428_),
    .Z(_05971_));
 MUX2_X1 _58735_ (.A(lce_data_cmd_i[48]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [48]),
    .S(_26428_),
    .Z(_05982_));
 MUX2_X1 _58736_ (.A(lce_data_cmd_i[49]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [49]),
    .S(_26428_),
    .Z(_05993_));
 MUX2_X1 _58737_ (.A(lce_data_cmd_i[50]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [50]),
    .S(_26428_),
    .Z(_06005_));
 MUX2_X1 _58738_ (.A(lce_data_cmd_i[51]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [51]),
    .S(_26428_),
    .Z(_06016_));
 MUX2_X1 _58739_ (.A(lce_data_cmd_i[52]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [52]),
    .S(_26428_),
    .Z(_06026_));
 MUX2_X1 _58740_ (.A(lce_data_cmd_i[53]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [53]),
    .S(_26428_),
    .Z(_06037_));
 MUX2_X1 _58741_ (.A(lce_data_cmd_i[54]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [54]),
    .S(_26428_),
    .Z(_06048_));
 BUF_X8 _58742_ (.A(_26382_),
    .Z(_26429_));
 MUX2_X1 _58743_ (.A(lce_data_cmd_i[55]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [55]),
    .S(_26429_),
    .Z(_06059_));
 MUX2_X1 _58744_ (.A(lce_data_cmd_i[56]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [56]),
    .S(_26429_),
    .Z(_06070_));
 MUX2_X1 _58745_ (.A(lce_data_cmd_i[57]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [57]),
    .S(_26429_),
    .Z(_06081_));
 MUX2_X1 _58746_ (.A(lce_data_cmd_i[58]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [58]),
    .S(_26429_),
    .Z(_06092_));
 MUX2_X1 _58747_ (.A(lce_data_cmd_i[59]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [59]),
    .S(_26429_),
    .Z(_06103_));
 MUX2_X1 _58748_ (.A(lce_data_cmd_i[60]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [60]),
    .S(_26429_),
    .Z(_06114_));
 MUX2_X1 _58749_ (.A(lce_data_cmd_i[61]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [61]),
    .S(_26429_),
    .Z(_06125_));
 MUX2_X1 _58750_ (.A(lce_data_cmd_i[62]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [62]),
    .S(_26429_),
    .Z(_06136_));
 MUX2_X1 _58751_ (.A(lce_data_cmd_i[63]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [63]),
    .S(_26429_),
    .Z(_06147_));
 MUX2_X1 _58752_ (.A(lce_data_cmd_i[64]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [64]),
    .S(_26429_),
    .Z(_06158_));
 BUF_X16 _58753_ (.A(_26382_),
    .Z(_26430_));
 MUX2_X1 _58754_ (.A(lce_data_cmd_i[65]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [65]),
    .S(_26430_),
    .Z(_06169_));
 MUX2_X1 _58755_ (.A(lce_data_cmd_i[66]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [66]),
    .S(_26430_),
    .Z(_06180_));
 MUX2_X1 _58756_ (.A(lce_data_cmd_i[67]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [67]),
    .S(_26430_),
    .Z(_06191_));
 MUX2_X1 _58757_ (.A(lce_data_cmd_i[68]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [68]),
    .S(_26430_),
    .Z(_06202_));
 MUX2_X1 _58758_ (.A(lce_data_cmd_i[69]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [69]),
    .S(_26430_),
    .Z(_06213_));
 MUX2_X1 _58759_ (.A(lce_data_cmd_i[70]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [70]),
    .S(_26430_),
    .Z(_06225_));
 MUX2_X1 _58760_ (.A(lce_data_cmd_i[71]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [71]),
    .S(_26430_),
    .Z(_06236_));
 MUX2_X1 _58761_ (.A(lce_data_cmd_i[72]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [72]),
    .S(_26430_),
    .Z(_06247_));
 MUX2_X1 _58762_ (.A(lce_data_cmd_i[73]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [73]),
    .S(_26430_),
    .Z(_06258_));
 MUX2_X1 _58763_ (.A(lce_data_cmd_i[74]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [74]),
    .S(_26430_),
    .Z(_06269_));
 BUF_X16 _58764_ (.A(_26382_),
    .Z(_26431_));
 MUX2_X1 _58765_ (.A(lce_data_cmd_i[75]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [75]),
    .S(_26431_),
    .Z(_06280_));
 MUX2_X1 _58766_ (.A(lce_data_cmd_i[76]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [76]),
    .S(_26431_),
    .Z(_06291_));
 MUX2_X1 _58767_ (.A(lce_data_cmd_i[77]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [77]),
    .S(_26431_),
    .Z(_06302_));
 MUX2_X1 _58768_ (.A(lce_data_cmd_i[78]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [78]),
    .S(_26431_),
    .Z(_06313_));
 MUX2_X1 _58769_ (.A(lce_data_cmd_i[79]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [79]),
    .S(_26431_),
    .Z(_06324_));
 MUX2_X1 _58770_ (.A(lce_data_cmd_i[80]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [80]),
    .S(_26431_),
    .Z(_06336_));
 MUX2_X1 _58771_ (.A(lce_data_cmd_i[81]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [81]),
    .S(_26431_),
    .Z(_06347_));
 MUX2_X1 _58772_ (.A(lce_data_cmd_i[82]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [82]),
    .S(_26431_),
    .Z(_06358_));
 MUX2_X1 _58773_ (.A(lce_data_cmd_i[83]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [83]),
    .S(_26431_),
    .Z(_06369_));
 MUX2_X1 _58774_ (.A(lce_data_cmd_i[84]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [84]),
    .S(_26431_),
    .Z(_06380_));
 BUF_X8 _58775_ (.A(_26382_),
    .Z(_26432_));
 MUX2_X1 _58776_ (.A(lce_data_cmd_i[85]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [85]),
    .S(_26432_),
    .Z(_06391_));
 MUX2_X1 _58777_ (.A(lce_data_cmd_i[86]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [86]),
    .S(_26432_),
    .Z(_06402_));
 MUX2_X1 _58778_ (.A(lce_data_cmd_i[87]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [87]),
    .S(_26432_),
    .Z(_06413_));
 MUX2_X1 _58779_ (.A(lce_data_cmd_i[88]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [88]),
    .S(_26432_),
    .Z(_06424_));
 MUX2_X1 _58780_ (.A(lce_data_cmd_i[89]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [89]),
    .S(_26432_),
    .Z(_06435_));
 MUX2_X1 _58781_ (.A(lce_data_cmd_i[90]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [90]),
    .S(_26432_),
    .Z(_06447_));
 MUX2_X1 _58782_ (.A(lce_data_cmd_i[91]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [91]),
    .S(_26432_),
    .Z(_06458_));
 MUX2_X1 _58783_ (.A(lce_data_cmd_i[92]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [92]),
    .S(_26432_),
    .Z(_06469_));
 MUX2_X1 _58784_ (.A(lce_data_cmd_i[93]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [93]),
    .S(_26432_),
    .Z(_06480_));
 MUX2_X1 _58785_ (.A(lce_data_cmd_i[94]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [94]),
    .S(_26432_),
    .Z(_06491_));
 BUF_X8 _58786_ (.A(_26382_),
    .Z(_26433_));
 MUX2_X1 _58787_ (.A(lce_data_cmd_i[95]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [95]),
    .S(_26433_),
    .Z(_06502_));
 MUX2_X1 _58788_ (.A(lce_data_cmd_i[96]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [96]),
    .S(_26433_),
    .Z(_06513_));
 MUX2_X1 _58789_ (.A(lce_data_cmd_i[97]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [97]),
    .S(_26433_),
    .Z(_06524_));
 MUX2_X1 _58790_ (.A(lce_data_cmd_i[98]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [98]),
    .S(_26433_),
    .Z(_06535_));
 MUX2_X1 _58791_ (.A(lce_data_cmd_i[99]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [99]),
    .S(_26433_),
    .Z(_06546_));
 MUX2_X1 _58792_ (.A(lce_data_cmd_i[100]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [100]),
    .S(_26433_),
    .Z(_05525_));
 MUX2_X1 _58793_ (.A(lce_data_cmd_i[101]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [101]),
    .S(_26433_),
    .Z(_05536_));
 MUX2_X1 _58794_ (.A(lce_data_cmd_i[102]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [102]),
    .S(_26433_),
    .Z(_05547_));
 MUX2_X1 _58795_ (.A(lce_data_cmd_i[103]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [103]),
    .S(_26433_),
    .Z(_05554_));
 MUX2_X1 _58796_ (.A(lce_data_cmd_i[104]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [104]),
    .S(_26433_),
    .Z(_05555_));
 BUF_X8 _58797_ (.A(_26382_),
    .Z(_26434_));
 MUX2_X1 _58798_ (.A(lce_data_cmd_i[105]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [105]),
    .S(_26434_),
    .Z(_05556_));
 MUX2_X1 _58799_ (.A(lce_data_cmd_i[106]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [106]),
    .S(_26434_),
    .Z(_05557_));
 MUX2_X1 _58800_ (.A(lce_data_cmd_i[107]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [107]),
    .S(_26434_),
    .Z(_05558_));
 MUX2_X1 _58801_ (.A(lce_data_cmd_i[108]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [108]),
    .S(_26434_),
    .Z(_05559_));
 MUX2_X1 _58802_ (.A(lce_data_cmd_i[109]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [109]),
    .S(_26434_),
    .Z(_05560_));
 MUX2_X1 _58803_ (.A(lce_data_cmd_i[110]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [110]),
    .S(_26434_),
    .Z(_05562_));
 MUX2_X1 _58804_ (.A(lce_data_cmd_i[111]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [111]),
    .S(_26434_),
    .Z(_05563_));
 MUX2_X1 _58805_ (.A(lce_data_cmd_i[112]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [112]),
    .S(_26434_),
    .Z(_05564_));
 MUX2_X1 _58806_ (.A(lce_data_cmd_i[113]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [113]),
    .S(_26434_),
    .Z(_05565_));
 MUX2_X1 _58807_ (.A(lce_data_cmd_i[114]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [114]),
    .S(_26434_),
    .Z(_05566_));
 MUX2_X1 _58808_ (.A(lce_data_cmd_i[115]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [115]),
    .S(_26378_),
    .Z(_05567_));
 MUX2_X1 _58809_ (.A(lce_data_cmd_i[116]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [116]),
    .S(_26378_),
    .Z(_05568_));
 MUX2_X1 _58810_ (.A(lce_data_cmd_i[117]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [117]),
    .S(_26378_),
    .Z(_05569_));
 MUX2_X1 _58811_ (.A(lce_data_cmd_i[118]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [118]),
    .S(_26378_),
    .Z(_05570_));
 MUX2_X1 _58812_ (.A(lce_data_cmd_i[119]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [119]),
    .S(_26378_),
    .Z(_05571_));
 MUX2_X1 _58813_ (.A(lce_data_cmd_i[120]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [120]),
    .S(_26378_),
    .Z(_05573_));
 MUX2_X1 _58814_ (.A(lce_data_cmd_i[121]),
    .B(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [121]),
    .S(_26378_),
    .Z(_05574_));
 AND4_X1 _58815_ (.A1(fe_cmd_v_i),
    .A2(_08028_),
    .A3(_21337_),
    .A4(_08662_),
    .ZN(N8));
 BUF_X8 _58816_ (.A(_08518_),
    .Z(_26435_));
 MUX2_X1 _58817_ (.A(\bp_fe_pc_gen_1.icache_pc_gen_i [0]),
    .B(\icache.vaddr_tl_r [0]),
    .S(_26435_),
    .Z(_03997_));
 MUX2_X1 _58818_ (.A(\bp_fe_pc_gen_1.icache_pc_gen_i [1]),
    .B(\icache.vaddr_tl_r [1]),
    .S(_26435_),
    .Z(_04008_));
 BUF_X8 _58819_ (.A(_08518_),
    .Z(_26436_));
 NAND2_X2 _58820_ (.A1(_26436_),
    .A2(\icache.vaddr_tl_r [2]),
    .ZN(_26437_));
 OAI21_X1 _58821_ (.A(_26437_),
    .B1(_11222_),
    .B2(\icache.N29 ),
    .ZN(_04019_));
 MUX2_X1 _58822_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [12]),
    .B(\icache.vaddr_tl_r [3]),
    .S(_26435_),
    .Z(_04029_));
 MUX2_X1 _58823_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [13]),
    .B(\icache.vaddr_tl_r [4]),
    .S(_26435_),
    .Z(_04030_));
 NAND2_X1 _58824_ (.A1(_26436_),
    .A2(\icache.vaddr_tl_r [5]),
    .ZN(_26438_));
 OAI21_X1 _58825_ (.A(_26438_),
    .B1(_11226_),
    .B2(\icache.N29 ),
    .ZN(_04031_));
 NAND2_X1 _58826_ (.A1(_26436_),
    .A2(\icache.vaddr_tl_r [6]),
    .ZN(_26439_));
 OAI21_X1 _58827_ (.A(_26439_),
    .B1(_11227_),
    .B2(\icache.N29 ),
    .ZN(_04032_));
 NAND2_X1 _58828_ (.A1(_26435_),
    .A2(\icache.vaddr_tl_r [7]),
    .ZN(_26440_));
 OAI21_X1 _58829_ (.A(_26440_),
    .B1(_11228_),
    .B2(\icache.N29 ),
    .ZN(_04033_));
 NAND2_X1 _58830_ (.A1(_26435_),
    .A2(\icache.vaddr_tl_r [8]),
    .ZN(_26441_));
 OAI21_X1 _58831_ (.A(_26441_),
    .B1(_11229_),
    .B2(\icache.N29 ),
    .ZN(_04034_));
 NAND2_X1 _58832_ (.A1(_26435_),
    .A2(\icache.vaddr_tl_r [9]),
    .ZN(_26442_));
 OAI21_X1 _58833_ (.A(_26442_),
    .B1(_11230_),
    .B2(\icache.N29 ),
    .ZN(_04035_));
 NAND2_X2 _58834_ (.A1(_26435_),
    .A2(\icache.vaddr_tl_r [10]),
    .ZN(_26443_));
 OAI21_X1 _58835_ (.A(_26443_),
    .B1(_11231_),
    .B2(\icache.N29 ),
    .ZN(_03998_));
 NAND2_X2 _58836_ (.A1(_26435_),
    .A2(\icache.vaddr_tl_r [11]),
    .ZN(_26444_));
 OAI21_X1 _58837_ (.A(_26444_),
    .B1(_11232_),
    .B2(\icache.N29 ),
    .ZN(_03999_));
 MUX2_X1 _58838_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [21]),
    .B(\icache.vaddr_tl_r [12]),
    .S(_26435_),
    .Z(_04000_));
 BUF_X8 _58839_ (.A(_08518_),
    .Z(_26445_));
 MUX2_X1 _58840_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [22]),
    .B(\icache.vaddr_tl_r [13]),
    .S(_26445_),
    .Z(_04001_));
 MUX2_X1 _58841_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [23]),
    .B(\icache.vaddr_tl_r [14]),
    .S(_26445_),
    .Z(_04002_));
 MUX2_X1 _58842_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [24]),
    .B(\icache.vaddr_tl_r [15]),
    .S(_26445_),
    .Z(_04003_));
 MUX2_X1 _58843_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [25]),
    .B(\icache.vaddr_tl_r [16]),
    .S(_26445_),
    .Z(_04004_));
 MUX2_X1 _58844_ (.A(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [26]),
    .B(\icache.vaddr_tl_r [17]),
    .S(_26445_),
    .Z(_04005_));
 MUX2_X1 _58845_ (.A(\bp_fe_pc_gen_1.icache_pc_gen_i [18]),
    .B(\icache.vaddr_tl_r [18]),
    .S(_26445_),
    .Z(_04006_));
 MUX2_X1 _58846_ (.A(\bp_fe_pc_gen_1.icache_pc_gen_i [19]),
    .B(\icache.vaddr_tl_r [19]),
    .S(_26445_),
    .Z(_04007_));
 MUX2_X1 _58847_ (.A(\bp_fe_pc_gen_1.icache_pc_gen_i [20]),
    .B(\icache.vaddr_tl_r [20]),
    .S(_26445_),
    .Z(_04009_));
 MUX2_X1 _58848_ (.A(\bp_fe_pc_gen_1.icache_pc_gen_i [21]),
    .B(\icache.vaddr_tl_r [21]),
    .S(_26445_),
    .Z(_04010_));
 MUX2_X1 _58849_ (.A(\bp_fe_pc_gen_1.icache_pc_gen_i [22]),
    .B(\icache.vaddr_tl_r [22]),
    .S(_26445_),
    .Z(_04011_));
 BUF_X8 _58850_ (.A(_08518_),
    .Z(_26446_));
 MUX2_X1 _58851_ (.A(\bp_fe_pc_gen_1.icache_pc_gen_i [23]),
    .B(\icache.vaddr_tl_r [23]),
    .S(_26446_),
    .Z(_04012_));
 MUX2_X1 _58852_ (.A(\bp_fe_pc_gen_1.icache_pc_gen_i [24]),
    .B(\icache.vaddr_tl_r [24]),
    .S(_26446_),
    .Z(_04013_));
 MUX2_X1 _58853_ (.A(\bp_fe_pc_gen_1.icache_pc_gen_i [25]),
    .B(\icache.vaddr_tl_r [25]),
    .S(_26446_),
    .Z(_04014_));
 MUX2_X1 _58854_ (.A(\bp_fe_pc_gen_1.icache_pc_gen_i [26]),
    .B(\icache.vaddr_tl_r [26]),
    .S(_26446_),
    .Z(_04015_));
 MUX2_X1 _58855_ (.A(\bp_fe_pc_gen_1.icache_pc_gen_i [27]),
    .B(\icache.vaddr_tl_r [27]),
    .S(_26446_),
    .Z(_04016_));
 MUX2_X1 _58856_ (.A(\bp_fe_pc_gen_1.icache_pc_gen_i [28]),
    .B(\icache.vaddr_tl_r [28]),
    .S(_26446_),
    .Z(_04017_));
 MUX2_X1 _58857_ (.A(\bp_fe_pc_gen_1.icache_pc_gen_i [29]),
    .B(\icache.vaddr_tl_r [29]),
    .S(_26446_),
    .Z(_04018_));
 MUX2_X1 _58858_ (.A(\bp_fe_pc_gen_1.icache_pc_gen_i [30]),
    .B(\icache.vaddr_tl_r [30]),
    .S(_26446_),
    .Z(_04020_));
 MUX2_X1 _58859_ (.A(\bp_fe_pc_gen_1.icache_pc_gen_i [31]),
    .B(\icache.vaddr_tl_r [31]),
    .S(_26446_),
    .Z(_04021_));
 MUX2_X1 _58860_ (.A(\bp_fe_pc_gen_1.icache_pc_gen_i [32]),
    .B(\icache.vaddr_tl_r [32]),
    .S(_26446_),
    .Z(_04022_));
 BUF_X16 _58861_ (.A(_08518_),
    .Z(_26447_));
 MUX2_X1 _58862_ (.A(\bp_fe_pc_gen_1.icache_pc_gen_i [33]),
    .B(\icache.vaddr_tl_r [33]),
    .S(_26447_),
    .Z(_04023_));
 MUX2_X1 _58863_ (.A(\bp_fe_pc_gen_1.icache_pc_gen_i [34]),
    .B(\icache.vaddr_tl_r [34]),
    .S(_26447_),
    .Z(_04024_));
 MUX2_X1 _58864_ (.A(\bp_fe_pc_gen_1.icache_pc_gen_i [35]),
    .B(\icache.vaddr_tl_r [35]),
    .S(_26447_),
    .Z(_04025_));
 MUX2_X1 _58865_ (.A(\bp_fe_pc_gen_1.icache_pc_gen_i [36]),
    .B(\icache.vaddr_tl_r [36]),
    .S(_26447_),
    .Z(_04026_));
 MUX2_X1 _58866_ (.A(\bp_fe_pc_gen_1.icache_pc_gen_i [37]),
    .B(\icache.vaddr_tl_r [37]),
    .S(_26447_),
    .Z(_04027_));
 MUX2_X1 _58867_ (.A(\bp_fe_pc_gen_1.icache_pc_gen_i [38]),
    .B(\icache.vaddr_tl_r [38]),
    .S(_26447_),
    .Z(_04028_));
 AOI21_X1 _58868_ (.A(\icache.vaddr_tl_r [0]),
    .B1(_08037_),
    .B2(_08727_),
    .ZN(_26448_));
 AOI21_X1 _58869_ (.A(_26448_),
    .B1(_08738_),
    .B2(\icache.N25 ),
    .ZN(_04849_));
 NAND3_X1 _58870_ (.A1(_08740_),
    .A2(\icache.N25 ),
    .A3(_08741_),
    .ZN(_26449_));
 OR2_X1 _58871_ (.A1(_08521_),
    .A2(\icache.vaddr_tl_r [1]),
    .ZN(_26450_));
 AND2_X1 _58872_ (.A1(_26449_),
    .A2(_26450_),
    .ZN(_04860_));
 OAI21_X1 _58873_ (.A(\icache.vaddr_tl_r [2]),
    .B1(_08481_),
    .B2(_21279_),
    .ZN(_26451_));
 BUF_X4 _58874_ (.A(_10634_),
    .Z(_26452_));
 OAI21_X1 _58875_ (.A(_26451_),
    .B1(_11215_),
    .B2(_26452_),
    .ZN(_04871_));
 OAI21_X1 _58876_ (.A(\icache.vaddr_tl_r [3]),
    .B1(_08481_),
    .B2(_21279_),
    .ZN(_26453_));
 OAI21_X1 _58877_ (.A(_26453_),
    .B1(_08752_),
    .B2(_26452_),
    .ZN(_04881_));
 OAI21_X1 _58878_ (.A(\icache.vaddr_tl_r [4]),
    .B1(_08481_),
    .B2(_21279_),
    .ZN(_26454_));
 OAI21_X1 _58879_ (.A(_26454_),
    .B1(_08755_),
    .B2(_26452_),
    .ZN(_04882_));
 OAI21_X1 _58880_ (.A(\icache.vaddr_tl_r [5]),
    .B1(_08481_),
    .B2(_21279_),
    .ZN(_26455_));
 OAI21_X1 _58881_ (.A(_26455_),
    .B1(_08757_),
    .B2(_26452_),
    .ZN(_04883_));
 OAI21_X1 _58882_ (.A(\icache.vaddr_tl_r [6]),
    .B1(_08481_),
    .B2(_21279_),
    .ZN(_26456_));
 OAI21_X1 _58883_ (.A(_26456_),
    .B1(_08759_),
    .B2(_26452_),
    .ZN(_04884_));
 OAI21_X1 _58884_ (.A(\icache.vaddr_tl_r [7]),
    .B1(_08481_),
    .B2(_21279_),
    .ZN(_26457_));
 OAI21_X1 _58885_ (.A(_26457_),
    .B1(_08762_),
    .B2(_26452_),
    .ZN(_04885_));
 BUF_X8 _58886_ (.A(_08480_),
    .Z(_26458_));
 OAI21_X1 _58887_ (.A(\icache.vaddr_tl_r [8]),
    .B1(_26458_),
    .B2(_21279_),
    .ZN(_26459_));
 OAI21_X1 _58888_ (.A(_26459_),
    .B1(_08764_),
    .B2(_26452_),
    .ZN(_04886_));
 OAI21_X1 _58889_ (.A(\icache.vaddr_tl_r [9]),
    .B1(_26458_),
    .B2(_21279_),
    .ZN(_26460_));
 OAI21_X1 _58890_ (.A(_26460_),
    .B1(_11216_),
    .B2(_26452_),
    .ZN(_04887_));
 OAI21_X1 _58891_ (.A(\icache.vaddr_tl_r [10]),
    .B1(_26458_),
    .B2(_08998_),
    .ZN(_26461_));
 OAI21_X1 _58892_ (.A(_26461_),
    .B1(_08767_),
    .B2(_26452_),
    .ZN(_04850_));
 OAI21_X1 _58893_ (.A(\icache.vaddr_tl_r [11]),
    .B1(_26458_),
    .B2(_08998_),
    .ZN(_26462_));
 OAI21_X1 _58894_ (.A(_26462_),
    .B1(_08769_),
    .B2(_26452_),
    .ZN(_04851_));
 MUX2_X1 _58895_ (.A(\icache.vaddr_tl_r [12]),
    .B(_10233_),
    .S(\icache.N25 ),
    .Z(_04852_));
 OAI21_X1 _58896_ (.A(\icache.vaddr_tl_r [13]),
    .B1(_26458_),
    .B2(_08998_),
    .ZN(_26463_));
 OAI21_X1 _58897_ (.A(_26463_),
    .B1(_10077_),
    .B2(_10634_),
    .ZN(_04853_));
 OAI21_X1 _58898_ (.A(\icache.vaddr_tl_r [14]),
    .B1(_26458_),
    .B2(_08998_),
    .ZN(_26464_));
 OAI21_X1 _58899_ (.A(_26464_),
    .B1(_08805_),
    .B2(_10634_),
    .ZN(_04854_));
 MUX2_X1 _58900_ (.A(\icache.vaddr_tl_r [15]),
    .B(_10171_),
    .S(\icache.N25 ),
    .Z(_04855_));
 MUX2_X1 _58901_ (.A(\icache.vaddr_tl_r [16]),
    .B(_10330_),
    .S(\icache.N25 ),
    .Z(_04856_));
 OAI21_X1 _58902_ (.A(\icache.vaddr_tl_r [17]),
    .B1(_26458_),
    .B2(_08998_),
    .ZN(_26465_));
 OAI21_X1 _58903_ (.A(_26465_),
    .B1(_10100_),
    .B2(_10634_),
    .ZN(_04857_));
 MUX2_X1 _58904_ (.A(\icache.vaddr_tl_r [18]),
    .B(_10449_),
    .S(\icache.N25 ),
    .Z(_04858_));
 OAI21_X1 _58905_ (.A(\icache.vaddr_tl_r [19]),
    .B1(_26458_),
    .B2(_08998_),
    .ZN(_26466_));
 OAI21_X1 _58906_ (.A(_26466_),
    .B1(_10101_),
    .B2(_10634_),
    .ZN(_04859_));
 OAI21_X1 _58907_ (.A(\icache.vaddr_tl_r [20]),
    .B1(_26458_),
    .B2(_08998_),
    .ZN(_26467_));
 OAI21_X1 _58908_ (.A(_26467_),
    .B1(_08853_),
    .B2(_10634_),
    .ZN(_04861_));
 MUX2_X1 _58909_ (.A(\icache.vaddr_tl_r [21]),
    .B(_10037_),
    .S(\icache.N25 ),
    .Z(_04862_));
 MUX2_X1 _58910_ (.A(\icache.vaddr_tl_r [22]),
    .B(_10088_),
    .S(\icache.N25 ),
    .Z(_04863_));
 AOI21_X1 _58911_ (.A(\icache.vaddr_tl_r [23]),
    .B1(_08037_),
    .B2(_08674_),
    .ZN(_26468_));
 AOI21_X1 _58912_ (.A(_26468_),
    .B1(_10064_),
    .B2(\icache.N25 ),
    .ZN(_04864_));
 BUF_X8 _58913_ (.A(_08521_),
    .Z(_26469_));
 MUX2_X1 _58914_ (.A(\icache.vaddr_tl_r [24]),
    .B(_10455_),
    .S(_26469_),
    .Z(_04865_));
 MUX2_X1 _58915_ (.A(\icache.vaddr_tl_r [25]),
    .B(_10283_),
    .S(_26469_),
    .Z(_04866_));
 OAI21_X1 _58916_ (.A(\icache.vaddr_tl_r [26]),
    .B1(_26458_),
    .B2(_08998_),
    .ZN(_26470_));
 OAI21_X1 _58917_ (.A(_26470_),
    .B1(_08901_),
    .B2(_10634_),
    .ZN(_04867_));
 MUX2_X1 _58918_ (.A(\icache.vaddr_tl_r [27]),
    .B(_10350_),
    .S(_26469_),
    .Z(_04868_));
 MUX2_X1 _58919_ (.A(\icache.vaddr_tl_r [28]),
    .B(_10106_),
    .S(_26469_),
    .Z(_04869_));
 MUX2_X1 _58920_ (.A(\icache.vaddr_tl_r [29]),
    .B(_10162_),
    .S(_26469_),
    .Z(_04870_));
 MUX2_X1 _58921_ (.A(\icache.vaddr_tl_r [30]),
    .B(_10193_),
    .S(_26469_),
    .Z(_04872_));
 MUX2_X1 _58922_ (.A(\icache.vaddr_tl_r [31]),
    .B(_10043_),
    .S(_26469_),
    .Z(_04873_));
 MUX2_X1 _58923_ (.A(\icache.vaddr_tl_r [32]),
    .B(_10123_),
    .S(_26469_),
    .Z(_04874_));
 MUX2_X1 _58924_ (.A(\icache.vaddr_tl_r [33]),
    .B(_10164_),
    .S(_26469_),
    .Z(_04875_));
 MUX2_X1 _58925_ (.A(\icache.vaddr_tl_r [34]),
    .B(_10381_),
    .S(_26469_),
    .Z(_04876_));
 MUX2_X1 _58926_ (.A(\icache.vaddr_tl_r [35]),
    .B(_10326_),
    .S(_08521_),
    .Z(_04877_));
 MUX2_X1 _58927_ (.A(\icache.vaddr_tl_r [36]),
    .B(_10117_),
    .S(_08521_),
    .Z(_04878_));
 MUX2_X1 _58928_ (.A(\icache.vaddr_tl_r [37]),
    .B(_10179_),
    .S(_08521_),
    .Z(_04879_));
 MUX2_X1 _58929_ (.A(\icache.vaddr_tl_r [38]),
    .B(_10268_),
    .S(_08521_),
    .Z(_04880_));
 MUX2_X1 _58930_ (.A(\icache.data_set_select_mux.data_i [414]),
    .B(\icache.data_mems_6__data_mem.data_o [30]),
    .S(_26447_),
    .Z(_04388_));
 MUX2_X1 _58931_ (.A(\icache.data_set_select_mux.data_i [415]),
    .B(\icache.data_mems_6__data_mem.data_o [31]),
    .S(_26447_),
    .Z(_04389_));
 MUX2_X1 _58932_ (.A(\icache.data_set_select_mux.data_i [416]),
    .B(\icache.data_mems_6__data_mem.data_o [32]),
    .S(_26447_),
    .Z(_04390_));
 MUX2_X1 _58933_ (.A(\icache.data_set_select_mux.data_i [417]),
    .B(\icache.data_mems_6__data_mem.data_o [33]),
    .S(_26447_),
    .Z(_04391_));
 BUF_X4 _58934_ (.A(_08518_),
    .Z(_26471_));
 MUX2_X1 _58935_ (.A(\icache.data_set_select_mux.data_i [418]),
    .B(\icache.data_mems_6__data_mem.data_o [34]),
    .S(_26471_),
    .Z(_04392_));
 MUX2_X1 _58936_ (.A(\icache.data_set_select_mux.data_i [419]),
    .B(\icache.data_mems_6__data_mem.data_o [35]),
    .S(_26471_),
    .Z(_04393_));
 MUX2_X1 _58937_ (.A(\icache.data_set_select_mux.data_i [420]),
    .B(\icache.data_mems_6__data_mem.data_o [36]),
    .S(_26471_),
    .Z(_04395_));
 MUX2_X1 _58938_ (.A(\icache.data_set_select_mux.data_i [421]),
    .B(\icache.data_mems_6__data_mem.data_o [37]),
    .S(_26471_),
    .Z(_04396_));
 MUX2_X1 _58939_ (.A(\icache.data_set_select_mux.data_i [422]),
    .B(\icache.data_mems_6__data_mem.data_o [38]),
    .S(_26471_),
    .Z(_04397_));
 MUX2_X1 _58940_ (.A(\icache.data_set_select_mux.data_i [423]),
    .B(\icache.data_mems_6__data_mem.data_o [39]),
    .S(_26471_),
    .Z(_04398_));
 MUX2_X1 _58941_ (.A(\icache.data_set_select_mux.data_i [424]),
    .B(\icache.data_mems_6__data_mem.data_o [40]),
    .S(_26471_),
    .Z(_04399_));
 MUX2_X1 _58942_ (.A(\icache.data_set_select_mux.data_i [425]),
    .B(\icache.data_mems_6__data_mem.data_o [41]),
    .S(_26471_),
    .Z(_04400_));
 MUX2_X1 _58943_ (.A(\icache.data_set_select_mux.data_i [426]),
    .B(\icache.data_mems_6__data_mem.data_o [42]),
    .S(_26471_),
    .Z(_04401_));
 MUX2_X1 _58944_ (.A(\icache.data_set_select_mux.data_i [427]),
    .B(\icache.data_mems_6__data_mem.data_o [43]),
    .S(_26471_),
    .Z(_04402_));
 BUF_X8 _58945_ (.A(_08518_),
    .Z(_26472_));
 MUX2_X1 _58946_ (.A(\icache.data_set_select_mux.data_i [428]),
    .B(\icache.data_mems_6__data_mem.data_o [44]),
    .S(_26472_),
    .Z(_04403_));
 MUX2_X1 _58947_ (.A(\icache.data_set_select_mux.data_i [429]),
    .B(\icache.data_mems_6__data_mem.data_o [45]),
    .S(_26472_),
    .Z(_04404_));
 MUX2_X1 _58948_ (.A(\icache.data_set_select_mux.data_i [430]),
    .B(\icache.data_mems_6__data_mem.data_o [46]),
    .S(_26472_),
    .Z(_04406_));
 MUX2_X1 _58949_ (.A(\icache.data_set_select_mux.data_i [431]),
    .B(\icache.data_mems_6__data_mem.data_o [47]),
    .S(_26472_),
    .Z(_04407_));
 MUX2_X1 _58950_ (.A(\icache.data_set_select_mux.data_i [432]),
    .B(\icache.data_mems_6__data_mem.data_o [48]),
    .S(_26472_),
    .Z(_04408_));
 MUX2_X1 _58951_ (.A(\icache.data_set_select_mux.data_i [433]),
    .B(\icache.data_mems_6__data_mem.data_o [49]),
    .S(_26472_),
    .Z(_04409_));
 MUX2_X1 _58952_ (.A(\icache.data_set_select_mux.data_i [434]),
    .B(\icache.data_mems_6__data_mem.data_o [50]),
    .S(_26472_),
    .Z(_04410_));
 MUX2_X1 _58953_ (.A(\icache.data_set_select_mux.data_i [435]),
    .B(\icache.data_mems_6__data_mem.data_o [51]),
    .S(_26472_),
    .Z(_04411_));
 MUX2_X1 _58954_ (.A(\icache.data_set_select_mux.data_i [436]),
    .B(\icache.data_mems_6__data_mem.data_o [52]),
    .S(_26472_),
    .Z(_04412_));
 MUX2_X1 _58955_ (.A(\icache.data_set_select_mux.data_i [437]),
    .B(\icache.data_mems_6__data_mem.data_o [53]),
    .S(_26472_),
    .Z(_04413_));
 BUF_X32 _58956_ (.A(_08517_),
    .Z(_26473_));
 BUF_X16 _58957_ (.A(_26473_),
    .Z(_26474_));
 BUF_X8 _58958_ (.A(_26474_),
    .Z(_26475_));
 MUX2_X1 _58959_ (.A(\icache.data_set_select_mux.data_i [438]),
    .B(\icache.data_mems_6__data_mem.data_o [54]),
    .S(_26475_),
    .Z(_04414_));
 MUX2_X1 _58960_ (.A(\icache.data_set_select_mux.data_i [439]),
    .B(\icache.data_mems_6__data_mem.data_o [55]),
    .S(_26475_),
    .Z(_04415_));
 MUX2_X1 _58961_ (.A(\icache.data_set_select_mux.data_i [440]),
    .B(\icache.data_mems_6__data_mem.data_o [56]),
    .S(_26475_),
    .Z(_04417_));
 MUX2_X1 _58962_ (.A(\icache.data_set_select_mux.data_i [441]),
    .B(\icache.data_mems_6__data_mem.data_o [57]),
    .S(_26475_),
    .Z(_04418_));
 MUX2_X1 _58963_ (.A(\icache.data_set_select_mux.data_i [442]),
    .B(\icache.data_mems_6__data_mem.data_o [58]),
    .S(_26475_),
    .Z(_04419_));
 MUX2_X1 _58964_ (.A(\icache.data_set_select_mux.data_i [443]),
    .B(\icache.data_mems_6__data_mem.data_o [59]),
    .S(_26475_),
    .Z(_04420_));
 MUX2_X1 _58965_ (.A(\icache.data_set_select_mux.data_i [444]),
    .B(\icache.data_mems_6__data_mem.data_o [60]),
    .S(_26475_),
    .Z(_04421_));
 MUX2_X1 _58966_ (.A(\icache.data_set_select_mux.data_i [445]),
    .B(\icache.data_mems_6__data_mem.data_o [61]),
    .S(_26475_),
    .Z(_04422_));
 MUX2_X1 _58967_ (.A(\icache.data_set_select_mux.data_i [446]),
    .B(\icache.data_mems_6__data_mem.data_o [62]),
    .S(_26475_),
    .Z(_04423_));
 MUX2_X1 _58968_ (.A(\icache.data_set_select_mux.data_i [447]),
    .B(\icache.data_mems_6__data_mem.data_o [63]),
    .S(_26475_),
    .Z(_04424_));
 BUF_X4 _58969_ (.A(_26474_),
    .Z(_26476_));
 MUX2_X1 _58970_ (.A(\icache.data_set_select_mux.data_i [448]),
    .B(\icache.data_mems_7__data_mem.data_o [0]),
    .S(_26476_),
    .Z(_04425_));
 MUX2_X1 _58971_ (.A(\icache.data_set_select_mux.data_i [449]),
    .B(\icache.data_mems_7__data_mem.data_o [1]),
    .S(_26476_),
    .Z(_04426_));
 MUX2_X1 _58972_ (.A(\icache.data_set_select_mux.data_i [450]),
    .B(\icache.data_mems_7__data_mem.data_o [2]),
    .S(_26476_),
    .Z(_04428_));
 MUX2_X1 _58973_ (.A(\icache.data_set_select_mux.data_i [451]),
    .B(\icache.data_mems_7__data_mem.data_o [3]),
    .S(_26476_),
    .Z(_04429_));
 MUX2_X1 _58974_ (.A(\icache.data_set_select_mux.data_i [452]),
    .B(\icache.data_mems_7__data_mem.data_o [4]),
    .S(_26476_),
    .Z(_04430_));
 MUX2_X1 _58975_ (.A(\icache.data_set_select_mux.data_i [453]),
    .B(\icache.data_mems_7__data_mem.data_o [5]),
    .S(_26476_),
    .Z(_04431_));
 MUX2_X1 _58976_ (.A(\icache.data_set_select_mux.data_i [454]),
    .B(\icache.data_mems_7__data_mem.data_o [6]),
    .S(_26476_),
    .Z(_04432_));
 MUX2_X1 _58977_ (.A(\icache.data_set_select_mux.data_i [455]),
    .B(\icache.data_mems_7__data_mem.data_o [7]),
    .S(_26476_),
    .Z(_04433_));
 MUX2_X1 _58978_ (.A(\icache.data_set_select_mux.data_i [456]),
    .B(\icache.data_mems_7__data_mem.data_o [8]),
    .S(_26476_),
    .Z(_04434_));
 MUX2_X1 _58979_ (.A(\icache.data_set_select_mux.data_i [457]),
    .B(\icache.data_mems_7__data_mem.data_o [9]),
    .S(_26476_),
    .Z(_04435_));
 BUF_X4 _58980_ (.A(_26474_),
    .Z(_26477_));
 MUX2_X1 _58981_ (.A(\icache.data_set_select_mux.data_i [458]),
    .B(\icache.data_mems_7__data_mem.data_o [10]),
    .S(_26477_),
    .Z(_04436_));
 MUX2_X1 _58982_ (.A(\icache.data_set_select_mux.data_i [459]),
    .B(\icache.data_mems_7__data_mem.data_o [11]),
    .S(_26477_),
    .Z(_04437_));
 MUX2_X1 _58983_ (.A(\icache.data_set_select_mux.data_i [460]),
    .B(\icache.data_mems_7__data_mem.data_o [12]),
    .S(_26477_),
    .Z(_04439_));
 MUX2_X1 _58984_ (.A(\icache.data_set_select_mux.data_i [461]),
    .B(\icache.data_mems_7__data_mem.data_o [13]),
    .S(_26477_),
    .Z(_04440_));
 MUX2_X1 _58985_ (.A(\icache.data_set_select_mux.data_i [462]),
    .B(\icache.data_mems_7__data_mem.data_o [14]),
    .S(_26477_),
    .Z(_04441_));
 MUX2_X1 _58986_ (.A(\icache.data_set_select_mux.data_i [463]),
    .B(\icache.data_mems_7__data_mem.data_o [15]),
    .S(_26477_),
    .Z(_04442_));
 MUX2_X1 _58987_ (.A(\icache.data_set_select_mux.data_i [464]),
    .B(\icache.data_mems_7__data_mem.data_o [16]),
    .S(_26477_),
    .Z(_04443_));
 MUX2_X1 _58988_ (.A(\icache.data_set_select_mux.data_i [465]),
    .B(\icache.data_mems_7__data_mem.data_o [17]),
    .S(_26477_),
    .Z(_04444_));
 MUX2_X1 _58989_ (.A(\icache.data_set_select_mux.data_i [466]),
    .B(\icache.data_mems_7__data_mem.data_o [18]),
    .S(_26477_),
    .Z(_04445_));
 MUX2_X1 _58990_ (.A(\icache.data_set_select_mux.data_i [467]),
    .B(\icache.data_mems_7__data_mem.data_o [19]),
    .S(_26477_),
    .Z(_04446_));
 BUF_X4 _58991_ (.A(_26474_),
    .Z(_26478_));
 MUX2_X1 _58992_ (.A(\icache.data_set_select_mux.data_i [468]),
    .B(\icache.data_mems_7__data_mem.data_o [20]),
    .S(_26478_),
    .Z(_04447_));
 MUX2_X1 _58993_ (.A(\icache.data_set_select_mux.data_i [469]),
    .B(\icache.data_mems_7__data_mem.data_o [21]),
    .S(_26478_),
    .Z(_04448_));
 MUX2_X1 _58994_ (.A(\icache.data_set_select_mux.data_i [470]),
    .B(\icache.data_mems_7__data_mem.data_o [22]),
    .S(_26478_),
    .Z(_04450_));
 MUX2_X1 _58995_ (.A(\icache.data_set_select_mux.data_i [471]),
    .B(\icache.data_mems_7__data_mem.data_o [23]),
    .S(_26478_),
    .Z(_04451_));
 MUX2_X1 _58996_ (.A(\icache.data_set_select_mux.data_i [472]),
    .B(\icache.data_mems_7__data_mem.data_o [24]),
    .S(_26478_),
    .Z(_04452_));
 MUX2_X1 _58997_ (.A(\icache.data_set_select_mux.data_i [473]),
    .B(\icache.data_mems_7__data_mem.data_o [25]),
    .S(_26478_),
    .Z(_04453_));
 MUX2_X1 _58998_ (.A(\icache.data_set_select_mux.data_i [474]),
    .B(\icache.data_mems_7__data_mem.data_o [26]),
    .S(_26478_),
    .Z(_04454_));
 MUX2_X1 _58999_ (.A(\icache.data_set_select_mux.data_i [475]),
    .B(\icache.data_mems_7__data_mem.data_o [27]),
    .S(_26478_),
    .Z(_04455_));
 MUX2_X1 _59000_ (.A(\icache.data_set_select_mux.data_i [476]),
    .B(\icache.data_mems_7__data_mem.data_o [28]),
    .S(_26478_),
    .Z(_04456_));
 MUX2_X1 _59001_ (.A(\icache.data_set_select_mux.data_i [477]),
    .B(\icache.data_mems_7__data_mem.data_o [29]),
    .S(_26478_),
    .Z(_04457_));
 BUF_X4 _59002_ (.A(_26474_),
    .Z(_26479_));
 MUX2_X1 _59003_ (.A(\icache.data_set_select_mux.data_i [478]),
    .B(\icache.data_mems_7__data_mem.data_o [30]),
    .S(_26479_),
    .Z(_04458_));
 MUX2_X1 _59004_ (.A(\icache.data_set_select_mux.data_i [479]),
    .B(\icache.data_mems_7__data_mem.data_o [31]),
    .S(_26479_),
    .Z(_04459_));
 MUX2_X1 _59005_ (.A(\icache.data_set_select_mux.data_i [480]),
    .B(\icache.data_mems_7__data_mem.data_o [32]),
    .S(_26479_),
    .Z(_04461_));
 MUX2_X1 _59006_ (.A(\icache.data_set_select_mux.data_i [481]),
    .B(\icache.data_mems_7__data_mem.data_o [33]),
    .S(_26479_),
    .Z(_04462_));
 MUX2_X1 _59007_ (.A(\icache.data_set_select_mux.data_i [482]),
    .B(\icache.data_mems_7__data_mem.data_o [34]),
    .S(_26479_),
    .Z(_04463_));
 MUX2_X1 _59008_ (.A(\icache.data_set_select_mux.data_i [483]),
    .B(\icache.data_mems_7__data_mem.data_o [35]),
    .S(_26479_),
    .Z(_04464_));
 MUX2_X1 _59009_ (.A(\icache.data_set_select_mux.data_i [484]),
    .B(\icache.data_mems_7__data_mem.data_o [36]),
    .S(_26479_),
    .Z(_04465_));
 MUX2_X1 _59010_ (.A(\icache.data_set_select_mux.data_i [485]),
    .B(\icache.data_mems_7__data_mem.data_o [37]),
    .S(_26479_),
    .Z(_04466_));
 MUX2_X1 _59011_ (.A(\icache.data_set_select_mux.data_i [486]),
    .B(\icache.data_mems_7__data_mem.data_o [38]),
    .S(_26479_),
    .Z(_04467_));
 MUX2_X1 _59012_ (.A(\icache.data_set_select_mux.data_i [487]),
    .B(\icache.data_mems_7__data_mem.data_o [39]),
    .S(_26479_),
    .Z(_04468_));
 BUF_X8 _59013_ (.A(_26474_),
    .Z(_26480_));
 MUX2_X1 _59014_ (.A(\icache.data_set_select_mux.data_i [488]),
    .B(\icache.data_mems_7__data_mem.data_o [40]),
    .S(_26480_),
    .Z(_04469_));
 MUX2_X1 _59015_ (.A(\icache.data_set_select_mux.data_i [489]),
    .B(\icache.data_mems_7__data_mem.data_o [41]),
    .S(_26480_),
    .Z(_04470_));
 MUX2_X1 _59016_ (.A(\icache.data_set_select_mux.data_i [490]),
    .B(\icache.data_mems_7__data_mem.data_o [42]),
    .S(_26480_),
    .Z(_04472_));
 MUX2_X1 _59017_ (.A(\icache.data_set_select_mux.data_i [491]),
    .B(\icache.data_mems_7__data_mem.data_o [43]),
    .S(_26480_),
    .Z(_04473_));
 MUX2_X1 _59018_ (.A(\icache.data_set_select_mux.data_i [492]),
    .B(\icache.data_mems_7__data_mem.data_o [44]),
    .S(_26480_),
    .Z(_04474_));
 MUX2_X1 _59019_ (.A(\icache.data_set_select_mux.data_i [493]),
    .B(\icache.data_mems_7__data_mem.data_o [45]),
    .S(_26480_),
    .Z(_04475_));
 MUX2_X1 _59020_ (.A(\icache.data_set_select_mux.data_i [494]),
    .B(\icache.data_mems_7__data_mem.data_o [46]),
    .S(_26480_),
    .Z(_04476_));
 MUX2_X1 _59021_ (.A(\icache.data_set_select_mux.data_i [495]),
    .B(\icache.data_mems_7__data_mem.data_o [47]),
    .S(_26480_),
    .Z(_04477_));
 MUX2_X1 _59022_ (.A(\icache.data_set_select_mux.data_i [496]),
    .B(\icache.data_mems_7__data_mem.data_o [48]),
    .S(_26480_),
    .Z(_04478_));
 MUX2_X1 _59023_ (.A(\icache.data_set_select_mux.data_i [497]),
    .B(\icache.data_mems_7__data_mem.data_o [49]),
    .S(_26480_),
    .Z(_04479_));
 BUF_X8 _59024_ (.A(_26474_),
    .Z(_26481_));
 MUX2_X1 _59025_ (.A(\icache.data_set_select_mux.data_i [498]),
    .B(\icache.data_mems_7__data_mem.data_o [50]),
    .S(_26481_),
    .Z(_04480_));
 MUX2_X1 _59026_ (.A(\icache.data_set_select_mux.data_i [499]),
    .B(\icache.data_mems_7__data_mem.data_o [51]),
    .S(_26481_),
    .Z(_04481_));
 MUX2_X1 _59027_ (.A(\icache.data_set_select_mux.data_i [500]),
    .B(\icache.data_mems_7__data_mem.data_o [52]),
    .S(_26481_),
    .Z(_04484_));
 MUX2_X1 _59028_ (.A(\icache.data_set_select_mux.data_i [501]),
    .B(\icache.data_mems_7__data_mem.data_o [53]),
    .S(_26481_),
    .Z(_04485_));
 MUX2_X1 _59029_ (.A(\icache.data_set_select_mux.data_i [502]),
    .B(\icache.data_mems_7__data_mem.data_o [54]),
    .S(_26481_),
    .Z(_04486_));
 MUX2_X1 _59030_ (.A(\icache.data_set_select_mux.data_i [503]),
    .B(\icache.data_mems_7__data_mem.data_o [55]),
    .S(_26481_),
    .Z(_04487_));
 MUX2_X1 _59031_ (.A(\icache.data_set_select_mux.data_i [504]),
    .B(\icache.data_mems_7__data_mem.data_o [56]),
    .S(_26481_),
    .Z(_04488_));
 MUX2_X1 _59032_ (.A(\icache.data_set_select_mux.data_i [505]),
    .B(\icache.data_mems_7__data_mem.data_o [57]),
    .S(_26481_),
    .Z(_04489_));
 MUX2_X1 _59033_ (.A(\icache.data_set_select_mux.data_i [506]),
    .B(\icache.data_mems_7__data_mem.data_o [58]),
    .S(_26481_),
    .Z(_04490_));
 MUX2_X1 _59034_ (.A(\icache.data_set_select_mux.data_i [507]),
    .B(\icache.data_mems_7__data_mem.data_o [59]),
    .S(_26481_),
    .Z(_04491_));
 BUF_X8 _59035_ (.A(_26474_),
    .Z(_26482_));
 MUX2_X1 _59036_ (.A(\icache.data_set_select_mux.data_i [508]),
    .B(\icache.data_mems_7__data_mem.data_o [60]),
    .S(_26482_),
    .Z(_04492_));
 MUX2_X1 _59037_ (.A(\icache.data_set_select_mux.data_i [509]),
    .B(\icache.data_mems_7__data_mem.data_o [61]),
    .S(_26482_),
    .Z(_04493_));
 MUX2_X1 _59038_ (.A(\icache.data_set_select_mux.data_i [510]),
    .B(\icache.data_mems_7__data_mem.data_o [62]),
    .S(_26482_),
    .Z(_04495_));
 MUX2_X1 _59039_ (.A(\icache.data_set_select_mux.data_i [511]),
    .B(\icache.data_mems_7__data_mem.data_o [63]),
    .S(_26482_),
    .Z(_04496_));
 MUX2_X1 _59040_ (.A(\icache.N8 ),
    .B(\icache.uncached_i ),
    .S(_26482_),
    .Z(_04848_));
 OAI21_X1 _59041_ (.A(_07580_),
    .B1(_08017_),
    .B2(_08024_),
    .ZN(_26483_));
 MUX2_X1 _59042_ (.A(_00003_),
    .B(_26483_),
    .S(_21265_),
    .Z(_26484_));
 OAI211_X1 _59043_ (.A(_09118_),
    .B(_08727_),
    .C1(_26484_),
    .C2(_00000_),
    .ZN(_26485_));
 OAI21_X1 _59044_ (.A(_26485_),
    .B1(_09000_),
    .B2(_15277_),
    .ZN(_04847_));
 AND2_X2 _59045_ (.A1(_15276_),
    .A2(_08519_),
    .ZN(_26486_));
 BUF_X16 _59046_ (.A(_26486_),
    .Z(_26487_));
 BUF_X4 _59047_ (.A(_26487_),
    .Z(_26488_));
 MUX2_X1 _59048_ (.A(\icache.final_data_mux.data_i [64]),
    .B(_11246_),
    .S(_26488_),
    .Z(_04783_));
 MUX2_X1 _59049_ (.A(\icache.final_data_mux.data_i [65]),
    .B(_11314_),
    .S(_26488_),
    .Z(_04794_));
 MUX2_X1 _59050_ (.A(\icache.final_data_mux.data_i [66]),
    .B(_11349_),
    .S(_26488_),
    .Z(_04805_));
 MUX2_X1 _59051_ (.A(\icache.final_data_mux.data_i [67]),
    .B(_11382_),
    .S(_26488_),
    .Z(_04816_));
 MUX2_X1 _59052_ (.A(\icache.final_data_mux.data_i [68]),
    .B(_11416_),
    .S(_26488_),
    .Z(_04827_));
 MUX2_X1 _59053_ (.A(\icache.final_data_mux.data_i [69]),
    .B(_11450_),
    .S(_26488_),
    .Z(_04838_));
 MUX2_X1 _59054_ (.A(\icache.final_data_mux.data_i [70]),
    .B(_11483_),
    .S(_26488_),
    .Z(_04843_));
 MUX2_X1 _59055_ (.A(\icache.final_data_mux.data_i [71]),
    .B(_11498_),
    .S(_26488_),
    .Z(_04844_));
 MUX2_X1 _59056_ (.A(\icache.final_data_mux.data_i [72]),
    .B(_11549_),
    .S(_26488_),
    .Z(_04845_));
 MUX2_X1 _59057_ (.A(\icache.final_data_mux.data_i [73]),
    .B(_11566_),
    .S(_26488_),
    .Z(_04846_));
 BUF_X4 _59058_ (.A(_26487_),
    .Z(_26489_));
 MUX2_X1 _59059_ (.A(\icache.final_data_mux.data_i [74]),
    .B(_11599_),
    .S(_26489_),
    .Z(_04784_));
 MUX2_X1 _59060_ (.A(\icache.final_data_mux.data_i [75]),
    .B(_11632_),
    .S(_26489_),
    .Z(_04785_));
 MUX2_X1 _59061_ (.A(\icache.final_data_mux.data_i [76]),
    .B(_11688_),
    .S(_26489_),
    .Z(_04786_));
 MUX2_X1 _59062_ (.A(\icache.final_data_mux.data_i [77]),
    .B(_11722_),
    .S(_26489_),
    .Z(_04787_));
 MUX2_X1 _59063_ (.A(\icache.final_data_mux.data_i [78]),
    .B(_11755_),
    .S(_26489_),
    .Z(_04788_));
 MUX2_X1 _59064_ (.A(\icache.final_data_mux.data_i [79]),
    .B(_11789_),
    .S(_26489_),
    .Z(_04789_));
 MUX2_X1 _59065_ (.A(\icache.final_data_mux.data_i [80]),
    .B(_11804_),
    .S(_26489_),
    .Z(_04790_));
 MUX2_X1 _59066_ (.A(\icache.final_data_mux.data_i [81]),
    .B(_11856_),
    .S(_26489_),
    .Z(_04791_));
 MUX2_X1 _59067_ (.A(\icache.final_data_mux.data_i [82]),
    .B(_11888_),
    .S(_26489_),
    .Z(_04792_));
 MUX2_X1 _59068_ (.A(\icache.final_data_mux.data_i [83]),
    .B(_11921_),
    .S(_26489_),
    .Z(_04793_));
 BUF_X4 _59069_ (.A(_26487_),
    .Z(_26490_));
 MUX2_X1 _59070_ (.A(\icache.final_data_mux.data_i [84]),
    .B(_11937_),
    .S(_26490_),
    .Z(_04795_));
 MUX2_X1 _59071_ (.A(\icache.final_data_mux.data_i [85]),
    .B(_11988_),
    .S(_26490_),
    .Z(_04796_));
 MUX2_X1 _59072_ (.A(\icache.final_data_mux.data_i [86]),
    .B(_12005_),
    .S(_26490_),
    .Z(_04797_));
 MUX2_X1 _59073_ (.A(\icache.final_data_mux.data_i [87]),
    .B(_12054_),
    .S(_26490_),
    .Z(_04798_));
 MUX2_X1 _59074_ (.A(\icache.final_data_mux.data_i [88]),
    .B(_12089_),
    .S(_26490_),
    .Z(_04799_));
 MUX2_X1 _59075_ (.A(\icache.final_data_mux.data_i [89]),
    .B(_12121_),
    .S(_26490_),
    .Z(_04800_));
 MUX2_X1 _59076_ (.A(\icache.final_data_mux.data_i [90]),
    .B(_12156_),
    .S(_26490_),
    .Z(_04801_));
 MUX2_X1 _59077_ (.A(\icache.final_data_mux.data_i [91]),
    .B(_12188_),
    .S(_26490_),
    .Z(_04802_));
 MUX2_X1 _59078_ (.A(\icache.final_data_mux.data_i [92]),
    .B(_12222_),
    .S(_26490_),
    .Z(_04803_));
 MUX2_X1 _59079_ (.A(\icache.final_data_mux.data_i [93]),
    .B(_12255_),
    .S(_26490_),
    .Z(_04804_));
 BUF_X4 _59080_ (.A(_26487_),
    .Z(_26491_));
 MUX2_X1 _59081_ (.A(\icache.final_data_mux.data_i [94]),
    .B(_12286_),
    .S(_26491_),
    .Z(_04806_));
 MUX2_X1 _59082_ (.A(\icache.final_data_mux.data_i [95]),
    .B(_12307_),
    .S(_26491_),
    .Z(_04807_));
 MUX2_X1 _59083_ (.A(\icache.final_data_mux.data_i [96]),
    .B(_12340_),
    .S(_26491_),
    .Z(_04808_));
 MUX2_X1 _59084_ (.A(\icache.final_data_mux.data_i [97]),
    .B(_12391_),
    .S(_26491_),
    .Z(_04809_));
 MUX2_X1 _59085_ (.A(\icache.final_data_mux.data_i [98]),
    .B(_12425_),
    .S(_26491_),
    .Z(_04810_));
 MUX2_X1 _59086_ (.A(\icache.final_data_mux.data_i [99]),
    .B(_12456_),
    .S(_26491_),
    .Z(_04811_));
 MUX2_X1 _59087_ (.A(\icache.final_data_mux.data_i [100]),
    .B(_12492_),
    .S(_26491_),
    .Z(_04812_));
 MUX2_X1 _59088_ (.A(\icache.final_data_mux.data_i [101]),
    .B(_12525_),
    .S(_26491_),
    .Z(_04813_));
 MUX2_X1 _59089_ (.A(\icache.final_data_mux.data_i [102]),
    .B(_12557_),
    .S(_26491_),
    .Z(_04814_));
 MUX2_X1 _59090_ (.A(\icache.final_data_mux.data_i [103]),
    .B(_12573_),
    .S(_26491_),
    .Z(_04815_));
 BUF_X4 _59091_ (.A(_26487_),
    .Z(_26492_));
 MUX2_X1 _59092_ (.A(\icache.final_data_mux.data_i [104]),
    .B(_12626_),
    .S(_26492_),
    .Z(_04817_));
 MUX2_X1 _59093_ (.A(\icache.final_data_mux.data_i [105]),
    .B(_12644_),
    .S(_26492_),
    .Z(_04818_));
 MUX2_X1 _59094_ (.A(\icache.final_data_mux.data_i [106]),
    .B(_12677_),
    .S(_26492_),
    .Z(_04819_));
 MUX2_X1 _59095_ (.A(\icache.final_data_mux.data_i [107]),
    .B(_12711_),
    .S(_26492_),
    .Z(_04820_));
 MUX2_X1 _59096_ (.A(\icache.final_data_mux.data_i [108]),
    .B(_12760_),
    .S(_26492_),
    .Z(_04821_));
 MUX2_X1 _59097_ (.A(\icache.final_data_mux.data_i [109]),
    .B(_12794_),
    .S(_26492_),
    .Z(_04822_));
 MUX2_X1 _59098_ (.A(\icache.final_data_mux.data_i [110]),
    .B(_12826_),
    .S(_26492_),
    .Z(_04823_));
 MUX2_X1 _59099_ (.A(\icache.final_data_mux.data_i [111]),
    .B(_12859_),
    .S(_26492_),
    .Z(_04824_));
 MUX2_X1 _59100_ (.A(\icache.final_data_mux.data_i [112]),
    .B(_12874_),
    .S(_26492_),
    .Z(_04825_));
 MUX2_X1 _59101_ (.A(\icache.final_data_mux.data_i [113]),
    .B(_12925_),
    .S(_26492_),
    .Z(_04826_));
 BUF_X4 _59102_ (.A(_26487_),
    .Z(_26493_));
 MUX2_X1 _59103_ (.A(\icache.final_data_mux.data_i [114]),
    .B(_12957_),
    .S(_26493_),
    .Z(_04828_));
 MUX2_X1 _59104_ (.A(\icache.final_data_mux.data_i [115]),
    .B(_12992_),
    .S(_26493_),
    .Z(_04829_));
 MUX2_X1 _59105_ (.A(\icache.final_data_mux.data_i [116]),
    .B(_13009_),
    .S(_26493_),
    .Z(_04830_));
 MUX2_X1 _59106_ (.A(\icache.final_data_mux.data_i [117]),
    .B(_13058_),
    .S(_26493_),
    .Z(_04831_));
 MUX2_X1 _59107_ (.A(\icache.final_data_mux.data_i [118]),
    .B(_13074_),
    .S(_26493_),
    .Z(_04832_));
 MUX2_X1 _59108_ (.A(\icache.final_data_mux.data_i [119]),
    .B(_13122_),
    .S(_26493_),
    .Z(_04833_));
 MUX2_X1 _59109_ (.A(\icache.final_data_mux.data_i [120]),
    .B(_13157_),
    .S(_26493_),
    .Z(_04834_));
 MUX2_X1 _59110_ (.A(\icache.final_data_mux.data_i [121]),
    .B(_13192_),
    .S(_26493_),
    .Z(_04835_));
 MUX2_X1 _59111_ (.A(\icache.final_data_mux.data_i [122]),
    .B(_13224_),
    .S(_26493_),
    .Z(_04836_));
 MUX2_X1 _59112_ (.A(\icache.final_data_mux.data_i [123]),
    .B(_13256_),
    .S(_26493_),
    .Z(_04837_));
 MUX2_X1 _59113_ (.A(\icache.final_data_mux.data_i [124]),
    .B(_13288_),
    .S(_26487_),
    .Z(_04839_));
 MUX2_X1 _59114_ (.A(\icache.final_data_mux.data_i [125]),
    .B(_13322_),
    .S(_26487_),
    .Z(_04840_));
 MUX2_X1 _59115_ (.A(\icache.final_data_mux.data_i [126]),
    .B(_13357_),
    .S(_26487_),
    .Z(_04841_));
 MUX2_X1 _59116_ (.A(\icache.final_data_mux.data_i [127]),
    .B(_13372_),
    .S(_26487_),
    .Z(_04842_));
 MUX2_X1 _59117_ (.A(\icache.tag_tv_r [151]),
    .B(\icache.tag_mem.data_o [161]),
    .S(_26482_),
    .Z(_04624_));
 MUX2_X1 _59118_ (.A(\icache.tag_tv_r [152]),
    .B(\icache.tag_mem.data_o [162]),
    .S(_26482_),
    .Z(_04625_));
 MUX2_X1 _59119_ (.A(\icache.tag_tv_r [153]),
    .B(\icache.tag_mem.data_o [163]),
    .S(_26482_),
    .Z(_04626_));
 MUX2_X1 _59120_ (.A(\icache.tag_tv_r [154]),
    .B(\icache.tag_mem.data_o [164]),
    .S(_26482_),
    .Z(_04627_));
 MUX2_X1 _59121_ (.A(\icache.tag_tv_r [155]),
    .B(\icache.tag_mem.data_o [165]),
    .S(_26482_),
    .Z(_04628_));
 BUF_X4 _59122_ (.A(_26474_),
    .Z(_26494_));
 MUX2_X1 _59123_ (.A(\icache.tag_tv_r [156]),
    .B(\icache.tag_mem.data_o [166]),
    .S(_26494_),
    .Z(_04629_));
 MUX2_X1 _59124_ (.A(\icache.tag_tv_r [157]),
    .B(\icache.tag_mem.data_o [167]),
    .S(_26494_),
    .Z(_04630_));
 MUX2_X1 _59125_ (.A(\icache.tag_tv_r [158]),
    .B(\icache.tag_mem.data_o [168]),
    .S(_26494_),
    .Z(_04631_));
 MUX2_X1 _59126_ (.A(\icache.tag_tv_r [159]),
    .B(\icache.tag_mem.data_o [169]),
    .S(_26494_),
    .Z(_04632_));
 MUX2_X1 _59127_ (.A(\icache.tag_tv_r [160]),
    .B(\icache.tag_mem.data_o [170]),
    .S(_26494_),
    .Z(_04634_));
 MUX2_X1 _59128_ (.A(\icache.tag_tv_r [161]),
    .B(\icache.tag_mem.data_o [171]),
    .S(_26494_),
    .Z(_04635_));
 MUX2_X1 _59129_ (.A(\icache.tag_tv_r [162]),
    .B(\icache.tag_mem.data_o [174]),
    .S(_26494_),
    .Z(_04636_));
 MUX2_X1 _59130_ (.A(\icache.tag_tv_r [163]),
    .B(\icache.tag_mem.data_o [175]),
    .S(_26494_),
    .Z(_04637_));
 MUX2_X1 _59131_ (.A(\icache.tag_tv_r [164]),
    .B(\icache.tag_mem.data_o [176]),
    .S(_26494_),
    .Z(_04638_));
 MUX2_X1 _59132_ (.A(\icache.tag_tv_r [165]),
    .B(\icache.tag_mem.data_o [177]),
    .S(_26494_),
    .Z(_04639_));
 BUF_X4 _59133_ (.A(_26474_),
    .Z(_26495_));
 MUX2_X1 _59134_ (.A(\icache.tag_tv_r [166]),
    .B(\icache.tag_mem.data_o [178]),
    .S(_26495_),
    .Z(_04640_));
 MUX2_X1 _59135_ (.A(\icache.tag_tv_r [167]),
    .B(\icache.tag_mem.data_o [179]),
    .S(_26495_),
    .Z(_04641_));
 MUX2_X1 _59136_ (.A(\icache.tag_tv_r [168]),
    .B(\icache.tag_mem.data_o [180]),
    .S(_26495_),
    .Z(_04642_));
 MUX2_X1 _59137_ (.A(\icache.tag_tv_r [169]),
    .B(\icache.tag_mem.data_o [181]),
    .S(_26495_),
    .Z(_04643_));
 MUX2_X1 _59138_ (.A(\icache.tag_tv_r [170]),
    .B(\icache.tag_mem.data_o [182]),
    .S(_26495_),
    .Z(_04645_));
 MUX2_X1 _59139_ (.A(\icache.tag_tv_r [171]),
    .B(\icache.tag_mem.data_o [183]),
    .S(_26495_),
    .Z(_04646_));
 MUX2_X1 _59140_ (.A(\icache.tag_tv_r [172]),
    .B(\icache.tag_mem.data_o [184]),
    .S(_26495_),
    .Z(_04647_));
 MUX2_X1 _59141_ (.A(\icache.tag_tv_r [173]),
    .B(\icache.tag_mem.data_o [185]),
    .S(_26495_),
    .Z(_04648_));
 MUX2_X1 _59142_ (.A(\icache.tag_tv_r [174]),
    .B(\icache.tag_mem.data_o [186]),
    .S(_26495_),
    .Z(_04649_));
 MUX2_X1 _59143_ (.A(\icache.tag_tv_r [175]),
    .B(\icache.tag_mem.data_o [187]),
    .S(_26495_),
    .Z(_04650_));
 BUF_X16 _59144_ (.A(_26473_),
    .Z(_26496_));
 BUF_X4 _59145_ (.A(_26496_),
    .Z(_26497_));
 MUX2_X1 _59146_ (.A(\icache.tag_tv_r [176]),
    .B(\icache.tag_mem.data_o [188]),
    .S(_26497_),
    .Z(_04651_));
 MUX2_X1 _59147_ (.A(\icache.tag_tv_r [177]),
    .B(\icache.tag_mem.data_o [189]),
    .S(_26497_),
    .Z(_04652_));
 MUX2_X1 _59148_ (.A(\icache.tag_tv_r [178]),
    .B(\icache.tag_mem.data_o [190]),
    .S(_26497_),
    .Z(_04653_));
 MUX2_X1 _59149_ (.A(\icache.tag_tv_r [179]),
    .B(\icache.tag_mem.data_o [191]),
    .S(_26497_),
    .Z(_04654_));
 MUX2_X1 _59150_ (.A(\icache.tag_tv_r [180]),
    .B(\icache.tag_mem.data_o [192]),
    .S(_26497_),
    .Z(_04656_));
 MUX2_X1 _59151_ (.A(\icache.tag_tv_r [181]),
    .B(\icache.tag_mem.data_o [193]),
    .S(_26497_),
    .Z(_04657_));
 MUX2_X1 _59152_ (.A(\icache.tag_tv_r [182]),
    .B(\icache.tag_mem.data_o [194]),
    .S(_26497_),
    .Z(_04658_));
 MUX2_X1 _59153_ (.A(\icache.tag_tv_r [183]),
    .B(\icache.tag_mem.data_o [195]),
    .S(_26497_),
    .Z(_04659_));
 MUX2_X1 _59154_ (.A(\icache.tag_tv_r [184]),
    .B(\icache.tag_mem.data_o [196]),
    .S(_26497_),
    .Z(_04660_));
 MUX2_X1 _59155_ (.A(\icache.tag_tv_r [185]),
    .B(\icache.tag_mem.data_o [197]),
    .S(_26497_),
    .Z(_04661_));
 BUF_X4 _59156_ (.A(_26496_),
    .Z(_26498_));
 MUX2_X1 _59157_ (.A(\icache.tag_tv_r [186]),
    .B(\icache.tag_mem.data_o [198]),
    .S(_26498_),
    .Z(_04662_));
 MUX2_X1 _59158_ (.A(\icache.tag_tv_r [187]),
    .B(\icache.tag_mem.data_o [199]),
    .S(_26498_),
    .Z(_04663_));
 MUX2_X1 _59159_ (.A(\icache.tag_tv_r [188]),
    .B(\icache.tag_mem.data_o [200]),
    .S(_26498_),
    .Z(_04664_));
 MUX2_X1 _59160_ (.A(\icache.tag_tv_r [189]),
    .B(\icache.tag_mem.data_o [203]),
    .S(_26498_),
    .Z(_04665_));
 MUX2_X1 _59161_ (.A(\icache.tag_tv_r [190]),
    .B(\icache.tag_mem.data_o [204]),
    .S(_26498_),
    .Z(_04667_));
 MUX2_X1 _59162_ (.A(\icache.tag_tv_r [191]),
    .B(\icache.tag_mem.data_o [205]),
    .S(_26498_),
    .Z(_04668_));
 MUX2_X1 _59163_ (.A(\icache.tag_tv_r [192]),
    .B(\icache.tag_mem.data_o [206]),
    .S(_26498_),
    .Z(_04669_));
 MUX2_X1 _59164_ (.A(\icache.tag_tv_r [193]),
    .B(\icache.tag_mem.data_o [207]),
    .S(_26498_),
    .Z(_04670_));
 MUX2_X1 _59165_ (.A(\icache.tag_tv_r [194]),
    .B(\icache.tag_mem.data_o [208]),
    .S(_26498_),
    .Z(_04671_));
 MUX2_X1 _59166_ (.A(\icache.tag_tv_r [195]),
    .B(\icache.tag_mem.data_o [209]),
    .S(_26498_),
    .Z(_04672_));
 BUF_X4 _59167_ (.A(_26496_),
    .Z(_26499_));
 MUX2_X1 _59168_ (.A(\icache.tag_tv_r [196]),
    .B(\icache.tag_mem.data_o [210]),
    .S(_26499_),
    .Z(_04673_));
 MUX2_X1 _59169_ (.A(\icache.tag_tv_r [197]),
    .B(\icache.tag_mem.data_o [211]),
    .S(_26499_),
    .Z(_04674_));
 MUX2_X1 _59170_ (.A(\icache.tag_tv_r [198]),
    .B(\icache.tag_mem.data_o [212]),
    .S(_26499_),
    .Z(_04675_));
 MUX2_X1 _59171_ (.A(\icache.tag_tv_r [199]),
    .B(\icache.tag_mem.data_o [213]),
    .S(_26499_),
    .Z(_04676_));
 MUX2_X1 _59172_ (.A(\icache.tag_tv_r [200]),
    .B(\icache.tag_mem.data_o [214]),
    .S(_26499_),
    .Z(_04679_));
 MUX2_X1 _59173_ (.A(\icache.tag_tv_r [201]),
    .B(\icache.tag_mem.data_o [215]),
    .S(_26499_),
    .Z(_04680_));
 MUX2_X1 _59174_ (.A(\icache.tag_tv_r [202]),
    .B(\icache.tag_mem.data_o [216]),
    .S(_26499_),
    .Z(_04681_));
 MUX2_X1 _59175_ (.A(\icache.tag_tv_r [203]),
    .B(\icache.tag_mem.data_o [217]),
    .S(_26499_),
    .Z(_04682_));
 MUX2_X1 _59176_ (.A(\icache.tag_tv_r [204]),
    .B(\icache.tag_mem.data_o [218]),
    .S(_26499_),
    .Z(_04683_));
 MUX2_X1 _59177_ (.A(\icache.tag_tv_r [205]),
    .B(\icache.tag_mem.data_o [219]),
    .S(_26499_),
    .Z(_04684_));
 BUF_X4 _59178_ (.A(_26496_),
    .Z(_26500_));
 MUX2_X1 _59179_ (.A(\icache.tag_tv_r [206]),
    .B(\icache.tag_mem.data_o [220]),
    .S(_26500_),
    .Z(_04685_));
 MUX2_X1 _59180_ (.A(\icache.tag_tv_r [207]),
    .B(\icache.tag_mem.data_o [221]),
    .S(_26500_),
    .Z(_04686_));
 MUX2_X1 _59181_ (.A(\icache.tag_tv_r [208]),
    .B(\icache.tag_mem.data_o [222]),
    .S(_26500_),
    .Z(_04687_));
 MUX2_X1 _59182_ (.A(\icache.tag_tv_r [209]),
    .B(\icache.tag_mem.data_o [223]),
    .S(_26500_),
    .Z(_04688_));
 MUX2_X1 _59183_ (.A(\icache.tag_tv_r [210]),
    .B(\icache.tag_mem.data_o [224]),
    .S(_26500_),
    .Z(_04690_));
 MUX2_X1 _59184_ (.A(\icache.tag_tv_r [211]),
    .B(\icache.tag_mem.data_o [225]),
    .S(_26500_),
    .Z(_04691_));
 MUX2_X1 _59185_ (.A(\icache.tag_tv_r [212]),
    .B(\icache.tag_mem.data_o [226]),
    .S(_26500_),
    .Z(_04692_));
 MUX2_X1 _59186_ (.A(\icache.tag_tv_r [213]),
    .B(\icache.tag_mem.data_o [227]),
    .S(_26500_),
    .Z(_04693_));
 MUX2_X1 _59187_ (.A(\icache.tag_tv_r [214]),
    .B(\icache.tag_mem.data_o [228]),
    .S(_26500_),
    .Z(_04694_));
 MUX2_X1 _59188_ (.A(\icache.tag_tv_r [215]),
    .B(\icache.tag_mem.data_o [229]),
    .S(_26500_),
    .Z(_04695_));
 BUF_X16 _59189_ (.A(_26496_),
    .Z(_26501_));
 MUX2_X1 _59190_ (.A(\icache.state_tv_r [0]),
    .B(\icache.tag_mem.data_o [27]),
    .S(_26501_),
    .Z(_04551_));
 MUX2_X1 _59191_ (.A(\icache.state_tv_r [1]),
    .B(\icache.tag_mem.data_o [28]),
    .S(_26501_),
    .Z(_04558_));
 MUX2_X1 _59192_ (.A(\icache.state_tv_r [2]),
    .B(\icache.tag_mem.data_o [56]),
    .S(_26501_),
    .Z(_04559_));
 MUX2_X1 _59193_ (.A(\icache.state_tv_r [3]),
    .B(\icache.tag_mem.data_o [57]),
    .S(_26501_),
    .Z(_04560_));
 MUX2_X1 _59194_ (.A(\icache.state_tv_r [4]),
    .B(\icache.tag_mem.data_o [85]),
    .S(_26501_),
    .Z(_04561_));
 MUX2_X1 _59195_ (.A(\icache.state_tv_r [5]),
    .B(\icache.tag_mem.data_o [86]),
    .S(_26501_),
    .Z(_04562_));
 MUX2_X1 _59196_ (.A(\icache.state_tv_r [6]),
    .B(\icache.tag_mem.data_o [114]),
    .S(_26501_),
    .Z(_04563_));
 MUX2_X1 _59197_ (.A(\icache.state_tv_r [7]),
    .B(\icache.tag_mem.data_o [115]),
    .S(_26501_),
    .Z(_04564_));
 MUX2_X1 _59198_ (.A(\icache.state_tv_r [8]),
    .B(\icache.tag_mem.data_o [143]),
    .S(_26501_),
    .Z(_04565_));
 MUX2_X1 _59199_ (.A(\icache.state_tv_r [9]),
    .B(\icache.tag_mem.data_o [144]),
    .S(_26501_),
    .Z(_04566_));
 BUF_X16 _59200_ (.A(_26496_),
    .Z(_26502_));
 MUX2_X1 _59201_ (.A(\icache.state_tv_r [10]),
    .B(\icache.tag_mem.data_o [172]),
    .S(_26502_),
    .Z(_04552_));
 MUX2_X1 _59202_ (.A(\icache.state_tv_r [11]),
    .B(\icache.tag_mem.data_o [173]),
    .S(_26502_),
    .Z(_04553_));
 MUX2_X1 _59203_ (.A(\icache.state_tv_r [12]),
    .B(\icache.tag_mem.data_o [201]),
    .S(_26502_),
    .Z(_04554_));
 MUX2_X1 _59204_ (.A(\icache.state_tv_r [13]),
    .B(\icache.tag_mem.data_o [202]),
    .S(_26502_),
    .Z(_04555_));
 MUX2_X1 _59205_ (.A(\icache.state_tv_r [14]),
    .B(\icache.tag_mem.data_o [230]),
    .S(_26502_),
    .Z(_04556_));
 MUX2_X1 _59206_ (.A(\icache.state_tv_r [15]),
    .B(\icache.tag_mem.data_o [231]),
    .S(_26502_),
    .Z(_04557_));
 INV_X1 _59207_ (.A(_15279_),
    .ZN(_26503_));
 OAI211_X4 _59208_ (.A(_08499_),
    .B(_26503_),
    .C1(_08026_),
    .C2(_08035_),
    .ZN(_26504_));
 NOR2_X4 _59209_ (.A1(_26504_),
    .A2(_15274_),
    .ZN(_26505_));
 MUX2_X1 _59210_ (.A(_18116_),
    .B(_08492_),
    .S(_26505_),
    .Z(_04036_));
 MUX2_X1 _59211_ (.A(_16386_),
    .B(_08448_),
    .S(_26505_),
    .Z(_04037_));
 MUX2_X1 _59212_ (.A(_15580_),
    .B(_08434_),
    .S(_26505_),
    .Z(_04038_));
 MUX2_X1 _59213_ (.A(\icache.data_set_select_mux.data_i [315]),
    .B(\icache.data_mems_4__data_mem.data_o [59]),
    .S(_26502_),
    .Z(_04278_));
 MUX2_X1 _59214_ (.A(\icache.data_set_select_mux.data_i [316]),
    .B(\icache.data_mems_4__data_mem.data_o [60]),
    .S(_26502_),
    .Z(_04279_));
 MUX2_X1 _59215_ (.A(\icache.data_set_select_mux.data_i [317]),
    .B(\icache.data_mems_4__data_mem.data_o [61]),
    .S(_26502_),
    .Z(_04280_));
 MUX2_X1 _59216_ (.A(\icache.data_set_select_mux.data_i [318]),
    .B(\icache.data_mems_4__data_mem.data_o [62]),
    .S(_26502_),
    .Z(_04281_));
 BUF_X4 _59217_ (.A(_26496_),
    .Z(_26506_));
 MUX2_X1 _59218_ (.A(\icache.data_set_select_mux.data_i [319]),
    .B(\icache.data_mems_4__data_mem.data_o [63]),
    .S(_26506_),
    .Z(_04282_));
 MUX2_X1 _59219_ (.A(\icache.data_set_select_mux.data_i [320]),
    .B(\icache.data_mems_5__data_mem.data_o [0]),
    .S(_26506_),
    .Z(_04284_));
 MUX2_X1 _59220_ (.A(\icache.data_set_select_mux.data_i [321]),
    .B(\icache.data_mems_5__data_mem.data_o [1]),
    .S(_26506_),
    .Z(_04285_));
 MUX2_X1 _59221_ (.A(\icache.data_set_select_mux.data_i [322]),
    .B(\icache.data_mems_5__data_mem.data_o [2]),
    .S(_26506_),
    .Z(_04286_));
 MUX2_X1 _59222_ (.A(\icache.data_set_select_mux.data_i [323]),
    .B(\icache.data_mems_5__data_mem.data_o [3]),
    .S(_26506_),
    .Z(_04287_));
 MUX2_X1 _59223_ (.A(\icache.data_set_select_mux.data_i [324]),
    .B(\icache.data_mems_5__data_mem.data_o [4]),
    .S(_26506_),
    .Z(_04288_));
 MUX2_X1 _59224_ (.A(\icache.data_set_select_mux.data_i [325]),
    .B(\icache.data_mems_5__data_mem.data_o [5]),
    .S(_26506_),
    .Z(_04289_));
 MUX2_X1 _59225_ (.A(\icache.data_set_select_mux.data_i [326]),
    .B(\icache.data_mems_5__data_mem.data_o [6]),
    .S(_26506_),
    .Z(_04290_));
 MUX2_X1 _59226_ (.A(\icache.data_set_select_mux.data_i [327]),
    .B(\icache.data_mems_5__data_mem.data_o [7]),
    .S(_26506_),
    .Z(_04291_));
 MUX2_X1 _59227_ (.A(\icache.data_set_select_mux.data_i [328]),
    .B(\icache.data_mems_5__data_mem.data_o [8]),
    .S(_26506_),
    .Z(_04292_));
 BUF_X8 _59228_ (.A(_26496_),
    .Z(_26507_));
 MUX2_X1 _59229_ (.A(\icache.data_set_select_mux.data_i [329]),
    .B(\icache.data_mems_5__data_mem.data_o [9]),
    .S(_26507_),
    .Z(_04293_));
 MUX2_X1 _59230_ (.A(\icache.data_set_select_mux.data_i [330]),
    .B(\icache.data_mems_5__data_mem.data_o [10]),
    .S(_26507_),
    .Z(_04295_));
 MUX2_X1 _59231_ (.A(\icache.data_set_select_mux.data_i [331]),
    .B(\icache.data_mems_5__data_mem.data_o [11]),
    .S(_26507_),
    .Z(_04296_));
 MUX2_X1 _59232_ (.A(\icache.data_set_select_mux.data_i [332]),
    .B(\icache.data_mems_5__data_mem.data_o [12]),
    .S(_26507_),
    .Z(_04297_));
 MUX2_X1 _59233_ (.A(\icache.data_set_select_mux.data_i [333]),
    .B(\icache.data_mems_5__data_mem.data_o [13]),
    .S(_26507_),
    .Z(_04298_));
 MUX2_X1 _59234_ (.A(\icache.data_set_select_mux.data_i [334]),
    .B(\icache.data_mems_5__data_mem.data_o [14]),
    .S(_26507_),
    .Z(_04299_));
 MUX2_X1 _59235_ (.A(\icache.data_set_select_mux.data_i [335]),
    .B(\icache.data_mems_5__data_mem.data_o [15]),
    .S(_26507_),
    .Z(_04300_));
 MUX2_X1 _59236_ (.A(\icache.data_set_select_mux.data_i [336]),
    .B(\icache.data_mems_5__data_mem.data_o [16]),
    .S(_26507_),
    .Z(_04301_));
 MUX2_X1 _59237_ (.A(\icache.data_set_select_mux.data_i [337]),
    .B(\icache.data_mems_5__data_mem.data_o [17]),
    .S(_26507_),
    .Z(_04302_));
 MUX2_X1 _59238_ (.A(\icache.data_set_select_mux.data_i [338]),
    .B(\icache.data_mems_5__data_mem.data_o [18]),
    .S(_26507_),
    .Z(_04303_));
 BUF_X4 _59239_ (.A(_26496_),
    .Z(_26508_));
 MUX2_X1 _59240_ (.A(\icache.data_set_select_mux.data_i [339]),
    .B(\icache.data_mems_5__data_mem.data_o [19]),
    .S(_26508_),
    .Z(_04304_));
 MUX2_X1 _59241_ (.A(\icache.data_set_select_mux.data_i [340]),
    .B(\icache.data_mems_5__data_mem.data_o [20]),
    .S(_26508_),
    .Z(_04306_));
 MUX2_X1 _59242_ (.A(\icache.data_set_select_mux.data_i [341]),
    .B(\icache.data_mems_5__data_mem.data_o [21]),
    .S(_26508_),
    .Z(_04307_));
 MUX2_X1 _59243_ (.A(\icache.data_set_select_mux.data_i [342]),
    .B(\icache.data_mems_5__data_mem.data_o [22]),
    .S(_26508_),
    .Z(_04308_));
 MUX2_X1 _59244_ (.A(\icache.data_set_select_mux.data_i [343]),
    .B(\icache.data_mems_5__data_mem.data_o [23]),
    .S(_26508_),
    .Z(_04309_));
 MUX2_X1 _59245_ (.A(\icache.data_set_select_mux.data_i [344]),
    .B(\icache.data_mems_5__data_mem.data_o [24]),
    .S(_26508_),
    .Z(_04310_));
 MUX2_X1 _59246_ (.A(\icache.data_set_select_mux.data_i [345]),
    .B(\icache.data_mems_5__data_mem.data_o [25]),
    .S(_26508_),
    .Z(_04311_));
 MUX2_X1 _59247_ (.A(\icache.data_set_select_mux.data_i [346]),
    .B(\icache.data_mems_5__data_mem.data_o [26]),
    .S(_26508_),
    .Z(_04312_));
 MUX2_X1 _59248_ (.A(\icache.data_set_select_mux.data_i [347]),
    .B(\icache.data_mems_5__data_mem.data_o [27]),
    .S(_26508_),
    .Z(_04313_));
 MUX2_X1 _59249_ (.A(\icache.data_set_select_mux.data_i [348]),
    .B(\icache.data_mems_5__data_mem.data_o [28]),
    .S(_26508_),
    .Z(_04314_));
 BUF_X4 _59250_ (.A(_26496_),
    .Z(_26509_));
 MUX2_X1 _59251_ (.A(\icache.data_set_select_mux.data_i [349]),
    .B(\icache.data_mems_5__data_mem.data_o [29]),
    .S(_26509_),
    .Z(_04315_));
 MUX2_X1 _59252_ (.A(\icache.data_set_select_mux.data_i [350]),
    .B(\icache.data_mems_5__data_mem.data_o [30]),
    .S(_26509_),
    .Z(_04317_));
 MUX2_X1 _59253_ (.A(\icache.data_set_select_mux.data_i [351]),
    .B(\icache.data_mems_5__data_mem.data_o [31]),
    .S(_26509_),
    .Z(_04318_));
 MUX2_X1 _59254_ (.A(\icache.data_set_select_mux.data_i [352]),
    .B(\icache.data_mems_5__data_mem.data_o [32]),
    .S(_26509_),
    .Z(_04319_));
 MUX2_X1 _59255_ (.A(\icache.data_set_select_mux.data_i [353]),
    .B(\icache.data_mems_5__data_mem.data_o [33]),
    .S(_26509_),
    .Z(_04320_));
 MUX2_X1 _59256_ (.A(\icache.data_set_select_mux.data_i [354]),
    .B(\icache.data_mems_5__data_mem.data_o [34]),
    .S(_26509_),
    .Z(_04321_));
 MUX2_X1 _59257_ (.A(\icache.data_set_select_mux.data_i [355]),
    .B(\icache.data_mems_5__data_mem.data_o [35]),
    .S(_26509_),
    .Z(_04322_));
 MUX2_X1 _59258_ (.A(\icache.data_set_select_mux.data_i [356]),
    .B(\icache.data_mems_5__data_mem.data_o [36]),
    .S(_26509_),
    .Z(_04323_));
 MUX2_X1 _59259_ (.A(\icache.data_set_select_mux.data_i [357]),
    .B(\icache.data_mems_5__data_mem.data_o [37]),
    .S(_26509_),
    .Z(_04324_));
 MUX2_X1 _59260_ (.A(\icache.data_set_select_mux.data_i [358]),
    .B(\icache.data_mems_5__data_mem.data_o [38]),
    .S(_26509_),
    .Z(_04325_));
 BUF_X8 _59261_ (.A(_26473_),
    .Z(_26510_));
 BUF_X4 _59262_ (.A(_26510_),
    .Z(_26511_));
 MUX2_X1 _59263_ (.A(\icache.data_set_select_mux.data_i [359]),
    .B(\icache.data_mems_5__data_mem.data_o [39]),
    .S(_26511_),
    .Z(_04326_));
 MUX2_X1 _59264_ (.A(\icache.data_set_select_mux.data_i [360]),
    .B(\icache.data_mems_5__data_mem.data_o [40]),
    .S(_26511_),
    .Z(_04328_));
 MUX2_X1 _59265_ (.A(\icache.data_set_select_mux.data_i [361]),
    .B(\icache.data_mems_5__data_mem.data_o [41]),
    .S(_26511_),
    .Z(_04329_));
 MUX2_X1 _59266_ (.A(\icache.data_set_select_mux.data_i [362]),
    .B(\icache.data_mems_5__data_mem.data_o [42]),
    .S(_26511_),
    .Z(_04330_));
 MUX2_X1 _59267_ (.A(\icache.data_set_select_mux.data_i [363]),
    .B(\icache.data_mems_5__data_mem.data_o [43]),
    .S(_26511_),
    .Z(_04331_));
 MUX2_X1 _59268_ (.A(\icache.data_set_select_mux.data_i [364]),
    .B(\icache.data_mems_5__data_mem.data_o [44]),
    .S(_26511_),
    .Z(_04332_));
 MUX2_X1 _59269_ (.A(\icache.data_set_select_mux.data_i [365]),
    .B(\icache.data_mems_5__data_mem.data_o [45]),
    .S(_26511_),
    .Z(_04333_));
 MUX2_X1 _59270_ (.A(\icache.data_set_select_mux.data_i [366]),
    .B(\icache.data_mems_5__data_mem.data_o [46]),
    .S(_26511_),
    .Z(_04334_));
 MUX2_X1 _59271_ (.A(\icache.data_set_select_mux.data_i [367]),
    .B(\icache.data_mems_5__data_mem.data_o [47]),
    .S(_26511_),
    .Z(_04335_));
 MUX2_X1 _59272_ (.A(\icache.data_set_select_mux.data_i [368]),
    .B(\icache.data_mems_5__data_mem.data_o [48]),
    .S(_26511_),
    .Z(_04336_));
 BUF_X4 _59273_ (.A(_26510_),
    .Z(_26512_));
 MUX2_X1 _59274_ (.A(\icache.data_set_select_mux.data_i [369]),
    .B(\icache.data_mems_5__data_mem.data_o [49]),
    .S(_26512_),
    .Z(_04337_));
 MUX2_X1 _59275_ (.A(\icache.data_set_select_mux.data_i [370]),
    .B(\icache.data_mems_5__data_mem.data_o [50]),
    .S(_26512_),
    .Z(_04339_));
 MUX2_X1 _59276_ (.A(\icache.data_set_select_mux.data_i [371]),
    .B(\icache.data_mems_5__data_mem.data_o [51]),
    .S(_26512_),
    .Z(_04340_));
 MUX2_X1 _59277_ (.A(\icache.data_set_select_mux.data_i [372]),
    .B(\icache.data_mems_5__data_mem.data_o [52]),
    .S(_26512_),
    .Z(_04341_));
 MUX2_X1 _59278_ (.A(\icache.data_set_select_mux.data_i [373]),
    .B(\icache.data_mems_5__data_mem.data_o [53]),
    .S(_26512_),
    .Z(_04342_));
 MUX2_X1 _59279_ (.A(\icache.data_set_select_mux.data_i [374]),
    .B(\icache.data_mems_5__data_mem.data_o [54]),
    .S(_26512_),
    .Z(_04343_));
 MUX2_X1 _59280_ (.A(\icache.data_set_select_mux.data_i [375]),
    .B(\icache.data_mems_5__data_mem.data_o [55]),
    .S(_26512_),
    .Z(_04344_));
 MUX2_X1 _59281_ (.A(\icache.data_set_select_mux.data_i [376]),
    .B(\icache.data_mems_5__data_mem.data_o [56]),
    .S(_26512_),
    .Z(_04345_));
 MUX2_X1 _59282_ (.A(\icache.data_set_select_mux.data_i [377]),
    .B(\icache.data_mems_5__data_mem.data_o [57]),
    .S(_26512_),
    .Z(_04346_));
 MUX2_X1 _59283_ (.A(\icache.data_set_select_mux.data_i [378]),
    .B(\icache.data_mems_5__data_mem.data_o [58]),
    .S(_26512_),
    .Z(_04347_));
 BUF_X8 _59284_ (.A(_26510_),
    .Z(_26513_));
 MUX2_X1 _59285_ (.A(\icache.data_set_select_mux.data_i [379]),
    .B(\icache.data_mems_5__data_mem.data_o [59]),
    .S(_26513_),
    .Z(_04348_));
 MUX2_X1 _59286_ (.A(\icache.data_set_select_mux.data_i [380]),
    .B(\icache.data_mems_5__data_mem.data_o [60]),
    .S(_26513_),
    .Z(_04350_));
 MUX2_X1 _59287_ (.A(\icache.data_set_select_mux.data_i [381]),
    .B(\icache.data_mems_5__data_mem.data_o [61]),
    .S(_26513_),
    .Z(_04351_));
 MUX2_X1 _59288_ (.A(\icache.data_set_select_mux.data_i [382]),
    .B(\icache.data_mems_5__data_mem.data_o [62]),
    .S(_26513_),
    .Z(_04352_));
 MUX2_X1 _59289_ (.A(\icache.data_set_select_mux.data_i [383]),
    .B(\icache.data_mems_5__data_mem.data_o [63]),
    .S(_26513_),
    .Z(_04353_));
 MUX2_X1 _59290_ (.A(\icache.data_set_select_mux.data_i [384]),
    .B(\icache.data_mems_6__data_mem.data_o [0]),
    .S(_26513_),
    .Z(_04354_));
 MUX2_X1 _59291_ (.A(\icache.data_set_select_mux.data_i [385]),
    .B(\icache.data_mems_6__data_mem.data_o [1]),
    .S(_26513_),
    .Z(_04355_));
 MUX2_X1 _59292_ (.A(\icache.data_set_select_mux.data_i [386]),
    .B(\icache.data_mems_6__data_mem.data_o [2]),
    .S(_26513_),
    .Z(_04356_));
 MUX2_X1 _59293_ (.A(\icache.data_set_select_mux.data_i [387]),
    .B(\icache.data_mems_6__data_mem.data_o [3]),
    .S(_26513_),
    .Z(_04357_));
 MUX2_X1 _59294_ (.A(\icache.data_set_select_mux.data_i [388]),
    .B(\icache.data_mems_6__data_mem.data_o [4]),
    .S(_26513_),
    .Z(_04358_));
 BUF_X4 _59295_ (.A(_26510_),
    .Z(_26514_));
 MUX2_X1 _59296_ (.A(\icache.data_set_select_mux.data_i [389]),
    .B(\icache.data_mems_6__data_mem.data_o [5]),
    .S(_26514_),
    .Z(_04359_));
 MUX2_X1 _59297_ (.A(\icache.data_set_select_mux.data_i [390]),
    .B(\icache.data_mems_6__data_mem.data_o [6]),
    .S(_26514_),
    .Z(_04361_));
 MUX2_X1 _59298_ (.A(\icache.data_set_select_mux.data_i [391]),
    .B(\icache.data_mems_6__data_mem.data_o [7]),
    .S(_26514_),
    .Z(_04362_));
 MUX2_X1 _59299_ (.A(\icache.data_set_select_mux.data_i [392]),
    .B(\icache.data_mems_6__data_mem.data_o [8]),
    .S(_26514_),
    .Z(_04363_));
 MUX2_X1 _59300_ (.A(\icache.data_set_select_mux.data_i [393]),
    .B(\icache.data_mems_6__data_mem.data_o [9]),
    .S(_26514_),
    .Z(_04364_));
 MUX2_X1 _59301_ (.A(\icache.data_set_select_mux.data_i [394]),
    .B(\icache.data_mems_6__data_mem.data_o [10]),
    .S(_26514_),
    .Z(_04365_));
 MUX2_X1 _59302_ (.A(\icache.data_set_select_mux.data_i [395]),
    .B(\icache.data_mems_6__data_mem.data_o [11]),
    .S(_26514_),
    .Z(_04366_));
 MUX2_X1 _59303_ (.A(\icache.data_set_select_mux.data_i [396]),
    .B(\icache.data_mems_6__data_mem.data_o [12]),
    .S(_26514_),
    .Z(_04367_));
 MUX2_X1 _59304_ (.A(\icache.data_set_select_mux.data_i [397]),
    .B(\icache.data_mems_6__data_mem.data_o [13]),
    .S(_26514_),
    .Z(_04368_));
 MUX2_X1 _59305_ (.A(\icache.data_set_select_mux.data_i [398]),
    .B(\icache.data_mems_6__data_mem.data_o [14]),
    .S(_26514_),
    .Z(_04369_));
 BUF_X8 _59306_ (.A(_26510_),
    .Z(_26515_));
 MUX2_X1 _59307_ (.A(\icache.data_set_select_mux.data_i [399]),
    .B(\icache.data_mems_6__data_mem.data_o [15]),
    .S(_26515_),
    .Z(_04370_));
 MUX2_X1 _59308_ (.A(\icache.data_set_select_mux.data_i [400]),
    .B(\icache.data_mems_6__data_mem.data_o [16]),
    .S(_26515_),
    .Z(_04373_));
 MUX2_X1 _59309_ (.A(\icache.data_set_select_mux.data_i [401]),
    .B(\icache.data_mems_6__data_mem.data_o [17]),
    .S(_26515_),
    .Z(_04374_));
 MUX2_X1 _59310_ (.A(\icache.data_set_select_mux.data_i [402]),
    .B(\icache.data_mems_6__data_mem.data_o [18]),
    .S(_26515_),
    .Z(_04375_));
 MUX2_X1 _59311_ (.A(\icache.data_set_select_mux.data_i [403]),
    .B(\icache.data_mems_6__data_mem.data_o [19]),
    .S(_26515_),
    .Z(_04376_));
 MUX2_X1 _59312_ (.A(\icache.data_set_select_mux.data_i [404]),
    .B(\icache.data_mems_6__data_mem.data_o [20]),
    .S(_26515_),
    .Z(_04377_));
 MUX2_X1 _59313_ (.A(\icache.data_set_select_mux.data_i [405]),
    .B(\icache.data_mems_6__data_mem.data_o [21]),
    .S(_26515_),
    .Z(_04378_));
 MUX2_X1 _59314_ (.A(\icache.data_set_select_mux.data_i [406]),
    .B(\icache.data_mems_6__data_mem.data_o [22]),
    .S(_26515_),
    .Z(_04379_));
 MUX2_X1 _59315_ (.A(\icache.data_set_select_mux.data_i [407]),
    .B(\icache.data_mems_6__data_mem.data_o [23]),
    .S(_26515_),
    .Z(_04380_));
 MUX2_X1 _59316_ (.A(\icache.data_set_select_mux.data_i [408]),
    .B(\icache.data_mems_6__data_mem.data_o [24]),
    .S(_26515_),
    .Z(_04381_));
 BUF_X8 _59317_ (.A(_26510_),
    .Z(_26516_));
 MUX2_X1 _59318_ (.A(\icache.data_set_select_mux.data_i [409]),
    .B(\icache.data_mems_6__data_mem.data_o [25]),
    .S(_26516_),
    .Z(_04382_));
 MUX2_X1 _59319_ (.A(\icache.data_set_select_mux.data_i [410]),
    .B(\icache.data_mems_6__data_mem.data_o [26]),
    .S(_26516_),
    .Z(_04384_));
 MUX2_X1 _59320_ (.A(\icache.data_set_select_mux.data_i [411]),
    .B(\icache.data_mems_6__data_mem.data_o [27]),
    .S(_26516_),
    .Z(_04385_));
 MUX2_X1 _59321_ (.A(\icache.data_set_select_mux.data_i [412]),
    .B(\icache.data_mems_6__data_mem.data_o [28]),
    .S(_26516_),
    .Z(_04386_));
 MUX2_X1 _59322_ (.A(\icache.data_set_select_mux.data_i [413]),
    .B(\icache.data_mems_6__data_mem.data_o [29]),
    .S(_26516_),
    .Z(_04387_));
 MUX2_X1 _59323_ (.A(\icache.addr_tv_r [0]),
    .B(\icache.vaddr_tl_r [0]),
    .S(_26516_),
    .Z(_03958_));
 MUX2_X1 _59324_ (.A(\icache.data_set_select_mux.data_i [216]),
    .B(\icache.data_mems_3__data_mem.data_o [24]),
    .S(_26516_),
    .Z(_04168_));
 MUX2_X1 _59325_ (.A(\icache.data_set_select_mux.data_i [217]),
    .B(\icache.data_mems_3__data_mem.data_o [25]),
    .S(_26516_),
    .Z(_04169_));
 MUX2_X1 _59326_ (.A(\icache.data_set_select_mux.data_i [218]),
    .B(\icache.data_mems_3__data_mem.data_o [26]),
    .S(_26516_),
    .Z(_04170_));
 MUX2_X1 _59327_ (.A(\icache.data_set_select_mux.data_i [219]),
    .B(\icache.data_mems_3__data_mem.data_o [27]),
    .S(_26516_),
    .Z(_04171_));
 BUF_X8 _59328_ (.A(_26510_),
    .Z(_26517_));
 MUX2_X1 _59329_ (.A(\icache.data_set_select_mux.data_i [220]),
    .B(\icache.data_mems_3__data_mem.data_o [28]),
    .S(_26517_),
    .Z(_04173_));
 MUX2_X1 _59330_ (.A(\icache.data_set_select_mux.data_i [221]),
    .B(\icache.data_mems_3__data_mem.data_o [29]),
    .S(_26517_),
    .Z(_04174_));
 MUX2_X1 _59331_ (.A(\icache.data_set_select_mux.data_i [222]),
    .B(\icache.data_mems_3__data_mem.data_o [30]),
    .S(_26517_),
    .Z(_04175_));
 MUX2_X1 _59332_ (.A(\icache.data_set_select_mux.data_i [223]),
    .B(\icache.data_mems_3__data_mem.data_o [31]),
    .S(_26517_),
    .Z(_04176_));
 MUX2_X1 _59333_ (.A(\icache.data_set_select_mux.data_i [224]),
    .B(\icache.data_mems_3__data_mem.data_o [32]),
    .S(_26517_),
    .Z(_04177_));
 MUX2_X1 _59334_ (.A(\icache.data_set_select_mux.data_i [225]),
    .B(\icache.data_mems_3__data_mem.data_o [33]),
    .S(_26517_),
    .Z(_04178_));
 MUX2_X1 _59335_ (.A(\icache.data_set_select_mux.data_i [226]),
    .B(\icache.data_mems_3__data_mem.data_o [34]),
    .S(_26517_),
    .Z(_04179_));
 MUX2_X1 _59336_ (.A(\icache.data_set_select_mux.data_i [227]),
    .B(\icache.data_mems_3__data_mem.data_o [35]),
    .S(_26517_),
    .Z(_04180_));
 MUX2_X1 _59337_ (.A(\icache.data_set_select_mux.data_i [228]),
    .B(\icache.data_mems_3__data_mem.data_o [36]),
    .S(_26517_),
    .Z(_04181_));
 MUX2_X1 _59338_ (.A(\icache.data_set_select_mux.data_i [229]),
    .B(\icache.data_mems_3__data_mem.data_o [37]),
    .S(_26517_),
    .Z(_04182_));
 BUF_X4 _59339_ (.A(_26510_),
    .Z(_26518_));
 MUX2_X1 _59340_ (.A(\icache.data_set_select_mux.data_i [230]),
    .B(\icache.data_mems_3__data_mem.data_o [38]),
    .S(_26518_),
    .Z(_04184_));
 MUX2_X1 _59341_ (.A(\icache.data_set_select_mux.data_i [231]),
    .B(\icache.data_mems_3__data_mem.data_o [39]),
    .S(_26518_),
    .Z(_04185_));
 MUX2_X1 _59342_ (.A(\icache.data_set_select_mux.data_i [232]),
    .B(\icache.data_mems_3__data_mem.data_o [40]),
    .S(_26518_),
    .Z(_04186_));
 MUX2_X1 _59343_ (.A(\icache.data_set_select_mux.data_i [233]),
    .B(\icache.data_mems_3__data_mem.data_o [41]),
    .S(_26518_),
    .Z(_04187_));
 MUX2_X1 _59344_ (.A(\icache.data_set_select_mux.data_i [234]),
    .B(\icache.data_mems_3__data_mem.data_o [42]),
    .S(_26518_),
    .Z(_04188_));
 MUX2_X1 _59345_ (.A(\icache.data_set_select_mux.data_i [235]),
    .B(\icache.data_mems_3__data_mem.data_o [43]),
    .S(_26518_),
    .Z(_04189_));
 MUX2_X1 _59346_ (.A(\icache.data_set_select_mux.data_i [236]),
    .B(\icache.data_mems_3__data_mem.data_o [44]),
    .S(_26518_),
    .Z(_04190_));
 MUX2_X1 _59347_ (.A(\icache.data_set_select_mux.data_i [237]),
    .B(\icache.data_mems_3__data_mem.data_o [45]),
    .S(_26518_),
    .Z(_04191_));
 MUX2_X1 _59348_ (.A(\icache.data_set_select_mux.data_i [238]),
    .B(\icache.data_mems_3__data_mem.data_o [46]),
    .S(_26518_),
    .Z(_04192_));
 MUX2_X1 _59349_ (.A(\icache.data_set_select_mux.data_i [239]),
    .B(\icache.data_mems_3__data_mem.data_o [47]),
    .S(_26518_),
    .Z(_04193_));
 BUF_X8 _59350_ (.A(_26510_),
    .Z(_26519_));
 MUX2_X1 _59351_ (.A(\icache.data_set_select_mux.data_i [240]),
    .B(\icache.data_mems_3__data_mem.data_o [48]),
    .S(_26519_),
    .Z(_04195_));
 MUX2_X1 _59352_ (.A(\icache.data_set_select_mux.data_i [241]),
    .B(\icache.data_mems_3__data_mem.data_o [49]),
    .S(_26519_),
    .Z(_04196_));
 MUX2_X1 _59353_ (.A(\icache.data_set_select_mux.data_i [242]),
    .B(\icache.data_mems_3__data_mem.data_o [50]),
    .S(_26519_),
    .Z(_04197_));
 MUX2_X1 _59354_ (.A(\icache.data_set_select_mux.data_i [243]),
    .B(\icache.data_mems_3__data_mem.data_o [51]),
    .S(_26519_),
    .Z(_04198_));
 MUX2_X1 _59355_ (.A(\icache.data_set_select_mux.data_i [244]),
    .B(\icache.data_mems_3__data_mem.data_o [52]),
    .S(_26519_),
    .Z(_04199_));
 MUX2_X1 _59356_ (.A(\icache.data_set_select_mux.data_i [245]),
    .B(\icache.data_mems_3__data_mem.data_o [53]),
    .S(_26519_),
    .Z(_04200_));
 MUX2_X1 _59357_ (.A(\icache.data_set_select_mux.data_i [246]),
    .B(\icache.data_mems_3__data_mem.data_o [54]),
    .S(_26519_),
    .Z(_04201_));
 MUX2_X1 _59358_ (.A(\icache.data_set_select_mux.data_i [247]),
    .B(\icache.data_mems_3__data_mem.data_o [55]),
    .S(_26519_),
    .Z(_04202_));
 MUX2_X1 _59359_ (.A(\icache.data_set_select_mux.data_i [248]),
    .B(\icache.data_mems_3__data_mem.data_o [56]),
    .S(_26519_),
    .Z(_04203_));
 MUX2_X1 _59360_ (.A(\icache.data_set_select_mux.data_i [249]),
    .B(\icache.data_mems_3__data_mem.data_o [57]),
    .S(_26519_),
    .Z(_04204_));
 BUF_X8 _59361_ (.A(_26510_),
    .Z(_26520_));
 MUX2_X1 _59362_ (.A(\icache.data_set_select_mux.data_i [250]),
    .B(\icache.data_mems_3__data_mem.data_o [58]),
    .S(_26520_),
    .Z(_04206_));
 MUX2_X1 _59363_ (.A(\icache.data_set_select_mux.data_i [251]),
    .B(\icache.data_mems_3__data_mem.data_o [59]),
    .S(_26520_),
    .Z(_04207_));
 MUX2_X1 _59364_ (.A(\icache.data_set_select_mux.data_i [252]),
    .B(\icache.data_mems_3__data_mem.data_o [60]),
    .S(_26520_),
    .Z(_04208_));
 MUX2_X1 _59365_ (.A(\icache.data_set_select_mux.data_i [253]),
    .B(\icache.data_mems_3__data_mem.data_o [61]),
    .S(_26520_),
    .Z(_04209_));
 MUX2_X1 _59366_ (.A(\icache.data_set_select_mux.data_i [254]),
    .B(\icache.data_mems_3__data_mem.data_o [62]),
    .S(_26520_),
    .Z(_04210_));
 MUX2_X1 _59367_ (.A(\icache.data_set_select_mux.data_i [255]),
    .B(\icache.data_mems_3__data_mem.data_o [63]),
    .S(_26520_),
    .Z(_04211_));
 MUX2_X1 _59368_ (.A(\icache.data_set_select_mux.data_i [256]),
    .B(\icache.data_mems_4__data_mem.data_o [0]),
    .S(_26520_),
    .Z(_04212_));
 MUX2_X1 _59369_ (.A(\icache.data_set_select_mux.data_i [257]),
    .B(\icache.data_mems_4__data_mem.data_o [1]),
    .S(_26520_),
    .Z(_04213_));
 MUX2_X1 _59370_ (.A(\icache.data_set_select_mux.data_i [258]),
    .B(\icache.data_mems_4__data_mem.data_o [2]),
    .S(_26520_),
    .Z(_04214_));
 MUX2_X1 _59371_ (.A(\icache.data_set_select_mux.data_i [259]),
    .B(\icache.data_mems_4__data_mem.data_o [3]),
    .S(_26520_),
    .Z(_04215_));
 BUF_X16 _59372_ (.A(_26473_),
    .Z(_26521_));
 BUF_X4 _59373_ (.A(_26521_),
    .Z(_26522_));
 MUX2_X1 _59374_ (.A(\icache.data_set_select_mux.data_i [260]),
    .B(\icache.data_mems_4__data_mem.data_o [4]),
    .S(_26522_),
    .Z(_04217_));
 MUX2_X1 _59375_ (.A(\icache.data_set_select_mux.data_i [261]),
    .B(\icache.data_mems_4__data_mem.data_o [5]),
    .S(_26522_),
    .Z(_04218_));
 MUX2_X1 _59376_ (.A(\icache.data_set_select_mux.data_i [262]),
    .B(\icache.data_mems_4__data_mem.data_o [6]),
    .S(_26522_),
    .Z(_04219_));
 MUX2_X1 _59377_ (.A(\icache.data_set_select_mux.data_i [263]),
    .B(\icache.data_mems_4__data_mem.data_o [7]),
    .S(_26522_),
    .Z(_04220_));
 MUX2_X1 _59378_ (.A(\icache.data_set_select_mux.data_i [264]),
    .B(\icache.data_mems_4__data_mem.data_o [8]),
    .S(_26522_),
    .Z(_04221_));
 MUX2_X1 _59379_ (.A(\icache.data_set_select_mux.data_i [265]),
    .B(\icache.data_mems_4__data_mem.data_o [9]),
    .S(_26522_),
    .Z(_04222_));
 MUX2_X1 _59380_ (.A(\icache.data_set_select_mux.data_i [266]),
    .B(\icache.data_mems_4__data_mem.data_o [10]),
    .S(_26522_),
    .Z(_04223_));
 MUX2_X1 _59381_ (.A(\icache.data_set_select_mux.data_i [267]),
    .B(\icache.data_mems_4__data_mem.data_o [11]),
    .S(_26522_),
    .Z(_04224_));
 MUX2_X1 _59382_ (.A(\icache.data_set_select_mux.data_i [268]),
    .B(\icache.data_mems_4__data_mem.data_o [12]),
    .S(_26522_),
    .Z(_04225_));
 MUX2_X1 _59383_ (.A(\icache.data_set_select_mux.data_i [269]),
    .B(\icache.data_mems_4__data_mem.data_o [13]),
    .S(_26522_),
    .Z(_04226_));
 BUF_X4 _59384_ (.A(_26521_),
    .Z(_26523_));
 MUX2_X1 _59385_ (.A(\icache.data_set_select_mux.data_i [270]),
    .B(\icache.data_mems_4__data_mem.data_o [14]),
    .S(_26523_),
    .Z(_04228_));
 MUX2_X1 _59386_ (.A(\icache.data_set_select_mux.data_i [271]),
    .B(\icache.data_mems_4__data_mem.data_o [15]),
    .S(_26523_),
    .Z(_04229_));
 MUX2_X1 _59387_ (.A(\icache.data_set_select_mux.data_i [272]),
    .B(\icache.data_mems_4__data_mem.data_o [16]),
    .S(_26523_),
    .Z(_04230_));
 MUX2_X1 _59388_ (.A(\icache.data_set_select_mux.data_i [273]),
    .B(\icache.data_mems_4__data_mem.data_o [17]),
    .S(_26523_),
    .Z(_04231_));
 MUX2_X1 _59389_ (.A(\icache.data_set_select_mux.data_i [274]),
    .B(\icache.data_mems_4__data_mem.data_o [18]),
    .S(_26523_),
    .Z(_04232_));
 MUX2_X1 _59390_ (.A(\icache.data_set_select_mux.data_i [275]),
    .B(\icache.data_mems_4__data_mem.data_o [19]),
    .S(_26523_),
    .Z(_04233_));
 MUX2_X1 _59391_ (.A(\icache.data_set_select_mux.data_i [276]),
    .B(\icache.data_mems_4__data_mem.data_o [20]),
    .S(_26523_),
    .Z(_04234_));
 MUX2_X1 _59392_ (.A(\icache.data_set_select_mux.data_i [277]),
    .B(\icache.data_mems_4__data_mem.data_o [21]),
    .S(_26523_),
    .Z(_04235_));
 MUX2_X1 _59393_ (.A(\icache.data_set_select_mux.data_i [278]),
    .B(\icache.data_mems_4__data_mem.data_o [22]),
    .S(_26523_),
    .Z(_04236_));
 MUX2_X1 _59394_ (.A(\icache.data_set_select_mux.data_i [279]),
    .B(\icache.data_mems_4__data_mem.data_o [23]),
    .S(_26523_),
    .Z(_04237_));
 BUF_X4 _59395_ (.A(_26521_),
    .Z(_26524_));
 MUX2_X1 _59396_ (.A(\icache.data_set_select_mux.data_i [280]),
    .B(\icache.data_mems_4__data_mem.data_o [24]),
    .S(_26524_),
    .Z(_04239_));
 MUX2_X1 _59397_ (.A(\icache.data_set_select_mux.data_i [281]),
    .B(\icache.data_mems_4__data_mem.data_o [25]),
    .S(_26524_),
    .Z(_04240_));
 MUX2_X1 _59398_ (.A(\icache.data_set_select_mux.data_i [282]),
    .B(\icache.data_mems_4__data_mem.data_o [26]),
    .S(_26524_),
    .Z(_04241_));
 MUX2_X1 _59399_ (.A(\icache.data_set_select_mux.data_i [283]),
    .B(\icache.data_mems_4__data_mem.data_o [27]),
    .S(_26524_),
    .Z(_04242_));
 MUX2_X1 _59400_ (.A(\icache.data_set_select_mux.data_i [284]),
    .B(\icache.data_mems_4__data_mem.data_o [28]),
    .S(_26524_),
    .Z(_04243_));
 MUX2_X1 _59401_ (.A(\icache.data_set_select_mux.data_i [285]),
    .B(\icache.data_mems_4__data_mem.data_o [29]),
    .S(_26524_),
    .Z(_04244_));
 MUX2_X1 _59402_ (.A(\icache.data_set_select_mux.data_i [286]),
    .B(\icache.data_mems_4__data_mem.data_o [30]),
    .S(_26524_),
    .Z(_04245_));
 MUX2_X1 _59403_ (.A(\icache.data_set_select_mux.data_i [287]),
    .B(\icache.data_mems_4__data_mem.data_o [31]),
    .S(_26524_),
    .Z(_04246_));
 MUX2_X1 _59404_ (.A(\icache.data_set_select_mux.data_i [288]),
    .B(\icache.data_mems_4__data_mem.data_o [32]),
    .S(_26524_),
    .Z(_04247_));
 MUX2_X1 _59405_ (.A(\icache.data_set_select_mux.data_i [289]),
    .B(\icache.data_mems_4__data_mem.data_o [33]),
    .S(_26524_),
    .Z(_04248_));
 BUF_X4 _59406_ (.A(_26521_),
    .Z(_26525_));
 MUX2_X1 _59407_ (.A(\icache.data_set_select_mux.data_i [290]),
    .B(\icache.data_mems_4__data_mem.data_o [34]),
    .S(_26525_),
    .Z(_04250_));
 MUX2_X1 _59408_ (.A(\icache.data_set_select_mux.data_i [291]),
    .B(\icache.data_mems_4__data_mem.data_o [35]),
    .S(_26525_),
    .Z(_04251_));
 MUX2_X1 _59409_ (.A(\icache.data_set_select_mux.data_i [292]),
    .B(\icache.data_mems_4__data_mem.data_o [36]),
    .S(_26525_),
    .Z(_04252_));
 MUX2_X1 _59410_ (.A(\icache.data_set_select_mux.data_i [293]),
    .B(\icache.data_mems_4__data_mem.data_o [37]),
    .S(_26525_),
    .Z(_04253_));
 MUX2_X1 _59411_ (.A(\icache.data_set_select_mux.data_i [294]),
    .B(\icache.data_mems_4__data_mem.data_o [38]),
    .S(_26525_),
    .Z(_04254_));
 MUX2_X1 _59412_ (.A(\icache.data_set_select_mux.data_i [295]),
    .B(\icache.data_mems_4__data_mem.data_o [39]),
    .S(_26525_),
    .Z(_04255_));
 MUX2_X1 _59413_ (.A(\icache.data_set_select_mux.data_i [296]),
    .B(\icache.data_mems_4__data_mem.data_o [40]),
    .S(_26525_),
    .Z(_04256_));
 MUX2_X1 _59414_ (.A(\icache.data_set_select_mux.data_i [297]),
    .B(\icache.data_mems_4__data_mem.data_o [41]),
    .S(_26525_),
    .Z(_04257_));
 MUX2_X1 _59415_ (.A(\icache.data_set_select_mux.data_i [298]),
    .B(\icache.data_mems_4__data_mem.data_o [42]),
    .S(_26525_),
    .Z(_04258_));
 MUX2_X1 _59416_ (.A(\icache.data_set_select_mux.data_i [299]),
    .B(\icache.data_mems_4__data_mem.data_o [43]),
    .S(_26525_),
    .Z(_04259_));
 BUF_X4 _59417_ (.A(_26521_),
    .Z(_26526_));
 MUX2_X1 _59418_ (.A(\icache.data_set_select_mux.data_i [300]),
    .B(\icache.data_mems_4__data_mem.data_o [44]),
    .S(_26526_),
    .Z(_04262_));
 MUX2_X1 _59419_ (.A(\icache.data_set_select_mux.data_i [301]),
    .B(\icache.data_mems_4__data_mem.data_o [45]),
    .S(_26526_),
    .Z(_04263_));
 MUX2_X1 _59420_ (.A(\icache.data_set_select_mux.data_i [302]),
    .B(\icache.data_mems_4__data_mem.data_o [46]),
    .S(_26526_),
    .Z(_04264_));
 MUX2_X1 _59421_ (.A(\icache.data_set_select_mux.data_i [303]),
    .B(\icache.data_mems_4__data_mem.data_o [47]),
    .S(_26526_),
    .Z(_04265_));
 MUX2_X1 _59422_ (.A(\icache.data_set_select_mux.data_i [304]),
    .B(\icache.data_mems_4__data_mem.data_o [48]),
    .S(_26526_),
    .Z(_04266_));
 MUX2_X1 _59423_ (.A(\icache.data_set_select_mux.data_i [305]),
    .B(\icache.data_mems_4__data_mem.data_o [49]),
    .S(_26526_),
    .Z(_04267_));
 MUX2_X1 _59424_ (.A(\icache.data_set_select_mux.data_i [306]),
    .B(\icache.data_mems_4__data_mem.data_o [50]),
    .S(_26526_),
    .Z(_04268_));
 MUX2_X1 _59425_ (.A(\icache.data_set_select_mux.data_i [307]),
    .B(\icache.data_mems_4__data_mem.data_o [51]),
    .S(_26526_),
    .Z(_04269_));
 MUX2_X1 _59426_ (.A(\icache.data_set_select_mux.data_i [308]),
    .B(\icache.data_mems_4__data_mem.data_o [52]),
    .S(_26526_),
    .Z(_04270_));
 MUX2_X1 _59427_ (.A(\icache.data_set_select_mux.data_i [309]),
    .B(\icache.data_mems_4__data_mem.data_o [53]),
    .S(_26526_),
    .Z(_04271_));
 BUF_X8 _59428_ (.A(_26521_),
    .Z(_26527_));
 MUX2_X1 _59429_ (.A(\icache.data_set_select_mux.data_i [310]),
    .B(\icache.data_mems_4__data_mem.data_o [54]),
    .S(_26527_),
    .Z(_04273_));
 MUX2_X1 _59430_ (.A(\icache.data_set_select_mux.data_i [311]),
    .B(\icache.data_mems_4__data_mem.data_o [55]),
    .S(_26527_),
    .Z(_04274_));
 MUX2_X1 _59431_ (.A(\icache.data_set_select_mux.data_i [312]),
    .B(\icache.data_mems_4__data_mem.data_o [56]),
    .S(_26527_),
    .Z(_04275_));
 MUX2_X1 _59432_ (.A(\icache.data_set_select_mux.data_i [313]),
    .B(\icache.data_mems_4__data_mem.data_o [57]),
    .S(_26527_),
    .Z(_04276_));
 MUX2_X1 _59433_ (.A(\icache.data_set_select_mux.data_i [314]),
    .B(\icache.data_mems_4__data_mem.data_o [58]),
    .S(_26527_),
    .Z(_04277_));
 MUX2_X1 _59434_ (.A(\icache.addr_tv_r [1]),
    .B(\icache.vaddr_tl_r [1]),
    .S(_26527_),
    .Z(_03969_));
 MUX2_X1 _59435_ (.A(\icache.data_set_select_mux.data_i [117]),
    .B(\icache.data_mems_1__data_mem.data_o [53]),
    .S(_26527_),
    .Z(_04058_));
 MUX2_X1 _59436_ (.A(\icache.data_set_select_mux.data_i [118]),
    .B(\icache.data_mems_1__data_mem.data_o [54]),
    .S(_26527_),
    .Z(_04059_));
 MUX2_X1 _59437_ (.A(\icache.data_set_select_mux.data_i [119]),
    .B(\icache.data_mems_1__data_mem.data_o [55]),
    .S(_26527_),
    .Z(_04060_));
 MUX2_X1 _59438_ (.A(\icache.data_set_select_mux.data_i [120]),
    .B(\icache.data_mems_1__data_mem.data_o [56]),
    .S(_26527_),
    .Z(_04062_));
 BUF_X8 _59439_ (.A(_26521_),
    .Z(_26528_));
 MUX2_X1 _59440_ (.A(\icache.data_set_select_mux.data_i [121]),
    .B(\icache.data_mems_1__data_mem.data_o [57]),
    .S(_26528_),
    .Z(_04063_));
 MUX2_X1 _59441_ (.A(\icache.data_set_select_mux.data_i [122]),
    .B(\icache.data_mems_1__data_mem.data_o [58]),
    .S(_26528_),
    .Z(_04064_));
 MUX2_X1 _59442_ (.A(\icache.data_set_select_mux.data_i [123]),
    .B(\icache.data_mems_1__data_mem.data_o [59]),
    .S(_26528_),
    .Z(_04065_));
 MUX2_X1 _59443_ (.A(\icache.data_set_select_mux.data_i [124]),
    .B(\icache.data_mems_1__data_mem.data_o [60]),
    .S(_26528_),
    .Z(_04066_));
 MUX2_X1 _59444_ (.A(\icache.data_set_select_mux.data_i [125]),
    .B(\icache.data_mems_1__data_mem.data_o [61]),
    .S(_26528_),
    .Z(_04067_));
 MUX2_X1 _59445_ (.A(\icache.data_set_select_mux.data_i [126]),
    .B(\icache.data_mems_1__data_mem.data_o [62]),
    .S(_26528_),
    .Z(_04068_));
 MUX2_X1 _59446_ (.A(\icache.data_set_select_mux.data_i [127]),
    .B(\icache.data_mems_1__data_mem.data_o [63]),
    .S(_26528_),
    .Z(_04069_));
 MUX2_X1 _59447_ (.A(\icache.data_set_select_mux.data_i [128]),
    .B(\icache.data_mems_2__data_mem.data_o [0]),
    .S(_26528_),
    .Z(_04070_));
 MUX2_X1 _59448_ (.A(\icache.data_set_select_mux.data_i [129]),
    .B(\icache.data_mems_2__data_mem.data_o [1]),
    .S(_26528_),
    .Z(_04071_));
 MUX2_X1 _59449_ (.A(\icache.data_set_select_mux.data_i [130]),
    .B(\icache.data_mems_2__data_mem.data_o [2]),
    .S(_26528_),
    .Z(_04073_));
 BUF_X8 _59450_ (.A(_26521_),
    .Z(_26529_));
 MUX2_X1 _59451_ (.A(\icache.data_set_select_mux.data_i [131]),
    .B(\icache.data_mems_2__data_mem.data_o [3]),
    .S(_26529_),
    .Z(_04074_));
 MUX2_X1 _59452_ (.A(\icache.data_set_select_mux.data_i [132]),
    .B(\icache.data_mems_2__data_mem.data_o [4]),
    .S(_26529_),
    .Z(_04075_));
 MUX2_X1 _59453_ (.A(\icache.data_set_select_mux.data_i [133]),
    .B(\icache.data_mems_2__data_mem.data_o [5]),
    .S(_26529_),
    .Z(_04076_));
 MUX2_X1 _59454_ (.A(\icache.data_set_select_mux.data_i [134]),
    .B(\icache.data_mems_2__data_mem.data_o [6]),
    .S(_26529_),
    .Z(_04077_));
 MUX2_X1 _59455_ (.A(\icache.data_set_select_mux.data_i [135]),
    .B(\icache.data_mems_2__data_mem.data_o [7]),
    .S(_26529_),
    .Z(_04078_));
 MUX2_X1 _59456_ (.A(\icache.data_set_select_mux.data_i [136]),
    .B(\icache.data_mems_2__data_mem.data_o [8]),
    .S(_26529_),
    .Z(_04079_));
 MUX2_X1 _59457_ (.A(\icache.data_set_select_mux.data_i [137]),
    .B(\icache.data_mems_2__data_mem.data_o [9]),
    .S(_26529_),
    .Z(_04080_));
 MUX2_X1 _59458_ (.A(\icache.data_set_select_mux.data_i [138]),
    .B(\icache.data_mems_2__data_mem.data_o [10]),
    .S(_26529_),
    .Z(_04081_));
 MUX2_X1 _59459_ (.A(\icache.data_set_select_mux.data_i [139]),
    .B(\icache.data_mems_2__data_mem.data_o [11]),
    .S(_26529_),
    .Z(_04082_));
 MUX2_X1 _59460_ (.A(\icache.data_set_select_mux.data_i [140]),
    .B(\icache.data_mems_2__data_mem.data_o [12]),
    .S(_26529_),
    .Z(_04084_));
 BUF_X4 _59461_ (.A(_26521_),
    .Z(_26530_));
 MUX2_X1 _59462_ (.A(\icache.data_set_select_mux.data_i [141]),
    .B(\icache.data_mems_2__data_mem.data_o [13]),
    .S(_26530_),
    .Z(_04085_));
 MUX2_X1 _59463_ (.A(\icache.data_set_select_mux.data_i [142]),
    .B(\icache.data_mems_2__data_mem.data_o [14]),
    .S(_26530_),
    .Z(_04086_));
 MUX2_X1 _59464_ (.A(\icache.data_set_select_mux.data_i [143]),
    .B(\icache.data_mems_2__data_mem.data_o [15]),
    .S(_26530_),
    .Z(_04087_));
 MUX2_X1 _59465_ (.A(\icache.data_set_select_mux.data_i [144]),
    .B(\icache.data_mems_2__data_mem.data_o [16]),
    .S(_26530_),
    .Z(_04088_));
 MUX2_X1 _59466_ (.A(\icache.data_set_select_mux.data_i [145]),
    .B(\icache.data_mems_2__data_mem.data_o [17]),
    .S(_26530_),
    .Z(_04089_));
 MUX2_X1 _59467_ (.A(\icache.data_set_select_mux.data_i [146]),
    .B(\icache.data_mems_2__data_mem.data_o [18]),
    .S(_26530_),
    .Z(_04090_));
 MUX2_X1 _59468_ (.A(\icache.data_set_select_mux.data_i [147]),
    .B(\icache.data_mems_2__data_mem.data_o [19]),
    .S(_26530_),
    .Z(_04091_));
 MUX2_X1 _59469_ (.A(\icache.data_set_select_mux.data_i [148]),
    .B(\icache.data_mems_2__data_mem.data_o [20]),
    .S(_26530_),
    .Z(_04092_));
 MUX2_X1 _59470_ (.A(\icache.data_set_select_mux.data_i [149]),
    .B(\icache.data_mems_2__data_mem.data_o [21]),
    .S(_26530_),
    .Z(_04093_));
 MUX2_X1 _59471_ (.A(\icache.data_set_select_mux.data_i [150]),
    .B(\icache.data_mems_2__data_mem.data_o [22]),
    .S(_26530_),
    .Z(_04095_));
 BUF_X4 _59472_ (.A(_26521_),
    .Z(_26531_));
 MUX2_X1 _59473_ (.A(\icache.data_set_select_mux.data_i [151]),
    .B(\icache.data_mems_2__data_mem.data_o [23]),
    .S(_26531_),
    .Z(_04096_));
 MUX2_X1 _59474_ (.A(\icache.data_set_select_mux.data_i [152]),
    .B(\icache.data_mems_2__data_mem.data_o [24]),
    .S(_26531_),
    .Z(_04097_));
 MUX2_X1 _59475_ (.A(\icache.data_set_select_mux.data_i [153]),
    .B(\icache.data_mems_2__data_mem.data_o [25]),
    .S(_26531_),
    .Z(_04098_));
 MUX2_X1 _59476_ (.A(\icache.data_set_select_mux.data_i [154]),
    .B(\icache.data_mems_2__data_mem.data_o [26]),
    .S(_26531_),
    .Z(_04099_));
 MUX2_X1 _59477_ (.A(\icache.data_set_select_mux.data_i [155]),
    .B(\icache.data_mems_2__data_mem.data_o [27]),
    .S(_26531_),
    .Z(_04100_));
 MUX2_X1 _59478_ (.A(\icache.data_set_select_mux.data_i [156]),
    .B(\icache.data_mems_2__data_mem.data_o [28]),
    .S(_26531_),
    .Z(_04101_));
 MUX2_X1 _59479_ (.A(\icache.data_set_select_mux.data_i [157]),
    .B(\icache.data_mems_2__data_mem.data_o [29]),
    .S(_26531_),
    .Z(_04102_));
 MUX2_X1 _59480_ (.A(\icache.data_set_select_mux.data_i [158]),
    .B(\icache.data_mems_2__data_mem.data_o [30]),
    .S(_26531_),
    .Z(_04103_));
 MUX2_X1 _59481_ (.A(\icache.data_set_select_mux.data_i [159]),
    .B(\icache.data_mems_2__data_mem.data_o [31]),
    .S(_26531_),
    .Z(_04104_));
 MUX2_X1 _59482_ (.A(\icache.data_set_select_mux.data_i [160]),
    .B(\icache.data_mems_2__data_mem.data_o [32]),
    .S(_26531_),
    .Z(_04106_));
 BUF_X8 _59483_ (.A(_26473_),
    .Z(_26532_));
 BUF_X4 _59484_ (.A(_26532_),
    .Z(_26533_));
 MUX2_X1 _59485_ (.A(\icache.data_set_select_mux.data_i [161]),
    .B(\icache.data_mems_2__data_mem.data_o [33]),
    .S(_26533_),
    .Z(_04107_));
 MUX2_X1 _59486_ (.A(\icache.data_set_select_mux.data_i [162]),
    .B(\icache.data_mems_2__data_mem.data_o [34]),
    .S(_26533_),
    .Z(_04108_));
 MUX2_X1 _59487_ (.A(\icache.data_set_select_mux.data_i [163]),
    .B(\icache.data_mems_2__data_mem.data_o [35]),
    .S(_26533_),
    .Z(_04109_));
 MUX2_X1 _59488_ (.A(\icache.data_set_select_mux.data_i [164]),
    .B(\icache.data_mems_2__data_mem.data_o [36]),
    .S(_26533_),
    .Z(_04110_));
 MUX2_X1 _59489_ (.A(\icache.data_set_select_mux.data_i [165]),
    .B(\icache.data_mems_2__data_mem.data_o [37]),
    .S(_26533_),
    .Z(_04111_));
 MUX2_X1 _59490_ (.A(\icache.data_set_select_mux.data_i [166]),
    .B(\icache.data_mems_2__data_mem.data_o [38]),
    .S(_26533_),
    .Z(_04112_));
 MUX2_X1 _59491_ (.A(\icache.data_set_select_mux.data_i [167]),
    .B(\icache.data_mems_2__data_mem.data_o [39]),
    .S(_26533_),
    .Z(_04113_));
 MUX2_X1 _59492_ (.A(\icache.data_set_select_mux.data_i [168]),
    .B(\icache.data_mems_2__data_mem.data_o [40]),
    .S(_26533_),
    .Z(_04114_));
 MUX2_X1 _59493_ (.A(\icache.data_set_select_mux.data_i [169]),
    .B(\icache.data_mems_2__data_mem.data_o [41]),
    .S(_26533_),
    .Z(_04115_));
 MUX2_X1 _59494_ (.A(\icache.data_set_select_mux.data_i [170]),
    .B(\icache.data_mems_2__data_mem.data_o [42]),
    .S(_26533_),
    .Z(_04117_));
 BUF_X4 _59495_ (.A(_26532_),
    .Z(_26534_));
 MUX2_X1 _59496_ (.A(\icache.data_set_select_mux.data_i [171]),
    .B(\icache.data_mems_2__data_mem.data_o [43]),
    .S(_26534_),
    .Z(_04118_));
 MUX2_X1 _59497_ (.A(\icache.data_set_select_mux.data_i [172]),
    .B(\icache.data_mems_2__data_mem.data_o [44]),
    .S(_26534_),
    .Z(_04119_));
 MUX2_X1 _59498_ (.A(\icache.data_set_select_mux.data_i [173]),
    .B(\icache.data_mems_2__data_mem.data_o [45]),
    .S(_26534_),
    .Z(_04120_));
 MUX2_X1 _59499_ (.A(\icache.data_set_select_mux.data_i [174]),
    .B(\icache.data_mems_2__data_mem.data_o [46]),
    .S(_26534_),
    .Z(_04121_));
 MUX2_X1 _59500_ (.A(\icache.data_set_select_mux.data_i [175]),
    .B(\icache.data_mems_2__data_mem.data_o [47]),
    .S(_26534_),
    .Z(_04122_));
 MUX2_X1 _59501_ (.A(\icache.data_set_select_mux.data_i [176]),
    .B(\icache.data_mems_2__data_mem.data_o [48]),
    .S(_26534_),
    .Z(_04123_));
 MUX2_X1 _59502_ (.A(\icache.data_set_select_mux.data_i [177]),
    .B(\icache.data_mems_2__data_mem.data_o [49]),
    .S(_26534_),
    .Z(_04124_));
 MUX2_X1 _59503_ (.A(\icache.data_set_select_mux.data_i [178]),
    .B(\icache.data_mems_2__data_mem.data_o [50]),
    .S(_26534_),
    .Z(_04125_));
 MUX2_X1 _59504_ (.A(\icache.data_set_select_mux.data_i [179]),
    .B(\icache.data_mems_2__data_mem.data_o [51]),
    .S(_26534_),
    .Z(_04126_));
 MUX2_X1 _59505_ (.A(\icache.data_set_select_mux.data_i [180]),
    .B(\icache.data_mems_2__data_mem.data_o [52]),
    .S(_26534_),
    .Z(_04128_));
 BUF_X8 _59506_ (.A(_26532_),
    .Z(_26535_));
 MUX2_X1 _59507_ (.A(\icache.data_set_select_mux.data_i [181]),
    .B(\icache.data_mems_2__data_mem.data_o [53]),
    .S(_26535_),
    .Z(_04129_));
 MUX2_X1 _59508_ (.A(\icache.data_set_select_mux.data_i [182]),
    .B(\icache.data_mems_2__data_mem.data_o [54]),
    .S(_26535_),
    .Z(_04130_));
 MUX2_X1 _59509_ (.A(\icache.data_set_select_mux.data_i [183]),
    .B(\icache.data_mems_2__data_mem.data_o [55]),
    .S(_26535_),
    .Z(_04131_));
 MUX2_X1 _59510_ (.A(\icache.data_set_select_mux.data_i [184]),
    .B(\icache.data_mems_2__data_mem.data_o [56]),
    .S(_26535_),
    .Z(_04132_));
 MUX2_X1 _59511_ (.A(\icache.data_set_select_mux.data_i [185]),
    .B(\icache.data_mems_2__data_mem.data_o [57]),
    .S(_26535_),
    .Z(_04133_));
 MUX2_X1 _59512_ (.A(\icache.data_set_select_mux.data_i [186]),
    .B(\icache.data_mems_2__data_mem.data_o [58]),
    .S(_26535_),
    .Z(_04134_));
 MUX2_X1 _59513_ (.A(\icache.data_set_select_mux.data_i [187]),
    .B(\icache.data_mems_2__data_mem.data_o [59]),
    .S(_26535_),
    .Z(_04135_));
 MUX2_X1 _59514_ (.A(\icache.data_set_select_mux.data_i [188]),
    .B(\icache.data_mems_2__data_mem.data_o [60]),
    .S(_26535_),
    .Z(_04136_));
 MUX2_X1 _59515_ (.A(\icache.data_set_select_mux.data_i [189]),
    .B(\icache.data_mems_2__data_mem.data_o [61]),
    .S(_26535_),
    .Z(_04137_));
 MUX2_X1 _59516_ (.A(\icache.data_set_select_mux.data_i [190]),
    .B(\icache.data_mems_2__data_mem.data_o [62]),
    .S(_26535_),
    .Z(_04139_));
 BUF_X8 _59517_ (.A(_26532_),
    .Z(_26536_));
 MUX2_X1 _59518_ (.A(\icache.data_set_select_mux.data_i [191]),
    .B(\icache.data_mems_2__data_mem.data_o [63]),
    .S(_26536_),
    .Z(_04140_));
 MUX2_X1 _59519_ (.A(\icache.data_set_select_mux.data_i [192]),
    .B(\icache.data_mems_3__data_mem.data_o [0]),
    .S(_26536_),
    .Z(_04141_));
 MUX2_X1 _59520_ (.A(\icache.data_set_select_mux.data_i [193]),
    .B(\icache.data_mems_3__data_mem.data_o [1]),
    .S(_26536_),
    .Z(_04142_));
 MUX2_X1 _59521_ (.A(\icache.data_set_select_mux.data_i [194]),
    .B(\icache.data_mems_3__data_mem.data_o [2]),
    .S(_26536_),
    .Z(_04143_));
 MUX2_X1 _59522_ (.A(\icache.data_set_select_mux.data_i [195]),
    .B(\icache.data_mems_3__data_mem.data_o [3]),
    .S(_26536_),
    .Z(_04144_));
 MUX2_X1 _59523_ (.A(\icache.data_set_select_mux.data_i [196]),
    .B(\icache.data_mems_3__data_mem.data_o [4]),
    .S(_26536_),
    .Z(_04145_));
 MUX2_X1 _59524_ (.A(\icache.data_set_select_mux.data_i [197]),
    .B(\icache.data_mems_3__data_mem.data_o [5]),
    .S(_26536_),
    .Z(_04146_));
 MUX2_X1 _59525_ (.A(\icache.data_set_select_mux.data_i [198]),
    .B(\icache.data_mems_3__data_mem.data_o [6]),
    .S(_26536_),
    .Z(_04147_));
 MUX2_X1 _59526_ (.A(\icache.data_set_select_mux.data_i [199]),
    .B(\icache.data_mems_3__data_mem.data_o [7]),
    .S(_26536_),
    .Z(_04148_));
 MUX2_X1 _59527_ (.A(\icache.data_set_select_mux.data_i [200]),
    .B(\icache.data_mems_3__data_mem.data_o [8]),
    .S(_26536_),
    .Z(_04151_));
 BUF_X4 _59528_ (.A(_26532_),
    .Z(_26537_));
 MUX2_X1 _59529_ (.A(\icache.data_set_select_mux.data_i [201]),
    .B(\icache.data_mems_3__data_mem.data_o [9]),
    .S(_26537_),
    .Z(_04152_));
 MUX2_X1 _59530_ (.A(\icache.data_set_select_mux.data_i [202]),
    .B(\icache.data_mems_3__data_mem.data_o [10]),
    .S(_26537_),
    .Z(_04153_));
 MUX2_X1 _59531_ (.A(\icache.data_set_select_mux.data_i [203]),
    .B(\icache.data_mems_3__data_mem.data_o [11]),
    .S(_26537_),
    .Z(_04154_));
 MUX2_X1 _59532_ (.A(\icache.data_set_select_mux.data_i [204]),
    .B(\icache.data_mems_3__data_mem.data_o [12]),
    .S(_26537_),
    .Z(_04155_));
 MUX2_X1 _59533_ (.A(\icache.data_set_select_mux.data_i [205]),
    .B(\icache.data_mems_3__data_mem.data_o [13]),
    .S(_26537_),
    .Z(_04156_));
 MUX2_X1 _59534_ (.A(\icache.data_set_select_mux.data_i [206]),
    .B(\icache.data_mems_3__data_mem.data_o [14]),
    .S(_26537_),
    .Z(_04157_));
 MUX2_X1 _59535_ (.A(\icache.data_set_select_mux.data_i [207]),
    .B(\icache.data_mems_3__data_mem.data_o [15]),
    .S(_26537_),
    .Z(_04158_));
 MUX2_X1 _59536_ (.A(\icache.data_set_select_mux.data_i [208]),
    .B(\icache.data_mems_3__data_mem.data_o [16]),
    .S(_26537_),
    .Z(_04159_));
 MUX2_X1 _59537_ (.A(\icache.data_set_select_mux.data_i [209]),
    .B(\icache.data_mems_3__data_mem.data_o [17]),
    .S(_26537_),
    .Z(_04160_));
 MUX2_X1 _59538_ (.A(\icache.data_set_select_mux.data_i [210]),
    .B(\icache.data_mems_3__data_mem.data_o [18]),
    .S(_26537_),
    .Z(_04162_));
 BUF_X8 _59539_ (.A(_26532_),
    .Z(_26538_));
 MUX2_X1 _59540_ (.A(\icache.data_set_select_mux.data_i [211]),
    .B(\icache.data_mems_3__data_mem.data_o [19]),
    .S(_26538_),
    .Z(_04163_));
 MUX2_X1 _59541_ (.A(\icache.data_set_select_mux.data_i [212]),
    .B(\icache.data_mems_3__data_mem.data_o [20]),
    .S(_26538_),
    .Z(_04164_));
 MUX2_X1 _59542_ (.A(\icache.data_set_select_mux.data_i [213]),
    .B(\icache.data_mems_3__data_mem.data_o [21]),
    .S(_26538_),
    .Z(_04165_));
 MUX2_X1 _59543_ (.A(\icache.data_set_select_mux.data_i [214]),
    .B(\icache.data_mems_3__data_mem.data_o [22]),
    .S(_26538_),
    .Z(_04166_));
 MUX2_X1 _59544_ (.A(\icache.data_set_select_mux.data_i [215]),
    .B(\icache.data_mems_3__data_mem.data_o [23]),
    .S(_26538_),
    .Z(_04167_));
 OAI21_X1 _59545_ (.A(_26437_),
    .B1(_09039_),
    .B2(\icache.N29 ),
    .ZN(_03980_));
 MUX2_X1 _59546_ (.A(\icache.data_set_select_mux.data_i [18]),
    .B(\icache.data_mems_0__data_mem.data_o [18]),
    .S(_26538_),
    .Z(_04138_));
 MUX2_X1 _59547_ (.A(\icache.data_set_select_mux.data_i [19]),
    .B(\icache.data_mems_0__data_mem.data_o [19]),
    .S(_26538_),
    .Z(_04149_));
 MUX2_X1 _59548_ (.A(\icache.data_set_select_mux.data_i [20]),
    .B(\icache.data_mems_0__data_mem.data_o [20]),
    .S(_26538_),
    .Z(_04161_));
 MUX2_X1 _59549_ (.A(\icache.data_set_select_mux.data_i [21]),
    .B(\icache.data_mems_0__data_mem.data_o [21]),
    .S(_26538_),
    .Z(_04172_));
 MUX2_X1 _59550_ (.A(\icache.data_set_select_mux.data_i [22]),
    .B(\icache.data_mems_0__data_mem.data_o [22]),
    .S(_26538_),
    .Z(_04183_));
 BUF_X8 _59551_ (.A(_26532_),
    .Z(_26539_));
 MUX2_X1 _59552_ (.A(\icache.data_set_select_mux.data_i [23]),
    .B(\icache.data_mems_0__data_mem.data_o [23]),
    .S(_26539_),
    .Z(_04194_));
 MUX2_X1 _59553_ (.A(\icache.data_set_select_mux.data_i [24]),
    .B(\icache.data_mems_0__data_mem.data_o [24]),
    .S(_26539_),
    .Z(_04205_));
 MUX2_X1 _59554_ (.A(\icache.data_set_select_mux.data_i [25]),
    .B(\icache.data_mems_0__data_mem.data_o [25]),
    .S(_26539_),
    .Z(_04216_));
 MUX2_X1 _59555_ (.A(\icache.data_set_select_mux.data_i [26]),
    .B(\icache.data_mems_0__data_mem.data_o [26]),
    .S(_26539_),
    .Z(_04227_));
 MUX2_X1 _59556_ (.A(\icache.data_set_select_mux.data_i [27]),
    .B(\icache.data_mems_0__data_mem.data_o [27]),
    .S(_26539_),
    .Z(_04238_));
 MUX2_X1 _59557_ (.A(\icache.data_set_select_mux.data_i [28]),
    .B(\icache.data_mems_0__data_mem.data_o [28]),
    .S(_26539_),
    .Z(_04249_));
 MUX2_X1 _59558_ (.A(\icache.data_set_select_mux.data_i [29]),
    .B(\icache.data_mems_0__data_mem.data_o [29]),
    .S(_26539_),
    .Z(_04260_));
 MUX2_X1 _59559_ (.A(\icache.data_set_select_mux.data_i [30]),
    .B(\icache.data_mems_0__data_mem.data_o [30]),
    .S(_26539_),
    .Z(_04272_));
 MUX2_X1 _59560_ (.A(\icache.data_set_select_mux.data_i [31]),
    .B(\icache.data_mems_0__data_mem.data_o [31]),
    .S(_26539_),
    .Z(_04283_));
 MUX2_X1 _59561_ (.A(\icache.data_set_select_mux.data_i [32]),
    .B(\icache.data_mems_0__data_mem.data_o [32]),
    .S(_26539_),
    .Z(_04294_));
 BUF_X4 _59562_ (.A(_26532_),
    .Z(_26540_));
 MUX2_X1 _59563_ (.A(\icache.data_set_select_mux.data_i [33]),
    .B(\icache.data_mems_0__data_mem.data_o [33]),
    .S(_26540_),
    .Z(_04305_));
 MUX2_X1 _59564_ (.A(\icache.data_set_select_mux.data_i [34]),
    .B(\icache.data_mems_0__data_mem.data_o [34]),
    .S(_26540_),
    .Z(_04316_));
 MUX2_X1 _59565_ (.A(\icache.data_set_select_mux.data_i [35]),
    .B(\icache.data_mems_0__data_mem.data_o [35]),
    .S(_26540_),
    .Z(_04327_));
 MUX2_X1 _59566_ (.A(\icache.data_set_select_mux.data_i [36]),
    .B(\icache.data_mems_0__data_mem.data_o [36]),
    .S(_26540_),
    .Z(_04338_));
 MUX2_X1 _59567_ (.A(\icache.data_set_select_mux.data_i [37]),
    .B(\icache.data_mems_0__data_mem.data_o [37]),
    .S(_26540_),
    .Z(_04349_));
 MUX2_X1 _59568_ (.A(\icache.data_set_select_mux.data_i [38]),
    .B(\icache.data_mems_0__data_mem.data_o [38]),
    .S(_26540_),
    .Z(_04360_));
 MUX2_X1 _59569_ (.A(\icache.data_set_select_mux.data_i [39]),
    .B(\icache.data_mems_0__data_mem.data_o [39]),
    .S(_26540_),
    .Z(_04371_));
 MUX2_X1 _59570_ (.A(\icache.data_set_select_mux.data_i [40]),
    .B(\icache.data_mems_0__data_mem.data_o [40]),
    .S(_26540_),
    .Z(_04383_));
 MUX2_X1 _59571_ (.A(\icache.data_set_select_mux.data_i [41]),
    .B(\icache.data_mems_0__data_mem.data_o [41]),
    .S(_26540_),
    .Z(_04394_));
 MUX2_X1 _59572_ (.A(\icache.data_set_select_mux.data_i [42]),
    .B(\icache.data_mems_0__data_mem.data_o [42]),
    .S(_26540_),
    .Z(_04405_));
 BUF_X4 _59573_ (.A(_26532_),
    .Z(_26541_));
 MUX2_X1 _59574_ (.A(\icache.data_set_select_mux.data_i [43]),
    .B(\icache.data_mems_0__data_mem.data_o [43]),
    .S(_26541_),
    .Z(_04416_));
 MUX2_X1 _59575_ (.A(\icache.data_set_select_mux.data_i [44]),
    .B(\icache.data_mems_0__data_mem.data_o [44]),
    .S(_26541_),
    .Z(_04427_));
 MUX2_X1 _59576_ (.A(\icache.data_set_select_mux.data_i [45]),
    .B(\icache.data_mems_0__data_mem.data_o [45]),
    .S(_26541_),
    .Z(_04438_));
 MUX2_X1 _59577_ (.A(\icache.data_set_select_mux.data_i [46]),
    .B(\icache.data_mems_0__data_mem.data_o [46]),
    .S(_26541_),
    .Z(_04449_));
 MUX2_X1 _59578_ (.A(\icache.data_set_select_mux.data_i [47]),
    .B(\icache.data_mems_0__data_mem.data_o [47]),
    .S(_26541_),
    .Z(_04460_));
 MUX2_X1 _59579_ (.A(\icache.data_set_select_mux.data_i [48]),
    .B(\icache.data_mems_0__data_mem.data_o [48]),
    .S(_26541_),
    .Z(_04471_));
 MUX2_X1 _59580_ (.A(\icache.data_set_select_mux.data_i [49]),
    .B(\icache.data_mems_0__data_mem.data_o [49]),
    .S(_26541_),
    .Z(_04482_));
 MUX2_X1 _59581_ (.A(\icache.data_set_select_mux.data_i [50]),
    .B(\icache.data_mems_0__data_mem.data_o [50]),
    .S(_26541_),
    .Z(_04494_));
 MUX2_X1 _59582_ (.A(\icache.data_set_select_mux.data_i [51]),
    .B(\icache.data_mems_0__data_mem.data_o [51]),
    .S(_26541_),
    .Z(_04497_));
 MUX2_X1 _59583_ (.A(\icache.data_set_select_mux.data_i [52]),
    .B(\icache.data_mems_0__data_mem.data_o [52]),
    .S(_26541_),
    .Z(_04498_));
 BUF_X8 _59584_ (.A(_26532_),
    .Z(_26542_));
 MUX2_X1 _59585_ (.A(\icache.data_set_select_mux.data_i [53]),
    .B(\icache.data_mems_0__data_mem.data_o [53]),
    .S(_26542_),
    .Z(_04499_));
 MUX2_X1 _59586_ (.A(\icache.data_set_select_mux.data_i [54]),
    .B(\icache.data_mems_0__data_mem.data_o [54]),
    .S(_26542_),
    .Z(_04500_));
 MUX2_X1 _59587_ (.A(\icache.data_set_select_mux.data_i [55]),
    .B(\icache.data_mems_0__data_mem.data_o [55]),
    .S(_26542_),
    .Z(_04501_));
 MUX2_X1 _59588_ (.A(\icache.data_set_select_mux.data_i [56]),
    .B(\icache.data_mems_0__data_mem.data_o [56]),
    .S(_26542_),
    .Z(_04502_));
 MUX2_X1 _59589_ (.A(\icache.data_set_select_mux.data_i [57]),
    .B(\icache.data_mems_0__data_mem.data_o [57]),
    .S(_26542_),
    .Z(_04503_));
 MUX2_X1 _59590_ (.A(\icache.data_set_select_mux.data_i [58]),
    .B(\icache.data_mems_0__data_mem.data_o [58]),
    .S(_26542_),
    .Z(_04504_));
 MUX2_X1 _59591_ (.A(\icache.data_set_select_mux.data_i [59]),
    .B(\icache.data_mems_0__data_mem.data_o [59]),
    .S(_26542_),
    .Z(_04505_));
 MUX2_X1 _59592_ (.A(\icache.data_set_select_mux.data_i [60]),
    .B(\icache.data_mems_0__data_mem.data_o [60]),
    .S(_26542_),
    .Z(_04507_));
 MUX2_X1 _59593_ (.A(\icache.data_set_select_mux.data_i [61]),
    .B(\icache.data_mems_0__data_mem.data_o [61]),
    .S(_26542_),
    .Z(_04508_));
 MUX2_X1 _59594_ (.A(\icache.data_set_select_mux.data_i [62]),
    .B(\icache.data_mems_0__data_mem.data_o [62]),
    .S(_26542_),
    .Z(_04509_));
 BUF_X32 _59595_ (.A(_08517_),
    .Z(_26543_));
 BUF_X4 _59596_ (.A(_26543_),
    .Z(_26544_));
 MUX2_X1 _59597_ (.A(\icache.data_set_select_mux.data_i [63]),
    .B(\icache.data_mems_0__data_mem.data_o [63]),
    .S(_26544_),
    .Z(_04510_));
 MUX2_X1 _59598_ (.A(\icache.data_set_select_mux.data_i [64]),
    .B(\icache.data_mems_1__data_mem.data_o [0]),
    .S(_26544_),
    .Z(_04511_));
 MUX2_X1 _59599_ (.A(\icache.data_set_select_mux.data_i [65]),
    .B(\icache.data_mems_1__data_mem.data_o [1]),
    .S(_26544_),
    .Z(_04512_));
 MUX2_X1 _59600_ (.A(\icache.data_set_select_mux.data_i [66]),
    .B(\icache.data_mems_1__data_mem.data_o [2]),
    .S(_26544_),
    .Z(_04513_));
 MUX2_X1 _59601_ (.A(\icache.data_set_select_mux.data_i [67]),
    .B(\icache.data_mems_1__data_mem.data_o [3]),
    .S(_26544_),
    .Z(_04514_));
 MUX2_X1 _59602_ (.A(\icache.data_set_select_mux.data_i [68]),
    .B(\icache.data_mems_1__data_mem.data_o [4]),
    .S(_26544_),
    .Z(_04515_));
 MUX2_X1 _59603_ (.A(\icache.data_set_select_mux.data_i [69]),
    .B(\icache.data_mems_1__data_mem.data_o [5]),
    .S(_26544_),
    .Z(_04516_));
 MUX2_X1 _59604_ (.A(\icache.data_set_select_mux.data_i [70]),
    .B(\icache.data_mems_1__data_mem.data_o [6]),
    .S(_26544_),
    .Z(_04518_));
 MUX2_X1 _59605_ (.A(\icache.data_set_select_mux.data_i [71]),
    .B(\icache.data_mems_1__data_mem.data_o [7]),
    .S(_26544_),
    .Z(_04519_));
 MUX2_X1 _59606_ (.A(\icache.data_set_select_mux.data_i [72]),
    .B(\icache.data_mems_1__data_mem.data_o [8]),
    .S(_26544_),
    .Z(_04520_));
 BUF_X4 _59607_ (.A(_26543_),
    .Z(_26545_));
 MUX2_X1 _59608_ (.A(\icache.data_set_select_mux.data_i [73]),
    .B(\icache.data_mems_1__data_mem.data_o [9]),
    .S(_26545_),
    .Z(_04521_));
 MUX2_X1 _59609_ (.A(\icache.data_set_select_mux.data_i [74]),
    .B(\icache.data_mems_1__data_mem.data_o [10]),
    .S(_26545_),
    .Z(_04522_));
 MUX2_X1 _59610_ (.A(\icache.data_set_select_mux.data_i [75]),
    .B(\icache.data_mems_1__data_mem.data_o [11]),
    .S(_26545_),
    .Z(_04523_));
 MUX2_X1 _59611_ (.A(\icache.data_set_select_mux.data_i [76]),
    .B(\icache.data_mems_1__data_mem.data_o [12]),
    .S(_26545_),
    .Z(_04524_));
 MUX2_X1 _59612_ (.A(\icache.data_set_select_mux.data_i [77]),
    .B(\icache.data_mems_1__data_mem.data_o [13]),
    .S(_26545_),
    .Z(_04525_));
 MUX2_X1 _59613_ (.A(\icache.data_set_select_mux.data_i [78]),
    .B(\icache.data_mems_1__data_mem.data_o [14]),
    .S(_26545_),
    .Z(_04526_));
 MUX2_X1 _59614_ (.A(\icache.data_set_select_mux.data_i [79]),
    .B(\icache.data_mems_1__data_mem.data_o [15]),
    .S(_26545_),
    .Z(_04527_));
 MUX2_X1 _59615_ (.A(\icache.data_set_select_mux.data_i [80]),
    .B(\icache.data_mems_1__data_mem.data_o [16]),
    .S(_26545_),
    .Z(_04529_));
 MUX2_X1 _59616_ (.A(\icache.data_set_select_mux.data_i [81]),
    .B(\icache.data_mems_1__data_mem.data_o [17]),
    .S(_26545_),
    .Z(_04530_));
 MUX2_X1 _59617_ (.A(\icache.data_set_select_mux.data_i [82]),
    .B(\icache.data_mems_1__data_mem.data_o [18]),
    .S(_26545_),
    .Z(_04531_));
 BUF_X4 _59618_ (.A(_26543_),
    .Z(_26546_));
 MUX2_X1 _59619_ (.A(\icache.data_set_select_mux.data_i [83]),
    .B(\icache.data_mems_1__data_mem.data_o [19]),
    .S(_26546_),
    .Z(_04532_));
 MUX2_X1 _59620_ (.A(\icache.data_set_select_mux.data_i [84]),
    .B(\icache.data_mems_1__data_mem.data_o [20]),
    .S(_26546_),
    .Z(_04533_));
 MUX2_X1 _59621_ (.A(\icache.data_set_select_mux.data_i [85]),
    .B(\icache.data_mems_1__data_mem.data_o [21]),
    .S(_26546_),
    .Z(_04534_));
 MUX2_X1 _59622_ (.A(\icache.data_set_select_mux.data_i [86]),
    .B(\icache.data_mems_1__data_mem.data_o [22]),
    .S(_26546_),
    .Z(_04535_));
 MUX2_X1 _59623_ (.A(\icache.data_set_select_mux.data_i [87]),
    .B(\icache.data_mems_1__data_mem.data_o [23]),
    .S(_26546_),
    .Z(_04536_));
 MUX2_X1 _59624_ (.A(\icache.data_set_select_mux.data_i [88]),
    .B(\icache.data_mems_1__data_mem.data_o [24]),
    .S(_26546_),
    .Z(_04537_));
 MUX2_X1 _59625_ (.A(\icache.data_set_select_mux.data_i [89]),
    .B(\icache.data_mems_1__data_mem.data_o [25]),
    .S(_26546_),
    .Z(_04538_));
 MUX2_X1 _59626_ (.A(\icache.data_set_select_mux.data_i [90]),
    .B(\icache.data_mems_1__data_mem.data_o [26]),
    .S(_26546_),
    .Z(_04540_));
 MUX2_X1 _59627_ (.A(\icache.data_set_select_mux.data_i [91]),
    .B(\icache.data_mems_1__data_mem.data_o [27]),
    .S(_26546_),
    .Z(_04541_));
 MUX2_X1 _59628_ (.A(\icache.data_set_select_mux.data_i [92]),
    .B(\icache.data_mems_1__data_mem.data_o [28]),
    .S(_26546_),
    .Z(_04542_));
 BUF_X8 _59629_ (.A(_26543_),
    .Z(_26547_));
 MUX2_X1 _59630_ (.A(\icache.data_set_select_mux.data_i [93]),
    .B(\icache.data_mems_1__data_mem.data_o [29]),
    .S(_26547_),
    .Z(_04543_));
 MUX2_X1 _59631_ (.A(\icache.data_set_select_mux.data_i [94]),
    .B(\icache.data_mems_1__data_mem.data_o [30]),
    .S(_26547_),
    .Z(_04544_));
 MUX2_X1 _59632_ (.A(\icache.data_set_select_mux.data_i [95]),
    .B(\icache.data_mems_1__data_mem.data_o [31]),
    .S(_26547_),
    .Z(_04545_));
 MUX2_X1 _59633_ (.A(\icache.data_set_select_mux.data_i [96]),
    .B(\icache.data_mems_1__data_mem.data_o [32]),
    .S(_26547_),
    .Z(_04546_));
 MUX2_X1 _59634_ (.A(\icache.data_set_select_mux.data_i [97]),
    .B(\icache.data_mems_1__data_mem.data_o [33]),
    .S(_26547_),
    .Z(_04547_));
 MUX2_X1 _59635_ (.A(\icache.data_set_select_mux.data_i [98]),
    .B(\icache.data_mems_1__data_mem.data_o [34]),
    .S(_26547_),
    .Z(_04548_));
 MUX2_X1 _59636_ (.A(\icache.data_set_select_mux.data_i [99]),
    .B(\icache.data_mems_1__data_mem.data_o [35]),
    .S(_26547_),
    .Z(_04549_));
 MUX2_X1 _59637_ (.A(\icache.data_set_select_mux.data_i [100]),
    .B(\icache.data_mems_1__data_mem.data_o [36]),
    .S(_26547_),
    .Z(_04040_));
 MUX2_X1 _59638_ (.A(\icache.data_set_select_mux.data_i [101]),
    .B(\icache.data_mems_1__data_mem.data_o [37]),
    .S(_26547_),
    .Z(_04041_));
 MUX2_X1 _59639_ (.A(\icache.data_set_select_mux.data_i [102]),
    .B(\icache.data_mems_1__data_mem.data_o [38]),
    .S(_26547_),
    .Z(_04042_));
 BUF_X8 _59640_ (.A(_26543_),
    .Z(_26548_));
 MUX2_X1 _59641_ (.A(\icache.data_set_select_mux.data_i [103]),
    .B(\icache.data_mems_1__data_mem.data_o [39]),
    .S(_26548_),
    .Z(_04043_));
 MUX2_X1 _59642_ (.A(\icache.data_set_select_mux.data_i [104]),
    .B(\icache.data_mems_1__data_mem.data_o [40]),
    .S(_26548_),
    .Z(_04044_));
 MUX2_X1 _59643_ (.A(\icache.data_set_select_mux.data_i [105]),
    .B(\icache.data_mems_1__data_mem.data_o [41]),
    .S(_26548_),
    .Z(_04045_));
 MUX2_X1 _59644_ (.A(\icache.data_set_select_mux.data_i [106]),
    .B(\icache.data_mems_1__data_mem.data_o [42]),
    .S(_26548_),
    .Z(_04046_));
 MUX2_X1 _59645_ (.A(\icache.data_set_select_mux.data_i [107]),
    .B(\icache.data_mems_1__data_mem.data_o [43]),
    .S(_26548_),
    .Z(_04047_));
 MUX2_X1 _59646_ (.A(\icache.data_set_select_mux.data_i [108]),
    .B(\icache.data_mems_1__data_mem.data_o [44]),
    .S(_26548_),
    .Z(_04048_));
 MUX2_X1 _59647_ (.A(\icache.data_set_select_mux.data_i [109]),
    .B(\icache.data_mems_1__data_mem.data_o [45]),
    .S(_26548_),
    .Z(_04049_));
 MUX2_X1 _59648_ (.A(\icache.data_set_select_mux.data_i [110]),
    .B(\icache.data_mems_1__data_mem.data_o [46]),
    .S(_26548_),
    .Z(_04051_));
 MUX2_X1 _59649_ (.A(\icache.data_set_select_mux.data_i [111]),
    .B(\icache.data_mems_1__data_mem.data_o [47]),
    .S(_26548_),
    .Z(_04052_));
 MUX2_X1 _59650_ (.A(\icache.data_set_select_mux.data_i [112]),
    .B(\icache.data_mems_1__data_mem.data_o [48]),
    .S(_26548_),
    .Z(_04053_));
 BUF_X16 _59651_ (.A(_26543_),
    .Z(_26549_));
 MUX2_X1 _59652_ (.A(\icache.data_set_select_mux.data_i [113]),
    .B(\icache.data_mems_1__data_mem.data_o [49]),
    .S(_26549_),
    .Z(_04054_));
 MUX2_X1 _59653_ (.A(\icache.data_set_select_mux.data_i [114]),
    .B(\icache.data_mems_1__data_mem.data_o [50]),
    .S(_26549_),
    .Z(_04055_));
 MUX2_X1 _59654_ (.A(\icache.data_set_select_mux.data_i [115]),
    .B(\icache.data_mems_1__data_mem.data_o [51]),
    .S(_26549_),
    .Z(_04056_));
 MUX2_X1 _59655_ (.A(\icache.data_set_select_mux.data_i [116]),
    .B(\icache.data_mems_1__data_mem.data_o [52]),
    .S(_26549_),
    .Z(_04057_));
 MUX2_X1 _59656_ (.A(\icache.addr_tv_r [3]),
    .B(\icache.vaddr_tl_r [3]),
    .S(_26549_),
    .Z(_03990_));
 MUX2_X1 _59657_ (.A(\icache.data_set_select_mux.data_i [0]),
    .B(\icache.data_mems_0__data_mem.data_o [0]),
    .S(_26549_),
    .Z(_04039_));
 MUX2_X1 _59658_ (.A(\icache.data_set_select_mux.data_i [1]),
    .B(\icache.data_mems_0__data_mem.data_o [1]),
    .S(_26549_),
    .Z(_04150_));
 MUX2_X1 _59659_ (.A(\icache.data_set_select_mux.data_i [2]),
    .B(\icache.data_mems_0__data_mem.data_o [2]),
    .S(_26549_),
    .Z(_04261_));
 MUX2_X1 _59660_ (.A(\icache.data_set_select_mux.data_i [3]),
    .B(\icache.data_mems_0__data_mem.data_o [3]),
    .S(_26549_),
    .Z(_04372_));
 MUX2_X1 _59661_ (.A(\icache.data_set_select_mux.data_i [4]),
    .B(\icache.data_mems_0__data_mem.data_o [4]),
    .S(_26549_),
    .Z(_04483_));
 BUF_X4 _59662_ (.A(_26543_),
    .Z(_26550_));
 MUX2_X1 _59663_ (.A(\icache.data_set_select_mux.data_i [5]),
    .B(\icache.data_mems_0__data_mem.data_o [5]),
    .S(_26550_),
    .Z(_04506_));
 MUX2_X1 _59664_ (.A(\icache.data_set_select_mux.data_i [6]),
    .B(\icache.data_mems_0__data_mem.data_o [6]),
    .S(_26550_),
    .Z(_04517_));
 MUX2_X1 _59665_ (.A(\icache.data_set_select_mux.data_i [7]),
    .B(\icache.data_mems_0__data_mem.data_o [7]),
    .S(_26550_),
    .Z(_04528_));
 MUX2_X1 _59666_ (.A(\icache.data_set_select_mux.data_i [8]),
    .B(\icache.data_mems_0__data_mem.data_o [8]),
    .S(_26550_),
    .Z(_04539_));
 MUX2_X1 _59667_ (.A(\icache.data_set_select_mux.data_i [9]),
    .B(\icache.data_mems_0__data_mem.data_o [9]),
    .S(_26550_),
    .Z(_04550_));
 MUX2_X1 _59668_ (.A(\icache.data_set_select_mux.data_i [10]),
    .B(\icache.data_mems_0__data_mem.data_o [10]),
    .S(_26550_),
    .Z(_04050_));
 MUX2_X1 _59669_ (.A(\icache.data_set_select_mux.data_i [11]),
    .B(\icache.data_mems_0__data_mem.data_o [11]),
    .S(_26550_),
    .Z(_04061_));
 MUX2_X1 _59670_ (.A(\icache.data_set_select_mux.data_i [12]),
    .B(\icache.data_mems_0__data_mem.data_o [12]),
    .S(_26550_),
    .Z(_04072_));
 MUX2_X1 _59671_ (.A(\icache.data_set_select_mux.data_i [13]),
    .B(\icache.data_mems_0__data_mem.data_o [13]),
    .S(_26550_),
    .Z(_04083_));
 MUX2_X1 _59672_ (.A(\icache.data_set_select_mux.data_i [14]),
    .B(\icache.data_mems_0__data_mem.data_o [14]),
    .S(_26550_),
    .Z(_04094_));
 BUF_X16 _59673_ (.A(_26543_),
    .Z(_26551_));
 MUX2_X1 _59674_ (.A(\icache.data_set_select_mux.data_i [15]),
    .B(\icache.data_mems_0__data_mem.data_o [15]),
    .S(_26551_),
    .Z(_04105_));
 MUX2_X1 _59675_ (.A(\icache.data_set_select_mux.data_i [16]),
    .B(\icache.data_mems_0__data_mem.data_o [16]),
    .S(_26551_),
    .Z(_04116_));
 MUX2_X1 _59676_ (.A(\icache.data_set_select_mux.data_i [17]),
    .B(\icache.data_mems_0__data_mem.data_o [17]),
    .S(_26551_),
    .Z(_04127_));
 MUX2_X1 _59677_ (.A(\icache.addr_tv_r [4]),
    .B(\icache.vaddr_tl_r [4]),
    .S(_26551_),
    .Z(_03991_));
 OAI21_X1 _59678_ (.A(_26438_),
    .B1(_09051_),
    .B2(_26436_),
    .ZN(_03992_));
 MUX2_X1 _59679_ (.A(net1335),
    .B(\icache.itlb_icache_data_resp_i [19]),
    .S(_26551_),
    .Z(_03982_));
 MUX2_X1 _59680_ (.A(_07133_),
    .B(\icache.itlb_icache_data_resp_i [20]),
    .S(_26551_),
    .Z(_03983_));
 MUX2_X1 _59681_ (.A(net1330),
    .B(\icache.itlb_icache_data_resp_i [21]),
    .S(_26551_),
    .Z(_03984_));
 MUX2_X1 _59682_ (.A(_07156_),
    .B(\icache.itlb_icache_data_resp_i [22]),
    .S(_26551_),
    .Z(_03985_));
 MUX2_X1 _59683_ (.A(net1325),
    .B(\icache.itlb_icache_data_resp_i [23]),
    .S(_26551_),
    .Z(_03986_));
 MUX2_X1 _59684_ (.A(_07092_),
    .B(\icache.itlb_icache_data_resp_i [24]),
    .S(_26551_),
    .Z(_03987_));
 BUF_X4 _59685_ (.A(_26543_),
    .Z(_26552_));
 MUX2_X1 _59686_ (.A(net1319),
    .B(\icache.itlb_icache_data_resp_i [25]),
    .S(_26552_),
    .Z(_03988_));
 MUX2_X1 _59687_ (.A(_07160_),
    .B(\icache.itlb_icache_data_resp_i [26]),
    .S(_26552_),
    .Z(_03989_));
 OAI21_X1 _59688_ (.A(_26439_),
    .B1(_07628_),
    .B2(_26436_),
    .ZN(_03993_));
 OAI21_X1 _59689_ (.A(_26440_),
    .B1(_07634_),
    .B2(_26436_),
    .ZN(_03994_));
 OAI21_X1 _59690_ (.A(_26441_),
    .B1(_07639_),
    .B2(_26436_),
    .ZN(_03995_));
 OAI21_X1 _59691_ (.A(_26442_),
    .B1(_07644_),
    .B2(_26436_),
    .ZN(_03996_));
 OAI21_X1 _59692_ (.A(_26443_),
    .B1(_07649_),
    .B2(_26436_),
    .ZN(_03959_));
 OAI21_X1 _59693_ (.A(_26444_),
    .B1(_07654_),
    .B2(_26436_),
    .ZN(_03960_));
 MUX2_X1 _59694_ (.A(_07193_),
    .B(\icache.itlb_icache_data_resp_i [0]),
    .S(_26552_),
    .Z(_03961_));
 MUX2_X1 _59695_ (.A(net1380),
    .B(\icache.itlb_icache_data_resp_i [1]),
    .S(_26552_),
    .Z(_03962_));
 MUX2_X2 _59696_ (.A(_07370_),
    .B(\icache.itlb_icache_data_resp_i [2]),
    .S(_26552_),
    .Z(_03963_));
 MUX2_X1 _59697_ (.A(_07186_),
    .B(\icache.itlb_icache_data_resp_i [3]),
    .S(_26552_),
    .Z(_03964_));
 MUX2_X1 _59698_ (.A(_07123_),
    .B(\icache.itlb_icache_data_resp_i [4]),
    .S(_26552_),
    .Z(_03965_));
 MUX2_X1 _59699_ (.A(net1369),
    .B(\icache.itlb_icache_data_resp_i [5]),
    .S(_26552_),
    .Z(_03966_));
 MUX2_X1 _59700_ (.A(_07113_),
    .B(\icache.itlb_icache_data_resp_i [6]),
    .S(_26552_),
    .Z(_03967_));
 MUX2_X1 _59701_ (.A(net1361),
    .B(\icache.itlb_icache_data_resp_i [7]),
    .S(_26552_),
    .Z(_03968_));
 BUF_X4 _59702_ (.A(_26543_),
    .Z(_26553_));
 MUX2_X1 _59703_ (.A(_07128_),
    .B(\icache.itlb_icache_data_resp_i [8]),
    .S(_26553_),
    .Z(_03970_));
 MUX2_X1 _59704_ (.A(net1356),
    .B(\icache.itlb_icache_data_resp_i [9]),
    .S(_26553_),
    .Z(_03971_));
 MUX2_X1 _59705_ (.A(_07118_),
    .B(\icache.itlb_icache_data_resp_i [10]),
    .S(_26553_),
    .Z(_03972_));
 MUX2_X1 _59706_ (.A(net1353),
    .B(\icache.itlb_icache_data_resp_i [11]),
    .S(_26553_),
    .Z(_03973_));
 MUX2_X1 _59707_ (.A(_07105_),
    .B(\icache.itlb_icache_data_resp_i [12]),
    .S(_26553_),
    .Z(_03974_));
 MUX2_X1 _59708_ (.A(_07135_),
    .B(\icache.itlb_icache_data_resp_i [13]),
    .S(_26553_),
    .Z(_03975_));
 MUX2_X1 _59709_ (.A(_07107_),
    .B(\icache.itlb_icache_data_resp_i [14]),
    .S(_26553_),
    .Z(_03976_));
 MUX2_X1 _59710_ (.A(_07190_),
    .B(\icache.itlb_icache_data_resp_i [15]),
    .S(_26553_),
    .Z(_03977_));
 MUX2_X1 _59711_ (.A(net1344),
    .B(\icache.itlb_icache_data_resp_i [16]),
    .S(_26553_),
    .Z(_03978_));
 MUX2_X1 _59712_ (.A(_07248_),
    .B(\icache.itlb_icache_data_resp_i [17]),
    .S(_26553_),
    .Z(_03979_));
 BUF_X16 _59713_ (.A(_08517_),
    .Z(_26554_));
 BUF_X4 _59714_ (.A(_26554_),
    .Z(_26555_));
 MUX2_X1 _59715_ (.A(_07130_),
    .B(\icache.itlb_icache_data_resp_i [18]),
    .S(_26555_),
    .Z(_03981_));
 MUX2_X1 _59716_ (.A(\icache.tag_tv_r [0]),
    .B(\icache.tag_mem.data_o [0]),
    .S(_26555_),
    .Z(_04567_));
 MUX2_X1 _59717_ (.A(\icache.tag_tv_r [1]),
    .B(\icache.tag_mem.data_o [1]),
    .S(_26555_),
    .Z(_04678_));
 MUX2_X1 _59718_ (.A(\icache.tag_tv_r [2]),
    .B(\icache.tag_mem.data_o [2]),
    .S(_26555_),
    .Z(_04705_));
 MUX2_X1 _59719_ (.A(\icache.tag_tv_r [3]),
    .B(\icache.tag_mem.data_o [3]),
    .S(_26555_),
    .Z(_04716_));
 MUX2_X1 _59720_ (.A(\icache.tag_tv_r [4]),
    .B(\icache.tag_mem.data_o [4]),
    .S(_26555_),
    .Z(_04727_));
 MUX2_X1 _59721_ (.A(\icache.tag_tv_r [5]),
    .B(\icache.tag_mem.data_o [5]),
    .S(_26555_),
    .Z(_04738_));
 MUX2_X1 _59722_ (.A(\icache.tag_tv_r [6]),
    .B(\icache.tag_mem.data_o [6]),
    .S(_26555_),
    .Z(_04749_));
 MUX2_X1 _59723_ (.A(\icache.tag_tv_r [7]),
    .B(\icache.tag_mem.data_o [7]),
    .S(_26555_),
    .Z(_04760_));
 MUX2_X1 _59724_ (.A(\icache.tag_tv_r [8]),
    .B(\icache.tag_mem.data_o [8]),
    .S(_26555_),
    .Z(_04771_));
 BUF_X4 _59725_ (.A(_26554_),
    .Z(_26556_));
 MUX2_X1 _59726_ (.A(\icache.tag_tv_r [9]),
    .B(\icache.tag_mem.data_o [9]),
    .S(_26556_),
    .Z(_04782_));
 MUX2_X1 _59727_ (.A(\icache.tag_tv_r [10]),
    .B(\icache.tag_mem.data_o [10]),
    .S(_26556_),
    .Z(_04578_));
 MUX2_X1 _59728_ (.A(\icache.tag_tv_r [11]),
    .B(\icache.tag_mem.data_o [11]),
    .S(_26556_),
    .Z(_04589_));
 MUX2_X1 _59729_ (.A(\icache.tag_tv_r [12]),
    .B(\icache.tag_mem.data_o [12]),
    .S(_26556_),
    .Z(_04600_));
 MUX2_X1 _59730_ (.A(\icache.tag_tv_r [13]),
    .B(\icache.tag_mem.data_o [13]),
    .S(_26556_),
    .Z(_04611_));
 MUX2_X1 _59731_ (.A(\icache.tag_tv_r [14]),
    .B(\icache.tag_mem.data_o [14]),
    .S(_26556_),
    .Z(_04622_));
 MUX2_X1 _59732_ (.A(\icache.tag_tv_r [15]),
    .B(\icache.tag_mem.data_o [15]),
    .S(_26556_),
    .Z(_04633_));
 MUX2_X1 _59733_ (.A(\icache.tag_tv_r [16]),
    .B(\icache.tag_mem.data_o [16]),
    .S(_26556_),
    .Z(_04644_));
 MUX2_X1 _59734_ (.A(\icache.tag_tv_r [17]),
    .B(\icache.tag_mem.data_o [17]),
    .S(_26556_),
    .Z(_04655_));
 MUX2_X1 _59735_ (.A(\icache.tag_tv_r [18]),
    .B(\icache.tag_mem.data_o [18]),
    .S(_26556_),
    .Z(_04666_));
 BUF_X8 _59736_ (.A(_26554_),
    .Z(_26557_));
 MUX2_X1 _59737_ (.A(\icache.tag_tv_r [19]),
    .B(\icache.tag_mem.data_o [19]),
    .S(_26557_),
    .Z(_04677_));
 MUX2_X1 _59738_ (.A(\icache.tag_tv_r [20]),
    .B(\icache.tag_mem.data_o [20]),
    .S(_26557_),
    .Z(_04689_));
 MUX2_X1 _59739_ (.A(\icache.tag_tv_r [21]),
    .B(\icache.tag_mem.data_o [21]),
    .S(_26557_),
    .Z(_04696_));
 MUX2_X1 _59740_ (.A(\icache.tag_tv_r [22]),
    .B(\icache.tag_mem.data_o [22]),
    .S(_26557_),
    .Z(_04697_));
 MUX2_X1 _59741_ (.A(\icache.tag_tv_r [23]),
    .B(\icache.tag_mem.data_o [23]),
    .S(_26557_),
    .Z(_04698_));
 MUX2_X1 _59742_ (.A(\icache.tag_tv_r [24]),
    .B(\icache.tag_mem.data_o [24]),
    .S(_26557_),
    .Z(_04699_));
 MUX2_X1 _59743_ (.A(\icache.tag_tv_r [25]),
    .B(\icache.tag_mem.data_o [25]),
    .S(_26557_),
    .Z(_04700_));
 MUX2_X1 _59744_ (.A(\icache.tag_tv_r [26]),
    .B(\icache.tag_mem.data_o [26]),
    .S(_26557_),
    .Z(_04701_));
 MUX2_X1 _59745_ (.A(\icache.tag_tv_r [27]),
    .B(\icache.tag_mem.data_o [29]),
    .S(_26557_),
    .Z(_04702_));
 MUX2_X1 _59746_ (.A(\icache.tag_tv_r [28]),
    .B(\icache.tag_mem.data_o [30]),
    .S(_26557_),
    .Z(_04703_));
 BUF_X4 _59747_ (.A(_26554_),
    .Z(_26558_));
 MUX2_X1 _59748_ (.A(\icache.tag_tv_r [29]),
    .B(\icache.tag_mem.data_o [31]),
    .S(_26558_),
    .Z(_04704_));
 MUX2_X1 _59749_ (.A(\icache.tag_tv_r [30]),
    .B(\icache.tag_mem.data_o [32]),
    .S(_26558_),
    .Z(_04706_));
 MUX2_X1 _59750_ (.A(\icache.tag_tv_r [31]),
    .B(\icache.tag_mem.data_o [33]),
    .S(_26558_),
    .Z(_04707_));
 MUX2_X1 _59751_ (.A(\icache.tag_tv_r [32]),
    .B(\icache.tag_mem.data_o [34]),
    .S(_26558_),
    .Z(_04708_));
 MUX2_X1 _59752_ (.A(\icache.tag_tv_r [33]),
    .B(\icache.tag_mem.data_o [35]),
    .S(_26558_),
    .Z(_04709_));
 MUX2_X1 _59753_ (.A(\icache.tag_tv_r [34]),
    .B(\icache.tag_mem.data_o [36]),
    .S(_26558_),
    .Z(_04710_));
 MUX2_X1 _59754_ (.A(\icache.tag_tv_r [35]),
    .B(\icache.tag_mem.data_o [37]),
    .S(_26558_),
    .Z(_04711_));
 MUX2_X1 _59755_ (.A(\icache.tag_tv_r [36]),
    .B(\icache.tag_mem.data_o [38]),
    .S(_26558_),
    .Z(_04712_));
 MUX2_X1 _59756_ (.A(\icache.tag_tv_r [37]),
    .B(\icache.tag_mem.data_o [39]),
    .S(_26558_),
    .Z(_04713_));
 MUX2_X1 _59757_ (.A(\icache.tag_tv_r [38]),
    .B(\icache.tag_mem.data_o [40]),
    .S(_26558_),
    .Z(_04714_));
 BUF_X4 _59758_ (.A(_26554_),
    .Z(_26559_));
 MUX2_X1 _59759_ (.A(\icache.tag_tv_r [39]),
    .B(\icache.tag_mem.data_o [41]),
    .S(_26559_),
    .Z(_04715_));
 MUX2_X1 _59760_ (.A(\icache.tag_tv_r [40]),
    .B(\icache.tag_mem.data_o [42]),
    .S(_26559_),
    .Z(_04717_));
 MUX2_X1 _59761_ (.A(\icache.tag_tv_r [41]),
    .B(\icache.tag_mem.data_o [43]),
    .S(_26559_),
    .Z(_04718_));
 MUX2_X1 _59762_ (.A(\icache.tag_tv_r [42]),
    .B(\icache.tag_mem.data_o [44]),
    .S(_26559_),
    .Z(_04719_));
 MUX2_X1 _59763_ (.A(\icache.tag_tv_r [43]),
    .B(\icache.tag_mem.data_o [45]),
    .S(_26559_),
    .Z(_04720_));
 MUX2_X1 _59764_ (.A(\icache.tag_tv_r [44]),
    .B(\icache.tag_mem.data_o [46]),
    .S(_26559_),
    .Z(_04721_));
 MUX2_X1 _59765_ (.A(\icache.tag_tv_r [45]),
    .B(\icache.tag_mem.data_o [47]),
    .S(_26559_),
    .Z(_04722_));
 MUX2_X1 _59766_ (.A(\icache.tag_tv_r [46]),
    .B(\icache.tag_mem.data_o [48]),
    .S(_26559_),
    .Z(_04723_));
 MUX2_X1 _59767_ (.A(\icache.tag_tv_r [47]),
    .B(\icache.tag_mem.data_o [49]),
    .S(_26559_),
    .Z(_04724_));
 MUX2_X1 _59768_ (.A(\icache.tag_tv_r [48]),
    .B(\icache.tag_mem.data_o [50]),
    .S(_26559_),
    .Z(_04725_));
 BUF_X4 _59769_ (.A(_26554_),
    .Z(_26560_));
 MUX2_X1 _59770_ (.A(\icache.tag_tv_r [49]),
    .B(\icache.tag_mem.data_o [51]),
    .S(_26560_),
    .Z(_04726_));
 MUX2_X1 _59771_ (.A(\icache.tag_tv_r [50]),
    .B(\icache.tag_mem.data_o [52]),
    .S(_26560_),
    .Z(_04728_));
 MUX2_X1 _59772_ (.A(\icache.tag_tv_r [51]),
    .B(\icache.tag_mem.data_o [53]),
    .S(_26560_),
    .Z(_04729_));
 MUX2_X1 _59773_ (.A(\icache.tag_tv_r [52]),
    .B(\icache.tag_mem.data_o [54]),
    .S(_26560_),
    .Z(_04730_));
 MUX2_X1 _59774_ (.A(\icache.tag_tv_r [53]),
    .B(\icache.tag_mem.data_o [55]),
    .S(_26560_),
    .Z(_04731_));
 MUX2_X1 _59775_ (.A(\icache.tag_tv_r [54]),
    .B(\icache.tag_mem.data_o [58]),
    .S(_26560_),
    .Z(_04732_));
 MUX2_X1 _59776_ (.A(\icache.tag_tv_r [55]),
    .B(\icache.tag_mem.data_o [59]),
    .S(_26560_),
    .Z(_04733_));
 MUX2_X1 _59777_ (.A(\icache.tag_tv_r [56]),
    .B(\icache.tag_mem.data_o [60]),
    .S(_26560_),
    .Z(_04734_));
 MUX2_X1 _59778_ (.A(\icache.tag_tv_r [57]),
    .B(\icache.tag_mem.data_o [61]),
    .S(_26560_),
    .Z(_04735_));
 MUX2_X1 _59779_ (.A(\icache.tag_tv_r [58]),
    .B(\icache.tag_mem.data_o [62]),
    .S(_26560_),
    .Z(_04736_));
 BUF_X4 _59780_ (.A(_26554_),
    .Z(_26561_));
 MUX2_X1 _59781_ (.A(\icache.tag_tv_r [59]),
    .B(\icache.tag_mem.data_o [63]),
    .S(_26561_),
    .Z(_04737_));
 MUX2_X1 _59782_ (.A(\icache.tag_tv_r [60]),
    .B(\icache.tag_mem.data_o [64]),
    .S(_26561_),
    .Z(_04739_));
 MUX2_X1 _59783_ (.A(\icache.tag_tv_r [61]),
    .B(\icache.tag_mem.data_o [65]),
    .S(_26561_),
    .Z(_04740_));
 MUX2_X1 _59784_ (.A(\icache.tag_tv_r [62]),
    .B(\icache.tag_mem.data_o [66]),
    .S(_26561_),
    .Z(_04741_));
 MUX2_X1 _59785_ (.A(\icache.tag_tv_r [63]),
    .B(\icache.tag_mem.data_o [67]),
    .S(_26561_),
    .Z(_04742_));
 MUX2_X1 _59786_ (.A(\icache.tag_tv_r [64]),
    .B(\icache.tag_mem.data_o [68]),
    .S(_26561_),
    .Z(_04743_));
 MUX2_X1 _59787_ (.A(\icache.tag_tv_r [65]),
    .B(\icache.tag_mem.data_o [69]),
    .S(_26561_),
    .Z(_04744_));
 MUX2_X1 _59788_ (.A(\icache.tag_tv_r [66]),
    .B(\icache.tag_mem.data_o [70]),
    .S(_26561_),
    .Z(_04745_));
 MUX2_X1 _59789_ (.A(\icache.tag_tv_r [67]),
    .B(\icache.tag_mem.data_o [71]),
    .S(_26561_),
    .Z(_04746_));
 MUX2_X1 _59790_ (.A(\icache.tag_tv_r [68]),
    .B(\icache.tag_mem.data_o [72]),
    .S(_26561_),
    .Z(_04747_));
 BUF_X4 _59791_ (.A(_26554_),
    .Z(_26562_));
 MUX2_X1 _59792_ (.A(\icache.tag_tv_r [69]),
    .B(\icache.tag_mem.data_o [73]),
    .S(_26562_),
    .Z(_04748_));
 MUX2_X1 _59793_ (.A(\icache.tag_tv_r [70]),
    .B(\icache.tag_mem.data_o [74]),
    .S(_26562_),
    .Z(_04750_));
 MUX2_X1 _59794_ (.A(\icache.tag_tv_r [71]),
    .B(\icache.tag_mem.data_o [75]),
    .S(_26562_),
    .Z(_04751_));
 MUX2_X1 _59795_ (.A(\icache.tag_tv_r [72]),
    .B(\icache.tag_mem.data_o [76]),
    .S(_26562_),
    .Z(_04752_));
 MUX2_X1 _59796_ (.A(\icache.tag_tv_r [73]),
    .B(\icache.tag_mem.data_o [77]),
    .S(_26562_),
    .Z(_04753_));
 MUX2_X1 _59797_ (.A(\icache.tag_tv_r [74]),
    .B(\icache.tag_mem.data_o [78]),
    .S(_26562_),
    .Z(_04754_));
 MUX2_X1 _59798_ (.A(\icache.tag_tv_r [75]),
    .B(\icache.tag_mem.data_o [79]),
    .S(_26562_),
    .Z(_04755_));
 MUX2_X1 _59799_ (.A(\icache.tag_tv_r [76]),
    .B(\icache.tag_mem.data_o [80]),
    .S(_26562_),
    .Z(_04756_));
 MUX2_X1 _59800_ (.A(\icache.tag_tv_r [77]),
    .B(\icache.tag_mem.data_o [81]),
    .S(_26562_),
    .Z(_04757_));
 MUX2_X1 _59801_ (.A(\icache.tag_tv_r [78]),
    .B(\icache.tag_mem.data_o [82]),
    .S(_26562_),
    .Z(_04758_));
 BUF_X4 _59802_ (.A(_26554_),
    .Z(_26563_));
 MUX2_X1 _59803_ (.A(\icache.tag_tv_r [79]),
    .B(\icache.tag_mem.data_o [83]),
    .S(_26563_),
    .Z(_04759_));
 MUX2_X1 _59804_ (.A(\icache.tag_tv_r [80]),
    .B(\icache.tag_mem.data_o [84]),
    .S(_26563_),
    .Z(_04761_));
 MUX2_X1 _59805_ (.A(\icache.tag_tv_r [81]),
    .B(\icache.tag_mem.data_o [87]),
    .S(_26563_),
    .Z(_04762_));
 MUX2_X1 _59806_ (.A(\icache.tag_tv_r [82]),
    .B(\icache.tag_mem.data_o [88]),
    .S(_26563_),
    .Z(_04763_));
 MUX2_X1 _59807_ (.A(\icache.tag_tv_r [83]),
    .B(\icache.tag_mem.data_o [89]),
    .S(_26563_),
    .Z(_04764_));
 MUX2_X1 _59808_ (.A(\icache.tag_tv_r [84]),
    .B(\icache.tag_mem.data_o [90]),
    .S(_26563_),
    .Z(_04765_));
 MUX2_X1 _59809_ (.A(\icache.tag_tv_r [85]),
    .B(\icache.tag_mem.data_o [91]),
    .S(_26563_),
    .Z(_04766_));
 MUX2_X1 _59810_ (.A(\icache.tag_tv_r [86]),
    .B(\icache.tag_mem.data_o [92]),
    .S(_26563_),
    .Z(_04767_));
 MUX2_X1 _59811_ (.A(\icache.tag_tv_r [87]),
    .B(\icache.tag_mem.data_o [93]),
    .S(_26563_),
    .Z(_04768_));
 MUX2_X1 _59812_ (.A(\icache.tag_tv_r [88]),
    .B(\icache.tag_mem.data_o [94]),
    .S(_26563_),
    .Z(_04769_));
 BUF_X4 _59813_ (.A(_26554_),
    .Z(_26564_));
 MUX2_X1 _59814_ (.A(\icache.tag_tv_r [89]),
    .B(\icache.tag_mem.data_o [95]),
    .S(_26564_),
    .Z(_04770_));
 MUX2_X1 _59815_ (.A(\icache.tag_tv_r [90]),
    .B(\icache.tag_mem.data_o [96]),
    .S(_26564_),
    .Z(_04772_));
 MUX2_X1 _59816_ (.A(\icache.tag_tv_r [91]),
    .B(\icache.tag_mem.data_o [97]),
    .S(_26564_),
    .Z(_04773_));
 MUX2_X1 _59817_ (.A(\icache.tag_tv_r [92]),
    .B(\icache.tag_mem.data_o [98]),
    .S(_26564_),
    .Z(_04774_));
 MUX2_X1 _59818_ (.A(\icache.tag_tv_r [93]),
    .B(\icache.tag_mem.data_o [99]),
    .S(_26564_),
    .Z(_04775_));
 MUX2_X1 _59819_ (.A(\icache.tag_tv_r [94]),
    .B(\icache.tag_mem.data_o [100]),
    .S(_26564_),
    .Z(_04776_));
 MUX2_X1 _59820_ (.A(\icache.tag_tv_r [95]),
    .B(\icache.tag_mem.data_o [101]),
    .S(_26564_),
    .Z(_04777_));
 MUX2_X1 _59821_ (.A(\icache.tag_tv_r [96]),
    .B(\icache.tag_mem.data_o [102]),
    .S(_26564_),
    .Z(_04778_));
 MUX2_X1 _59822_ (.A(\icache.tag_tv_r [97]),
    .B(\icache.tag_mem.data_o [103]),
    .S(_26564_),
    .Z(_04779_));
 MUX2_X1 _59823_ (.A(\icache.tag_tv_r [98]),
    .B(\icache.tag_mem.data_o [104]),
    .S(_26564_),
    .Z(_04780_));
 BUF_X16 _59824_ (.A(_26473_),
    .Z(_26565_));
 MUX2_X1 _59825_ (.A(\icache.tag_tv_r [99]),
    .B(\icache.tag_mem.data_o [105]),
    .S(_26565_),
    .Z(_04781_));
 MUX2_X1 _59826_ (.A(\icache.tag_tv_r [100]),
    .B(\icache.tag_mem.data_o [106]),
    .S(_26565_),
    .Z(_04568_));
 MUX2_X1 _59827_ (.A(\icache.tag_tv_r [101]),
    .B(\icache.tag_mem.data_o [107]),
    .S(_26565_),
    .Z(_04569_));
 MUX2_X1 _59828_ (.A(\icache.tag_tv_r [102]),
    .B(\icache.tag_mem.data_o [108]),
    .S(_26565_),
    .Z(_04570_));
 MUX2_X1 _59829_ (.A(\icache.tag_tv_r [103]),
    .B(\icache.tag_mem.data_o [109]),
    .S(_26565_),
    .Z(_04571_));
 MUX2_X1 _59830_ (.A(\icache.tag_tv_r [104]),
    .B(\icache.tag_mem.data_o [110]),
    .S(_26565_),
    .Z(_04572_));
 MUX2_X1 _59831_ (.A(\icache.tag_tv_r [105]),
    .B(\icache.tag_mem.data_o [111]),
    .S(_26565_),
    .Z(_04573_));
 MUX2_X1 _59832_ (.A(\icache.tag_tv_r [106]),
    .B(\icache.tag_mem.data_o [112]),
    .S(_26565_),
    .Z(_04574_));
 MUX2_X1 _59833_ (.A(\icache.tag_tv_r [107]),
    .B(\icache.tag_mem.data_o [113]),
    .S(_26565_),
    .Z(_04575_));
 MUX2_X1 _59834_ (.A(\icache.tag_tv_r [108]),
    .B(\icache.tag_mem.data_o [116]),
    .S(_26565_),
    .Z(_04576_));
 BUF_X8 _59835_ (.A(_26473_),
    .Z(_26566_));
 MUX2_X1 _59836_ (.A(net1302),
    .B(\icache.tag_mem.data_o [117]),
    .S(_26566_),
    .Z(_04577_));
 MUX2_X1 _59837_ (.A(net1301),
    .B(\icache.tag_mem.data_o [118]),
    .S(_26566_),
    .Z(_04579_));
 MUX2_X1 _59838_ (.A(net1300),
    .B(\icache.tag_mem.data_o [119]),
    .S(_26566_),
    .Z(_04580_));
 MUX2_X1 _59839_ (.A(net1299),
    .B(\icache.tag_mem.data_o [120]),
    .S(_26566_),
    .Z(_04581_));
 MUX2_X1 _59840_ (.A(net1297),
    .B(\icache.tag_mem.data_o [121]),
    .S(_26566_),
    .Z(_04582_));
 MUX2_X1 _59841_ (.A(net1296),
    .B(\icache.tag_mem.data_o [122]),
    .S(_26566_),
    .Z(_04583_));
 MUX2_X1 _59842_ (.A(net1293),
    .B(\icache.tag_mem.data_o [123]),
    .S(_26566_),
    .Z(_04584_));
 MUX2_X1 _59843_ (.A(net1292),
    .B(\icache.tag_mem.data_o [124]),
    .S(_26566_),
    .Z(_04585_));
 MUX2_X1 _59844_ (.A(net1291),
    .B(\icache.tag_mem.data_o [125]),
    .S(_26566_),
    .Z(_04586_));
 MUX2_X1 _59845_ (.A(net1290),
    .B(\icache.tag_mem.data_o [126]),
    .S(_26566_),
    .Z(_04587_));
 BUF_X4 _59846_ (.A(_26473_),
    .Z(_26567_));
 MUX2_X1 _59847_ (.A(net1289),
    .B(\icache.tag_mem.data_o [127]),
    .S(_26567_),
    .Z(_04588_));
 MUX2_X1 _59848_ (.A(net1288),
    .B(\icache.tag_mem.data_o [128]),
    .S(_26567_),
    .Z(_04590_));
 MUX2_X1 _59849_ (.A(net1286),
    .B(\icache.tag_mem.data_o [129]),
    .S(_26567_),
    .Z(_04591_));
 MUX2_X1 _59850_ (.A(net1284),
    .B(\icache.tag_mem.data_o [130]),
    .S(_26567_),
    .Z(_04592_));
 MUX2_X1 _59851_ (.A(net1283),
    .B(\icache.tag_mem.data_o [131]),
    .S(_26567_),
    .Z(_04593_));
 MUX2_X1 _59852_ (.A(net1280),
    .B(\icache.tag_mem.data_o [132]),
    .S(_26567_),
    .Z(_04594_));
 MUX2_X1 _59853_ (.A(net1279),
    .B(\icache.tag_mem.data_o [133]),
    .S(_26567_),
    .Z(_04595_));
 MUX2_X1 _59854_ (.A(net1278),
    .B(\icache.tag_mem.data_o [134]),
    .S(_26567_),
    .Z(_04596_));
 MUX2_X1 _59855_ (.A(net1277),
    .B(\icache.tag_mem.data_o [135]),
    .S(_26567_),
    .Z(_04597_));
 MUX2_X1 _59856_ (.A(net1276),
    .B(\icache.tag_mem.data_o [136]),
    .S(_26567_),
    .Z(_04598_));
 BUF_X4 _59857_ (.A(_26473_),
    .Z(_26568_));
 MUX2_X1 _59858_ (.A(net1275),
    .B(\icache.tag_mem.data_o [137]),
    .S(_26568_),
    .Z(_04599_));
 MUX2_X1 _59859_ (.A(net1274),
    .B(\icache.tag_mem.data_o [138]),
    .S(_26568_),
    .Z(_04601_));
 MUX2_X1 _59860_ (.A(\icache.tag_tv_r [131]),
    .B(\icache.tag_mem.data_o [139]),
    .S(_26568_),
    .Z(_04602_));
 MUX2_X1 _59861_ (.A(net1273),
    .B(\icache.tag_mem.data_o [140]),
    .S(_26568_),
    .Z(_04603_));
 MUX2_X1 _59862_ (.A(net1272),
    .B(\icache.tag_mem.data_o [141]),
    .S(_26568_),
    .Z(_04604_));
 MUX2_X1 _59863_ (.A(net1271),
    .B(\icache.tag_mem.data_o [142]),
    .S(_26568_),
    .Z(_04605_));
 MUX2_X1 _59864_ (.A(net1270),
    .B(\icache.tag_mem.data_o [145]),
    .S(_26568_),
    .Z(_04606_));
 MUX2_X1 _59865_ (.A(net1269),
    .B(\icache.tag_mem.data_o [146]),
    .S(_26568_),
    .Z(_04607_));
 MUX2_X1 _59866_ (.A(net1268),
    .B(\icache.tag_mem.data_o [147]),
    .S(_26568_),
    .Z(_04608_));
 MUX2_X1 _59867_ (.A(net1267),
    .B(\icache.tag_mem.data_o [148]),
    .S(_26568_),
    .Z(_04609_));
 BUF_X4 _59868_ (.A(_26473_),
    .Z(_26569_));
 MUX2_X1 _59869_ (.A(\icache.tag_tv_r [139]),
    .B(\icache.tag_mem.data_o [149]),
    .S(_26569_),
    .Z(_04610_));
 MUX2_X1 _59870_ (.A(\icache.tag_tv_r [140]),
    .B(\icache.tag_mem.data_o [150]),
    .S(_26569_),
    .Z(_04612_));
 MUX2_X1 _59871_ (.A(\icache.tag_tv_r [141]),
    .B(\icache.tag_mem.data_o [151]),
    .S(_26569_),
    .Z(_04613_));
 MUX2_X1 _59872_ (.A(\icache.tag_tv_r [142]),
    .B(\icache.tag_mem.data_o [152]),
    .S(_26569_),
    .Z(_04614_));
 MUX2_X1 _59873_ (.A(\icache.tag_tv_r [143]),
    .B(\icache.tag_mem.data_o [153]),
    .S(_26569_),
    .Z(_04615_));
 MUX2_X1 _59874_ (.A(\icache.tag_tv_r [144]),
    .B(\icache.tag_mem.data_o [154]),
    .S(_26569_),
    .Z(_04616_));
 MUX2_X1 _59875_ (.A(\icache.tag_tv_r [145]),
    .B(\icache.tag_mem.data_o [155]),
    .S(_26569_),
    .Z(_04617_));
 MUX2_X1 _59876_ (.A(\icache.tag_tv_r [146]),
    .B(\icache.tag_mem.data_o [156]),
    .S(_26569_),
    .Z(_04618_));
 MUX2_X1 _59877_ (.A(\icache.tag_tv_r [147]),
    .B(\icache.tag_mem.data_o [157]),
    .S(_26569_),
    .Z(_04619_));
 MUX2_X1 _59878_ (.A(\icache.tag_tv_r [148]),
    .B(\icache.tag_mem.data_o [158]),
    .S(_26569_),
    .Z(_04620_));
 MUX2_X1 _59879_ (.A(\icache.tag_tv_r [149]),
    .B(\icache.tag_mem.data_o [159]),
    .S(_08518_),
    .Z(_04621_));
 MUX2_X1 _59880_ (.A(\icache.tag_tv_r [150]),
    .B(\icache.tag_mem.data_o [160]),
    .S(_08518_),
    .Z(_04623_));
 OAI211_X2 _59881_ (.A(_26503_),
    .B(_08727_),
    .C1(_08499_),
    .C2(_15275_),
    .ZN(_26570_));
 OAI21_X4 _59882_ (.A(_26570_),
    .B1(_08481_),
    .B2(_09000_),
    .ZN(\icache.data_mems_0__data_mem.v_i ));
 AOI21_X4 _59883_ (.A(_08651_),
    .B1(_08481_),
    .B2(_10729_),
    .ZN(\icache.n_0_net_ ));
 OAI211_X4 _59884_ (.A(_10657_),
    .B(_10730_),
    .C1(_10731_),
    .C2(_10717_),
    .ZN(lce_resp_v_o));
 OR2_X1 _59885_ (.A1(_21275_),
    .A2(\icache.lce.lce_cmd_inst.rv_adapter.full_r ),
    .ZN(_26571_));
 AOI21_X1 _59886_ (.A(_21259_),
    .B1(_26571_),
    .B2(_00001_),
    .ZN(_26572_));
 OR2_X1 _59887_ (.A1(_26572_),
    .A2(_21279_),
    .ZN(\icache.lce.lce_cmd_inst.rv_adapter.N13 ));
 AOI21_X1 _59888_ (.A(_15281_),
    .B1(_20982_),
    .B2(_21281_),
    .ZN(_26573_));
 OAI21_X1 _59889_ (.A(_08675_),
    .B1(_26573_),
    .B2(_21282_),
    .ZN(\icache.lce.lce_data_cmd.rv_adapter.N13 ));
 NOR4_X4 _59890_ (.A1(_08038_),
    .A2(_08499_),
    .A3(_15279_),
    .A4(_15274_),
    .ZN(\icache.data_mem_w_li ));
 AOI21_X4 _59891_ (.A(_08651_),
    .B1(_10722_),
    .B2(_21266_),
    .ZN(\icache.n_9_net_ ));
 DFF_X1 _59892_ (.D(_00610_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.N79 ),
    .QN(_26574_));
 DFF_X1 _59893_ (.D(_00621_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.N80 ),
    .QN(_26575_));
 DFF_X1 _59894_ (.D(_00632_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if1_r [2]),
    .QN(_26576_));
 DFF_X1 _59895_ (.D(_00642_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if1_r [3]),
    .QN(_26577_));
 DFF_X1 _59896_ (.D(_00643_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if1_r [4]),
    .QN(_26578_));
 DFF_X1 _59897_ (.D(_00644_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if1_r [5]),
    .QN(_26579_));
 DFF_X1 _59898_ (.D(_00645_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if1_r [6]),
    .QN(_00005_));
 DFF_X1 _59899_ (.D(_00646_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if1_r [7]),
    .QN(_26580_));
 DFF_X1 _59900_ (.D(_00647_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if1_r [8]),
    .QN(_00073_));
 DFF_X1 _59901_ (.D(_00648_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if1_r [9]),
    .QN(_26581_));
 DFF_X1 _59902_ (.D(_00611_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if1_r [10]),
    .QN(_00074_));
 DFF_X1 _59903_ (.D(_00612_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if1_r [11]),
    .QN(_26582_));
 DFF_X1 _59904_ (.D(_00613_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if1_r [12]),
    .QN(_00083_));
 DFF_X1 _59905_ (.D(_00614_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if1_r [13]),
    .QN(_26583_));
 DFF_X1 _59906_ (.D(_00615_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if1_r [14]),
    .QN(_00084_));
 DFF_X1 _59907_ (.D(_00616_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if1_r [15]),
    .QN(_26584_));
 DFF_X1 _59908_ (.D(_00617_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if1_r [16]),
    .QN(_00085_));
 DFF_X1 _59909_ (.D(_00618_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if1_r [17]),
    .QN(_26585_));
 DFF_X1 _59910_ (.D(_00619_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if1_r [18]),
    .QN(_00086_));
 DFF_X1 _59911_ (.D(_00620_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if1_r [19]),
    .QN(_26586_));
 DFF_X1 _59912_ (.D(_00622_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if1_r [20]),
    .QN(_00087_));
 DFF_X1 _59913_ (.D(_00623_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if1_r [21]),
    .QN(_26587_));
 DFF_X1 _59914_ (.D(_00624_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if1_r [22]),
    .QN(_00088_));
 DFF_X1 _59915_ (.D(_00625_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if1_r [23]),
    .QN(_26588_));
 DFF_X1 _59916_ (.D(_00626_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if1_r [24]),
    .QN(_00089_));
 DFF_X1 _59917_ (.D(_00627_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if1_r [25]),
    .QN(_26589_));
 DFF_X1 _59918_ (.D(_00628_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if1_r [26]),
    .QN(_00090_));
 DFF_X1 _59919_ (.D(_00629_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if1_r [27]),
    .QN(_26590_));
 DFF_X1 _59920_ (.D(_00630_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if1_r [28]),
    .QN(_00091_));
 DFF_X1 _59921_ (.D(_00631_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if1_r [29]),
    .QN(_26591_));
 DFF_X1 _59922_ (.D(_00633_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if1_r [30]),
    .QN(_00092_));
 DFF_X1 _59923_ (.D(_00634_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if1_r [31]),
    .QN(_26592_));
 DFF_X1 _59924_ (.D(_00635_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if1_r [32]),
    .QN(_00093_));
 DFF_X1 _59925_ (.D(_00636_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if1_r [33]),
    .QN(_26593_));
 DFF_X1 _59926_ (.D(_00637_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if1_r [34]),
    .QN(_00094_));
 DFF_X1 _59927_ (.D(_00638_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if1_r [35]),
    .QN(_26594_));
 DFF_X1 _59928_ (.D(_00639_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if1_r [36]),
    .QN(_00095_));
 DFF_X1 _59929_ (.D(_00640_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if1_r [37]),
    .QN(_26595_));
 DFF_X1 _59930_ (.D(_00641_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if1_r [38]),
    .QN(_26596_));
 DFF_X1 _59931_ (.D(_00728_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_v_if2_r ),
    .QN(_00080_));
 DFF_X1 _59932_ (.D(_00727_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_v_if1_r ),
    .QN(_26597_));
 DFF_X1 _59933_ (.D(_00609_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.itlb_miss_if2_r ),
    .QN(_26598_));
 DFF_X1 _59934_ (.D(_00729_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.state_r [0]),
    .QN(_26599_));
 DFF_X1 _59935_ (.D(_00730_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.state_r [1]),
    .QN(_26600_));
 DFF_X1 _59936_ (.D(_00649_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if2_r [0]),
    .QN(_00078_));
 DFF_X1 _59937_ (.D(_00660_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if2_r [1]),
    .QN(_00079_));
 DFF_X1 _59938_ (.D(_00671_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if2_r [2]),
    .QN(_26601_));
 DFF_X1 _59939_ (.D(_00681_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if2_r [3]),
    .QN(_26602_));
 DFF_X1 _59940_ (.D(_00682_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if2_r [4]),
    .QN(_26603_));
 DFF_X1 _59941_ (.D(_00683_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if2_r [5]),
    .QN(_26604_));
 DFF_X1 _59942_ (.D(_00684_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if2_r [6]),
    .QN(_26605_));
 DFF_X1 _59943_ (.D(_00685_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if2_r [7]),
    .QN(_26606_));
 DFF_X1 _59944_ (.D(_00686_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if2_r [8]),
    .QN(_26607_));
 DFF_X1 _59945_ (.D(_00687_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if2_r [9]),
    .QN(_26608_));
 DFF_X1 _59946_ (.D(_00650_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if2_r [10]),
    .QN(_26609_));
 DFF_X1 _59947_ (.D(_00651_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if2_r [11]),
    .QN(_26610_));
 DFF_X1 _59948_ (.D(_00652_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if2_r [12]),
    .QN(_26611_));
 DFF_X1 _59949_ (.D(_00653_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if2_r [13]),
    .QN(_26612_));
 DFF_X1 _59950_ (.D(_00654_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if2_r [14]),
    .QN(_26613_));
 DFF_X1 _59951_ (.D(_00655_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if2_r [15]),
    .QN(_26614_));
 DFF_X1 _59952_ (.D(_00656_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if2_r [16]),
    .QN(_26615_));
 DFF_X1 _59953_ (.D(_00657_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if2_r [17]),
    .QN(_26616_));
 DFF_X1 _59954_ (.D(_00658_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if2_r [18]),
    .QN(_26617_));
 DFF_X1 _59955_ (.D(_00659_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if2_r [19]),
    .QN(_26618_));
 DFF_X1 _59956_ (.D(_00661_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if2_r [20]),
    .QN(_26619_));
 DFF_X1 _59957_ (.D(_00662_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if2_r [21]),
    .QN(_26620_));
 DFF_X1 _59958_ (.D(_00663_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if2_r [22]),
    .QN(_26621_));
 DFF_X1 _59959_ (.D(_00664_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if2_r [23]),
    .QN(_26622_));
 DFF_X1 _59960_ (.D(_00665_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if2_r [24]),
    .QN(_26623_));
 DFF_X1 _59961_ (.D(_00666_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if2_r [25]),
    .QN(_26624_));
 DFF_X1 _59962_ (.D(_00667_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if2_r [26]),
    .QN(_26625_));
 DFF_X1 _59963_ (.D(_00668_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if2_r [27]),
    .QN(_26626_));
 DFF_X1 _59964_ (.D(_00669_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if2_r [28]),
    .QN(_26627_));
 DFF_X1 _59965_ (.D(_00670_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if2_r [29]),
    .QN(_26628_));
 DFF_X1 _59966_ (.D(_00672_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if2_r [30]),
    .QN(_26629_));
 DFF_X1 _59967_ (.D(_00673_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if2_r [31]),
    .QN(_26630_));
 DFF_X1 _59968_ (.D(_00674_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if2_r [32]),
    .QN(_26631_));
 DFF_X1 _59969_ (.D(_00675_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if2_r [33]),
    .QN(_26632_));
 DFF_X1 _59970_ (.D(_00676_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if2_r [34]),
    .QN(_26633_));
 DFF_X1 _59971_ (.D(_00677_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if2_r [35]),
    .QN(_26634_));
 DFF_X1 _59972_ (.D(_00678_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if2_r [36]),
    .QN(_26635_));
 DFF_X1 _59973_ (.D(_00679_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if2_r [37]),
    .QN(_26636_));
 DFF_X1 _59974_ (.D(_00680_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_if2_r [38]),
    .QN(_26637_));
 DFF_X1 _59975_ (.D(_00688_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_resume_r [0]),
    .QN(_26638_));
 DFF_X1 _59976_ (.D(_00699_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_resume_r [1]),
    .QN(_26639_));
 DFF_X1 _59977_ (.D(_00710_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_resume_r [2]),
    .QN(_00081_));
 DFF_X1 _59978_ (.D(_00720_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_resume_r [3]),
    .QN(_00076_));
 DFF_X1 _59979_ (.D(_00721_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_resume_r [4]),
    .QN(_26640_));
 DFF_X1 _59980_ (.D(_00722_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_resume_r [5]),
    .QN(_26641_));
 DFF_X1 _59981_ (.D(_00723_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_resume_r [6]),
    .QN(_26642_));
 DFF_X1 _59982_ (.D(_00724_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_resume_r [7]),
    .QN(_26643_));
 DFF_X1 _59983_ (.D(_00725_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_resume_r [8]),
    .QN(_26644_));
 DFF_X1 _59984_ (.D(_00726_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_resume_r [9]),
    .QN(_26645_));
 DFF_X1 _59985_ (.D(_00689_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_resume_r [10]),
    .QN(_26646_));
 DFF_X1 _59986_ (.D(_00690_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_resume_r [11]),
    .QN(_26647_));
 DFF_X1 _59987_ (.D(_00691_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_resume_r [12]),
    .QN(_26648_));
 DFF_X1 _59988_ (.D(_00692_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_resume_r [13]),
    .QN(_26649_));
 DFF_X1 _59989_ (.D(_00693_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_resume_r [14]),
    .QN(_26650_));
 DFF_X1 _59990_ (.D(_00694_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_resume_r [15]),
    .QN(_26651_));
 DFF_X1 _59991_ (.D(_00695_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_resume_r [16]),
    .QN(_26652_));
 DFF_X1 _59992_ (.D(_00696_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_resume_r [17]),
    .QN(_26653_));
 DFF_X1 _59993_ (.D(_00697_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_resume_r [18]),
    .QN(_26654_));
 DFF_X1 _59994_ (.D(_00698_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_resume_r [19]),
    .QN(_26655_));
 DFF_X1 _59995_ (.D(_00700_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_resume_r [20]),
    .QN(_26656_));
 DFF_X1 _59996_ (.D(_00701_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_resume_r [21]),
    .QN(_26657_));
 DFF_X1 _59997_ (.D(_00702_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_resume_r [22]),
    .QN(_26658_));
 DFF_X1 _59998_ (.D(_00703_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_resume_r [23]),
    .QN(_26659_));
 DFF_X1 _59999_ (.D(_00704_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_resume_r [24]),
    .QN(_26660_));
 DFF_X1 _60000_ (.D(_00705_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_resume_r [25]),
    .QN(_26661_));
 DFF_X1 _60001_ (.D(_00706_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_resume_r [26]),
    .QN(_26662_));
 DFF_X1 _60002_ (.D(_00707_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_resume_r [27]),
    .QN(_26663_));
 DFF_X1 _60003_ (.D(_00708_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_resume_r [28]),
    .QN(_26664_));
 DFF_X1 _60004_ (.D(_00709_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_resume_r [29]),
    .QN(_26665_));
 DFF_X1 _60005_ (.D(_00711_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_resume_r [30]),
    .QN(_26666_));
 DFF_X1 _60006_ (.D(_00712_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_resume_r [31]),
    .QN(_26667_));
 DFF_X1 _60007_ (.D(_00713_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_resume_r [32]),
    .QN(_26668_));
 DFF_X1 _60008_ (.D(_00714_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_resume_r [33]),
    .QN(_26669_));
 DFF_X1 _60009_ (.D(_00715_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_resume_r [34]),
    .QN(_26670_));
 DFF_X1 _60010_ (.D(_00716_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_resume_r [35]),
    .QN(_26671_));
 DFF_X1 _60011_ (.D(_00717_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_resume_r [36]),
    .QN(_26672_));
 DFF_X1 _60012_ (.D(_00718_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_resume_r [37]),
    .QN(_26673_));
 DFF_X1 _60013_ (.D(_00719_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.pc_resume_r [38]),
    .QN(_26674_));
 DFF_X1 _60014_ (.D(\itlb.entry_ram.z_s1r1w_data_lo [0]),
    .CK(clk_i),
    .Q(\icache.uncached_i ),
    .QN(_26675_));
 DFF_X1 _60015_ (.D(\itlb.entry_ram.z_s1r1w_data_lo [6]),
    .CK(clk_i),
    .Q(\icache.itlb_icache_data_resp_i [0]),
    .QN(_26676_));
 DFF_X1 _60016_ (.D(\itlb.entry_ram.z_s1r1w_data_lo [7]),
    .CK(clk_i),
    .Q(\icache.itlb_icache_data_resp_i [1]),
    .QN(_26677_));
 DFF_X1 _60017_ (.D(\itlb.entry_ram.z_s1r1w_data_lo [8]),
    .CK(clk_i),
    .Q(\icache.itlb_icache_data_resp_i [2]),
    .QN(_26678_));
 DFF_X1 _60018_ (.D(\itlb.entry_ram.z_s1r1w_data_lo [9]),
    .CK(clk_i),
    .Q(\icache.itlb_icache_data_resp_i [3]),
    .QN(_26679_));
 DFF_X1 _60019_ (.D(\itlb.entry_ram.z_s1r1w_data_lo [10]),
    .CK(clk_i),
    .Q(\icache.itlb_icache_data_resp_i [4]),
    .QN(_26680_));
 DFF_X1 _60020_ (.D(\itlb.entry_ram.z_s1r1w_data_lo [11]),
    .CK(clk_i),
    .Q(\icache.itlb_icache_data_resp_i [5]),
    .QN(_26681_));
 DFF_X1 _60021_ (.D(\itlb.entry_ram.z_s1r1w_data_lo [12]),
    .CK(clk_i),
    .Q(\icache.itlb_icache_data_resp_i [6]),
    .QN(_26682_));
 DFF_X1 _60022_ (.D(\itlb.entry_ram.z_s1r1w_data_lo [13]),
    .CK(clk_i),
    .Q(\icache.itlb_icache_data_resp_i [7]),
    .QN(_26683_));
 DFF_X1 _60023_ (.D(\itlb.entry_ram.z_s1r1w_data_lo [14]),
    .CK(clk_i),
    .Q(\icache.itlb_icache_data_resp_i [8]),
    .QN(_26684_));
 DFF_X1 _60024_ (.D(\itlb.entry_ram.z_s1r1w_data_lo [15]),
    .CK(clk_i),
    .Q(\icache.itlb_icache_data_resp_i [9]),
    .QN(_26685_));
 DFF_X1 _60025_ (.D(\itlb.entry_ram.z_s1r1w_data_lo [16]),
    .CK(clk_i),
    .Q(\icache.itlb_icache_data_resp_i [10]),
    .QN(_26686_));
 DFF_X1 _60026_ (.D(\itlb.entry_ram.z_s1r1w_data_lo [17]),
    .CK(clk_i),
    .Q(\icache.itlb_icache_data_resp_i [11]),
    .QN(_26687_));
 DFF_X1 _60027_ (.D(\itlb.entry_ram.z_s1r1w_data_lo [18]),
    .CK(clk_i),
    .Q(\icache.itlb_icache_data_resp_i [12]),
    .QN(_26688_));
 DFF_X1 _60028_ (.D(\itlb.entry_ram.z_s1r1w_data_lo [19]),
    .CK(clk_i),
    .Q(\icache.itlb_icache_data_resp_i [13]),
    .QN(_26689_));
 DFF_X1 _60029_ (.D(\itlb.entry_ram.z_s1r1w_data_lo [20]),
    .CK(clk_i),
    .Q(\icache.itlb_icache_data_resp_i [14]),
    .QN(_26690_));
 DFF_X1 _60030_ (.D(\itlb.entry_ram.z_s1r1w_data_lo [21]),
    .CK(clk_i),
    .Q(\icache.itlb_icache_data_resp_i [15]),
    .QN(_26691_));
 DFF_X1 _60031_ (.D(\itlb.entry_ram.z_s1r1w_data_lo [22]),
    .CK(clk_i),
    .Q(\icache.itlb_icache_data_resp_i [16]),
    .QN(_26692_));
 DFF_X1 _60032_ (.D(\itlb.entry_ram.z_s1r1w_data_lo [23]),
    .CK(clk_i),
    .Q(\icache.itlb_icache_data_resp_i [17]),
    .QN(_26693_));
 DFF_X1 _60033_ (.D(\itlb.entry_ram.z_s1r1w_data_lo [24]),
    .CK(clk_i),
    .Q(\icache.itlb_icache_data_resp_i [18]),
    .QN(_26694_));
 DFF_X1 _60034_ (.D(\itlb.entry_ram.z_s1r1w_data_lo [25]),
    .CK(clk_i),
    .Q(\icache.itlb_icache_data_resp_i [19]),
    .QN(_26695_));
 DFF_X1 _60035_ (.D(\itlb.entry_ram.z_s1r1w_data_lo [26]),
    .CK(clk_i),
    .Q(\icache.itlb_icache_data_resp_i [20]),
    .QN(_26696_));
 DFF_X1 _60036_ (.D(\itlb.entry_ram.z_s1r1w_data_lo [27]),
    .CK(clk_i),
    .Q(\icache.itlb_icache_data_resp_i [21]),
    .QN(_26697_));
 DFF_X1 _60037_ (.D(\itlb.entry_ram.z_s1r1w_data_lo [28]),
    .CK(clk_i),
    .Q(\icache.itlb_icache_data_resp_i [22]),
    .QN(_26698_));
 DFF_X1 _60038_ (.D(\itlb.entry_ram.z_s1r1w_data_lo [29]),
    .CK(clk_i),
    .Q(\icache.itlb_icache_data_resp_i [23]),
    .QN(_26699_));
 DFF_X1 _60039_ (.D(\itlb.entry_ram.z_s1r1w_data_lo [30]),
    .CK(clk_i),
    .Q(\icache.itlb_icache_data_resp_i [24]),
    .QN(_26700_));
 DFF_X1 _60040_ (.D(\itlb.entry_ram.z_s1r1w_data_lo [31]),
    .CK(clk_i),
    .Q(\icache.itlb_icache_data_resp_i [25]),
    .QN(_26701_));
 DFF_X1 _60041_ (.D(\itlb.entry_ram.z_s1r1w_data_lo [32]),
    .CK(clk_i),
    .Q(\icache.itlb_icache_data_resp_i [26]),
    .QN(_26702_));
 DFF_X1 _60042_ (.D(_06817_),
    .CK(clk_i),
    .Q(\itlb.plru.encoder.N1 ),
    .QN(_00582_));
 DFF_X1 _60043_ (.D(_06818_),
    .CK(clk_i),
    .Q(\itlb.plru.encoder.lru_i [1]),
    .QN(_00576_));
 DFF_X1 _60044_ (.D(_06819_),
    .CK(clk_i),
    .Q(\itlb.plru.encoder.lru_i [2]),
    .QN(_00577_));
 DFF_X1 _60045_ (.D(_06820_),
    .CK(clk_i),
    .Q(\itlb.plru.encoder.lru_i [3]),
    .QN(_00578_));
 DFF_X1 _60046_ (.D(_06821_),
    .CK(clk_i),
    .Q(\itlb.plru.encoder.lru_i [4]),
    .QN(_00579_));
 DFF_X1 _60047_ (.D(_06822_),
    .CK(clk_i),
    .Q(\itlb.plru.encoder.lru_i [5]),
    .QN(_00580_));
 DFF_X1 _60048_ (.D(_06823_),
    .CK(clk_i),
    .Q(\itlb.plru.encoder.lru_i [6]),
    .QN(_00581_));
 DFF_X1 _60049_ (.D(_07040_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.valid [0]),
    .QN(_26703_));
 DFF_X1 _60050_ (.D(_07041_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.valid [1]),
    .QN(_26704_));
 DFF_X1 _60051_ (.D(_07042_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.valid [2]),
    .QN(_26705_));
 DFF_X1 _60052_ (.D(_07043_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.valid [3]),
    .QN(_26706_));
 DFF_X1 _60053_ (.D(_07044_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.valid [4]),
    .QN(_26707_));
 DFF_X1 _60054_ (.D(_07045_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.valid [5]),
    .QN(_26708_));
 DFF_X1 _60055_ (.D(_07046_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.valid [6]),
    .QN(_26709_));
 DFF_X1 _60056_ (.D(_07047_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.valid [7]),
    .QN(_26710_));
 DFF_X1 _60057_ (.D(_06824_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [0]),
    .QN(_26711_));
 DFF_X1 _60058_ (.D(_06935_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [1]),
    .QN(_26712_));
 DFF_X1 _60059_ (.D(_06962_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [2]),
    .QN(_26713_));
 DFF_X1 _60060_ (.D(_06973_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [3]),
    .QN(_26714_));
 DFF_X1 _60061_ (.D(_06984_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [4]),
    .QN(_26715_));
 DFF_X1 _60062_ (.D(_06995_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [5]),
    .QN(_26716_));
 DFF_X1 _60063_ (.D(_07006_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [6]),
    .QN(_26717_));
 DFF_X1 _60064_ (.D(_07017_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [7]),
    .QN(_26718_));
 DFF_X1 _60065_ (.D(_07028_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [8]),
    .QN(_26719_));
 DFF_X1 _60066_ (.D(_07039_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [9]),
    .QN(_26720_));
 DFF_X1 _60067_ (.D(_06835_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [10]),
    .QN(_26721_));
 DFF_X1 _60068_ (.D(_06846_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [11]),
    .QN(_26722_));
 DFF_X1 _60069_ (.D(_06857_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [12]),
    .QN(_26723_));
 DFF_X1 _60070_ (.D(_06868_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [13]),
    .QN(_26724_));
 DFF_X1 _60071_ (.D(_06879_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [14]),
    .QN(_26725_));
 DFF_X1 _60072_ (.D(_06890_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [15]),
    .QN(_26726_));
 DFF_X1 _60073_ (.D(_06901_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [16]),
    .QN(_26727_));
 DFF_X1 _60074_ (.D(_06912_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [17]),
    .QN(_26728_));
 DFF_X1 _60075_ (.D(_06923_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [18]),
    .QN(_26729_));
 DFF_X1 _60076_ (.D(_06934_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [19]),
    .QN(_26730_));
 DFF_X1 _60077_ (.D(_06946_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [20]),
    .QN(_26731_));
 DFF_X1 _60078_ (.D(_06953_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [21]),
    .QN(_26732_));
 DFF_X1 _60079_ (.D(_06954_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [22]),
    .QN(_26733_));
 DFF_X1 _60080_ (.D(_06955_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [23]),
    .QN(_26734_));
 DFF_X1 _60081_ (.D(_06956_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [24]),
    .QN(_26735_));
 DFF_X1 _60082_ (.D(_06957_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [25]),
    .QN(_26736_));
 DFF_X1 _60083_ (.D(_06958_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [26]),
    .QN(_26737_));
 DFF_X1 _60084_ (.D(_06959_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [27]),
    .QN(_26738_));
 DFF_X1 _60085_ (.D(_06960_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [28]),
    .QN(_26739_));
 DFF_X1 _60086_ (.D(_06961_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [29]),
    .QN(_26740_));
 DFF_X1 _60087_ (.D(_06963_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [30]),
    .QN(_26741_));
 DFF_X1 _60088_ (.D(_06964_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [31]),
    .QN(_26742_));
 DFF_X1 _60089_ (.D(_06965_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [32]),
    .QN(_26743_));
 DFF_X1 _60090_ (.D(_06966_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [33]),
    .QN(_26744_));
 DFF_X1 _60091_ (.D(_06967_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [34]),
    .QN(_26745_));
 DFF_X1 _60092_ (.D(_06968_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [35]),
    .QN(_26746_));
 DFF_X1 _60093_ (.D(_06969_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [36]),
    .QN(_26747_));
 DFF_X1 _60094_ (.D(_06970_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [37]),
    .QN(_26748_));
 DFF_X1 _60095_ (.D(_06971_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [38]),
    .QN(_26749_));
 DFF_X1 _60096_ (.D(_06972_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [39]),
    .QN(_26750_));
 DFF_X1 _60097_ (.D(_06974_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [40]),
    .QN(_26751_));
 DFF_X1 _60098_ (.D(_06975_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [41]),
    .QN(_26752_));
 DFF_X1 _60099_ (.D(_06976_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [42]),
    .QN(_26753_));
 DFF_X1 _60100_ (.D(_06977_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [43]),
    .QN(_26754_));
 DFF_X1 _60101_ (.D(_06978_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [44]),
    .QN(_26755_));
 DFF_X1 _60102_ (.D(_06979_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [45]),
    .QN(_26756_));
 DFF_X1 _60103_ (.D(_06980_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [46]),
    .QN(_26757_));
 DFF_X1 _60104_ (.D(_06981_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [47]),
    .QN(_26758_));
 DFF_X1 _60105_ (.D(_06982_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [48]),
    .QN(_26759_));
 DFF_X1 _60106_ (.D(_06983_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [49]),
    .QN(_26760_));
 DFF_X1 _60107_ (.D(_06985_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [50]),
    .QN(_26761_));
 DFF_X1 _60108_ (.D(_06986_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [51]),
    .QN(_26762_));
 DFF_X1 _60109_ (.D(_06987_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [52]),
    .QN(_26763_));
 DFF_X1 _60110_ (.D(_06988_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [53]),
    .QN(_26764_));
 DFF_X1 _60111_ (.D(_06989_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [54]),
    .QN(_26765_));
 DFF_X1 _60112_ (.D(_06990_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [55]),
    .QN(_26766_));
 DFF_X1 _60113_ (.D(_06991_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [56]),
    .QN(_26767_));
 DFF_X1 _60114_ (.D(_06992_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [57]),
    .QN(_26768_));
 DFF_X1 _60115_ (.D(_06993_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [58]),
    .QN(_26769_));
 DFF_X1 _60116_ (.D(_06994_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [59]),
    .QN(_26770_));
 DFF_X1 _60117_ (.D(_06996_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [60]),
    .QN(_26771_));
 DFF_X1 _60118_ (.D(_06997_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [61]),
    .QN(_26772_));
 DFF_X1 _60119_ (.D(_06998_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [62]),
    .QN(_26773_));
 DFF_X1 _60120_ (.D(_06999_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [63]),
    .QN(_26774_));
 DFF_X1 _60121_ (.D(_07000_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [64]),
    .QN(_26775_));
 DFF_X1 _60122_ (.D(_07001_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [65]),
    .QN(_26776_));
 DFF_X1 _60123_ (.D(_07002_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [66]),
    .QN(_26777_));
 DFF_X1 _60124_ (.D(_07003_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [67]),
    .QN(_26778_));
 DFF_X1 _60125_ (.D(_07004_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [68]),
    .QN(_26779_));
 DFF_X1 _60126_ (.D(_07005_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [69]),
    .QN(_26780_));
 DFF_X1 _60127_ (.D(_07007_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [70]),
    .QN(_26781_));
 DFF_X1 _60128_ (.D(_07008_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [71]),
    .QN(_26782_));
 DFF_X1 _60129_ (.D(_07009_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [72]),
    .QN(_26783_));
 DFF_X1 _60130_ (.D(_07010_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [73]),
    .QN(_26784_));
 DFF_X1 _60131_ (.D(_07011_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [74]),
    .QN(_26785_));
 DFF_X1 _60132_ (.D(_07012_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [75]),
    .QN(_26786_));
 DFF_X1 _60133_ (.D(_07013_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [76]),
    .QN(_26787_));
 DFF_X1 _60134_ (.D(_07014_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [77]),
    .QN(_26788_));
 DFF_X1 _60135_ (.D(_07015_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [78]),
    .QN(_26789_));
 DFF_X1 _60136_ (.D(_07016_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [79]),
    .QN(_26790_));
 DFF_X1 _60137_ (.D(_07018_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [80]),
    .QN(_26791_));
 DFF_X1 _60138_ (.D(_07019_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [81]),
    .QN(_26792_));
 DFF_X1 _60139_ (.D(_07020_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [82]),
    .QN(_26793_));
 DFF_X1 _60140_ (.D(_07021_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [83]),
    .QN(_26794_));
 DFF_X1 _60141_ (.D(_07022_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [84]),
    .QN(_26795_));
 DFF_X1 _60142_ (.D(_07023_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [85]),
    .QN(_26796_));
 DFF_X1 _60143_ (.D(_07024_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [86]),
    .QN(_26797_));
 DFF_X1 _60144_ (.D(_07025_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [87]),
    .QN(_26798_));
 DFF_X1 _60145_ (.D(_07026_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [88]),
    .QN(_26799_));
 DFF_X1 _60146_ (.D(_07027_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [89]),
    .QN(_26800_));
 DFF_X1 _60147_ (.D(_07029_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [90]),
    .QN(_26801_));
 DFF_X1 _60148_ (.D(_07030_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [91]),
    .QN(_26802_));
 DFF_X1 _60149_ (.D(_07031_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [92]),
    .QN(_26803_));
 DFF_X1 _60150_ (.D(_07032_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [93]),
    .QN(_26804_));
 DFF_X1 _60151_ (.D(_07033_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [94]),
    .QN(_26805_));
 DFF_X1 _60152_ (.D(_07034_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [95]),
    .QN(_26806_));
 DFF_X1 _60153_ (.D(_07035_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [96]),
    .QN(_26807_));
 DFF_X1 _60154_ (.D(_07036_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [97]),
    .QN(_26808_));
 DFF_X1 _60155_ (.D(_07037_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [98]),
    .QN(_26809_));
 DFF_X1 _60156_ (.D(_07038_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [99]),
    .QN(_26810_));
 DFF_X1 _60157_ (.D(_06825_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [100]),
    .QN(_26811_));
 DFF_X1 _60158_ (.D(_06826_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [101]),
    .QN(_26812_));
 DFF_X1 _60159_ (.D(_06827_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [102]),
    .QN(_26813_));
 DFF_X1 _60160_ (.D(_06828_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [103]),
    .QN(_26814_));
 DFF_X1 _60161_ (.D(_06829_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [104]),
    .QN(_26815_));
 DFF_X1 _60162_ (.D(_06830_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [105]),
    .QN(_26816_));
 DFF_X1 _60163_ (.D(_06831_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [106]),
    .QN(_26817_));
 DFF_X1 _60164_ (.D(_06832_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [107]),
    .QN(_26818_));
 DFF_X1 _60165_ (.D(_06833_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [108]),
    .QN(_26819_));
 DFF_X1 _60166_ (.D(_06834_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [109]),
    .QN(_26820_));
 DFF_X1 _60167_ (.D(_06836_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [110]),
    .QN(_26821_));
 DFF_X1 _60168_ (.D(_06837_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [111]),
    .QN(_26822_));
 DFF_X1 _60169_ (.D(_06838_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [112]),
    .QN(_26823_));
 DFF_X1 _60170_ (.D(_06839_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [113]),
    .QN(_26824_));
 DFF_X1 _60171_ (.D(_06840_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [114]),
    .QN(_26825_));
 DFF_X1 _60172_ (.D(_06841_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [115]),
    .QN(_26826_));
 DFF_X1 _60173_ (.D(_06842_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [116]),
    .QN(_26827_));
 DFF_X1 _60174_ (.D(_06843_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [117]),
    .QN(_26828_));
 DFF_X1 _60175_ (.D(_06844_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [118]),
    .QN(_26829_));
 DFF_X1 _60176_ (.D(_06845_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [119]),
    .QN(_26830_));
 DFF_X1 _60177_ (.D(_06847_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [120]),
    .QN(_26831_));
 DFF_X1 _60178_ (.D(_06848_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [121]),
    .QN(_26832_));
 DFF_X1 _60179_ (.D(_06849_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [122]),
    .QN(_26833_));
 DFF_X1 _60180_ (.D(_06850_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [123]),
    .QN(_26834_));
 DFF_X1 _60181_ (.D(_06851_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [124]),
    .QN(_26835_));
 DFF_X1 _60182_ (.D(_06852_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [125]),
    .QN(_26836_));
 DFF_X1 _60183_ (.D(_06853_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [126]),
    .QN(_26837_));
 DFF_X1 _60184_ (.D(_06854_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [127]),
    .QN(_26838_));
 DFF_X1 _60185_ (.D(_06855_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [128]),
    .QN(_26839_));
 DFF_X1 _60186_ (.D(_06856_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [129]),
    .QN(_26840_));
 DFF_X1 _60187_ (.D(_06858_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [130]),
    .QN(_26841_));
 DFF_X1 _60188_ (.D(_06859_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [131]),
    .QN(_26842_));
 DFF_X1 _60189_ (.D(_06860_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [132]),
    .QN(_26843_));
 DFF_X1 _60190_ (.D(_06861_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [133]),
    .QN(_26844_));
 DFF_X1 _60191_ (.D(_06862_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [134]),
    .QN(_26845_));
 DFF_X1 _60192_ (.D(_06863_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [135]),
    .QN(_26846_));
 DFF_X1 _60193_ (.D(_06864_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [136]),
    .QN(_26847_));
 DFF_X1 _60194_ (.D(_06865_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [137]),
    .QN(_26848_));
 DFF_X1 _60195_ (.D(_06866_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [138]),
    .QN(_26849_));
 DFF_X1 _60196_ (.D(_06867_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [139]),
    .QN(_26850_));
 DFF_X1 _60197_ (.D(_06869_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [140]),
    .QN(_26851_));
 DFF_X1 _60198_ (.D(_06870_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [141]),
    .QN(_26852_));
 DFF_X1 _60199_ (.D(_06871_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [142]),
    .QN(_26853_));
 DFF_X1 _60200_ (.D(_06872_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [143]),
    .QN(_26854_));
 DFF_X1 _60201_ (.D(_06873_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [144]),
    .QN(_26855_));
 DFF_X1 _60202_ (.D(_06874_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [145]),
    .QN(_26856_));
 DFF_X1 _60203_ (.D(_06875_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [146]),
    .QN(_26857_));
 DFF_X1 _60204_ (.D(_06876_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [147]),
    .QN(_26858_));
 DFF_X1 _60205_ (.D(_06877_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [148]),
    .QN(_26859_));
 DFF_X1 _60206_ (.D(_06878_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [149]),
    .QN(_26860_));
 DFF_X1 _60207_ (.D(_06880_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [150]),
    .QN(_26861_));
 DFF_X1 _60208_ (.D(_06881_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [151]),
    .QN(_26862_));
 DFF_X1 _60209_ (.D(_06882_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [152]),
    .QN(_26863_));
 DFF_X1 _60210_ (.D(_06883_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [153]),
    .QN(_26864_));
 DFF_X1 _60211_ (.D(_06884_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [154]),
    .QN(_26865_));
 DFF_X1 _60212_ (.D(_06885_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [155]),
    .QN(_26866_));
 DFF_X1 _60213_ (.D(_06886_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [156]),
    .QN(_26867_));
 DFF_X1 _60214_ (.D(_06887_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [157]),
    .QN(_26868_));
 DFF_X1 _60215_ (.D(_06888_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [158]),
    .QN(_26869_));
 DFF_X1 _60216_ (.D(_06889_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [159]),
    .QN(_26870_));
 DFF_X1 _60217_ (.D(_06891_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [160]),
    .QN(_26871_));
 DFF_X1 _60218_ (.D(_06892_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [161]),
    .QN(_26872_));
 DFF_X1 _60219_ (.D(_06893_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [162]),
    .QN(_26873_));
 DFF_X1 _60220_ (.D(_06894_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [163]),
    .QN(_26874_));
 DFF_X1 _60221_ (.D(_06895_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [164]),
    .QN(_26875_));
 DFF_X1 _60222_ (.D(_06896_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [165]),
    .QN(_26876_));
 DFF_X1 _60223_ (.D(_06897_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [166]),
    .QN(_26877_));
 DFF_X1 _60224_ (.D(_06898_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [167]),
    .QN(_26878_));
 DFF_X1 _60225_ (.D(_06899_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [168]),
    .QN(_26879_));
 DFF_X1 _60226_ (.D(_06900_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [169]),
    .QN(_26880_));
 DFF_X1 _60227_ (.D(_06902_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [170]),
    .QN(_26881_));
 DFF_X1 _60228_ (.D(_06903_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [171]),
    .QN(_26882_));
 DFF_X1 _60229_ (.D(_06904_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [172]),
    .QN(_26883_));
 DFF_X1 _60230_ (.D(_06905_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [173]),
    .QN(_26884_));
 DFF_X1 _60231_ (.D(_06906_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [174]),
    .QN(_26885_));
 DFF_X1 _60232_ (.D(_06907_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [175]),
    .QN(_26886_));
 DFF_X1 _60233_ (.D(_06908_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [176]),
    .QN(_26887_));
 DFF_X1 _60234_ (.D(_06909_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [177]),
    .QN(_26888_));
 DFF_X1 _60235_ (.D(_06910_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [178]),
    .QN(_26889_));
 DFF_X1 _60236_ (.D(_06911_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [179]),
    .QN(_26890_));
 DFF_X1 _60237_ (.D(_06913_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [180]),
    .QN(_26891_));
 DFF_X1 _60238_ (.D(_06914_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [181]),
    .QN(_26892_));
 DFF_X1 _60239_ (.D(_06915_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [182]),
    .QN(_26893_));
 DFF_X1 _60240_ (.D(_06916_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [183]),
    .QN(_26894_));
 DFF_X1 _60241_ (.D(_06917_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [184]),
    .QN(_26895_));
 DFF_X1 _60242_ (.D(_06918_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [185]),
    .QN(_26896_));
 DFF_X1 _60243_ (.D(_06919_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [186]),
    .QN(_26897_));
 DFF_X1 _60244_ (.D(_06920_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [187]),
    .QN(_26898_));
 DFF_X1 _60245_ (.D(_06921_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [188]),
    .QN(_26899_));
 DFF_X1 _60246_ (.D(_06922_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [189]),
    .QN(_26900_));
 DFF_X1 _60247_ (.D(_06924_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [190]),
    .QN(_26901_));
 DFF_X1 _60248_ (.D(_06925_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [191]),
    .QN(_26902_));
 DFF_X1 _60249_ (.D(_06926_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [192]),
    .QN(_26903_));
 DFF_X1 _60250_ (.D(_06927_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [193]),
    .QN(_26904_));
 DFF_X1 _60251_ (.D(_06928_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [194]),
    .QN(_26905_));
 DFF_X1 _60252_ (.D(_06929_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [195]),
    .QN(_26906_));
 DFF_X1 _60253_ (.D(_06930_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [196]),
    .QN(_26907_));
 DFF_X1 _60254_ (.D(_06931_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [197]),
    .QN(_26908_));
 DFF_X1 _60255_ (.D(_06932_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [198]),
    .QN(_26909_));
 DFF_X1 _60256_ (.D(_06933_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [199]),
    .QN(_26910_));
 DFF_X1 _60257_ (.D(_06936_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [200]),
    .QN(_26911_));
 DFF_X1 _60258_ (.D(_06937_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [201]),
    .QN(_26912_));
 DFF_X1 _60259_ (.D(_06938_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [202]),
    .QN(_26913_));
 DFF_X1 _60260_ (.D(_06939_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [203]),
    .QN(_26914_));
 DFF_X1 _60261_ (.D(_06940_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [204]),
    .QN(_26915_));
 DFF_X1 _60262_ (.D(_06941_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [205]),
    .QN(_26916_));
 DFF_X1 _60263_ (.D(_06942_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [206]),
    .QN(_26917_));
 DFF_X1 _60264_ (.D(_06943_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [207]),
    .QN(_26918_));
 DFF_X1 _60265_ (.D(_06944_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [208]),
    .QN(_26919_));
 DFF_X1 _60266_ (.D(_06945_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [209]),
    .QN(_26920_));
 DFF_X1 _60267_ (.D(_06947_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [210]),
    .QN(_26921_));
 DFF_X1 _60268_ (.D(_06948_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [211]),
    .QN(_26922_));
 DFF_X1 _60269_ (.D(_06949_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [212]),
    .QN(_26923_));
 DFF_X1 _60270_ (.D(_06950_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [213]),
    .QN(_26924_));
 DFF_X1 _60271_ (.D(_06951_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [214]),
    .QN(_26925_));
 DFF_X1 _60272_ (.D(_06952_),
    .CK(clk_i),
    .Q(\itlb.vtag_cam.mem [215]),
    .QN(_26926_));
 DFF_X1 _60273_ (.D(\itlb.miss_v_reg.N3 ),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.itlb_miss_i ),
    .QN(_26927_));
 DFF_X1 _60274_ (.D(\itlb.r_v_reg.N3 ),
    .CK(clk_i),
    .Q(\icache.itlb_icache_data_resp_v_i ),
    .QN(_26928_));
 DFF_X1 _60275_ (.D(_04888_),
    .CK(clk_i),
    .Q(\icache.N7 ),
    .QN(_26929_));
 DFF_X1 _60276_ (.D(_00758_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [0]),
    .QN(_00006_));
 DFF_X1 _60277_ (.D(_00769_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [1]),
    .QN(_00007_));
 DFF_X1 _60278_ (.D(_00780_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [2]),
    .QN(_00008_));
 DFF_X1 _60279_ (.D(_00791_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [3]),
    .QN(_00009_));
 DFF_X1 _60280_ (.D(_00802_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [4]),
    .QN(_00010_));
 DFF_X1 _60281_ (.D(_00813_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [5]),
    .QN(_00011_));
 DFF_X1 _60282_ (.D(_00818_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [6]),
    .QN(_00012_));
 DFF_X1 _60283_ (.D(_00819_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [7]),
    .QN(_00013_));
 DFF_X1 _60284_ (.D(_00820_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [8]),
    .QN(_00014_));
 DFF_X1 _60285_ (.D(_00821_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [9]),
    .QN(_00015_));
 DFF_X1 _60286_ (.D(_00759_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [10]),
    .QN(_00016_));
 DFF_X1 _60287_ (.D(_00760_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [11]),
    .QN(_00017_));
 DFF_X1 _60288_ (.D(_00761_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [12]),
    .QN(_00018_));
 DFF_X1 _60289_ (.D(_00762_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [13]),
    .QN(_00019_));
 DFF_X1 _60290_ (.D(_00763_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [14]),
    .QN(_00020_));
 DFF_X1 _60291_ (.D(_00764_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [15]),
    .QN(_00021_));
 DFF_X1 _60292_ (.D(_00765_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [16]),
    .QN(_00022_));
 DFF_X1 _60293_ (.D(_00766_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [17]),
    .QN(_00023_));
 DFF_X1 _60294_ (.D(_00767_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [18]),
    .QN(_00024_));
 DFF_X1 _60295_ (.D(_00768_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [19]),
    .QN(_00025_));
 DFF_X1 _60296_ (.D(_00770_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [20]),
    .QN(_00026_));
 DFF_X1 _60297_ (.D(_00771_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [21]),
    .QN(_00027_));
 DFF_X1 _60298_ (.D(_00772_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [22]),
    .QN(_00028_));
 DFF_X1 _60299_ (.D(_00773_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [23]),
    .QN(_00029_));
 DFF_X1 _60300_ (.D(_00774_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [24]),
    .QN(_00030_));
 DFF_X1 _60301_ (.D(_00775_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [25]),
    .QN(_00031_));
 DFF_X1 _60302_ (.D(_00776_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [26]),
    .QN(_00032_));
 DFF_X1 _60303_ (.D(_00777_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [27]),
    .QN(_00033_));
 DFF_X1 _60304_ (.D(_00778_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [28]),
    .QN(_00034_));
 DFF_X1 _60305_ (.D(_00779_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [29]),
    .QN(_00035_));
 DFF_X1 _60306_ (.D(_00781_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [30]),
    .QN(_00036_));
 DFF_X1 _60307_ (.D(_00782_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [31]),
    .QN(_00037_));
 DFF_X1 _60308_ (.D(_00783_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [32]),
    .QN(_00038_));
 DFF_X1 _60309_ (.D(_00784_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [33]),
    .QN(_00039_));
 DFF_X1 _60310_ (.D(_00785_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [34]),
    .QN(_00040_));
 DFF_X1 _60311_ (.D(_00786_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [35]),
    .QN(_00041_));
 DFF_X1 _60312_ (.D(_00787_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [36]),
    .QN(_00042_));
 DFF_X1 _60313_ (.D(_00788_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [37]),
    .QN(_00043_));
 DFF_X1 _60314_ (.D(_00789_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [38]),
    .QN(_00044_));
 DFF_X1 _60315_ (.D(_00790_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [39]),
    .QN(_00045_));
 DFF_X1 _60316_ (.D(_00792_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [40]),
    .QN(_00046_));
 DFF_X1 _60317_ (.D(_00793_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [41]),
    .QN(_00047_));
 DFF_X1 _60318_ (.D(_00794_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [42]),
    .QN(_00048_));
 DFF_X1 _60319_ (.D(_00795_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [43]),
    .QN(_00049_));
 DFF_X1 _60320_ (.D(_00796_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [44]),
    .QN(_00050_));
 DFF_X1 _60321_ (.D(_00797_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [45]),
    .QN(_00051_));
 DFF_X1 _60322_ (.D(_00798_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [46]),
    .QN(_00052_));
 DFF_X1 _60323_ (.D(_00799_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [47]),
    .QN(_00053_));
 DFF_X1 _60324_ (.D(_00800_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [48]),
    .QN(_00054_));
 DFF_X1 _60325_ (.D(_00801_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [49]),
    .QN(_00055_));
 DFF_X1 _60326_ (.D(_00803_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [50]),
    .QN(_00056_));
 DFF_X1 _60327_ (.D(_00804_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [51]),
    .QN(_00057_));
 DFF_X1 _60328_ (.D(_00805_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [52]),
    .QN(_00058_));
 DFF_X1 _60329_ (.D(_00806_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [53]),
    .QN(_00059_));
 DFF_X1 _60330_ (.D(_00807_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [54]),
    .QN(_00060_));
 DFF_X1 _60331_ (.D(_00808_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [55]),
    .QN(_00061_));
 DFF_X1 _60332_ (.D(_00809_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [56]),
    .QN(_00062_));
 DFF_X1 _60333_ (.D(_00810_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [57]),
    .QN(_00063_));
 DFF_X1 _60334_ (.D(_00811_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [58]),
    .QN(_00064_));
 DFF_X1 _60335_ (.D(_00812_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [59]),
    .QN(_00065_));
 DFF_X1 _60336_ (.D(_00814_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [60]),
    .QN(_00066_));
 DFF_X1 _60337_ (.D(_00815_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [61]),
    .QN(_00067_));
 DFF_X1 _60338_ (.D(_00816_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [62]),
    .QN(_00068_));
 DFF_X1 _60339_ (.D(_00817_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.v_r [63]),
    .QN(_26930_));
 DFF_X1 _60340_ (.D(\bp_fe_pc_gen_1.btb.N150 ),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.r_tag_r [0]),
    .QN(_26931_));
 DFF_X1 _60341_ (.D(\bp_fe_pc_gen_1.btb.N151 ),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.r_tag_r [1]),
    .QN(_26932_));
 DFF_X1 _60342_ (.D(\bp_fe_pc_gen_1.btb.N152 ),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.r_tag_r [2]),
    .QN(_26933_));
 DFF_X1 _60343_ (.D(\bp_fe_pc_gen_1.btb.N153 ),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.r_tag_r [3]),
    .QN(_26934_));
 DFF_X1 _60344_ (.D(\bp_fe_pc_gen_1.btb.N154 ),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.r_tag_r [4]),
    .QN(_26935_));
 DFF_X1 _60345_ (.D(\bp_fe_pc_gen_1.btb.N155 ),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.r_tag_r [5]),
    .QN(_26936_));
 DFF_X1 _60346_ (.D(\bp_fe_pc_gen_1.btb.N156 ),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.r_tag_r [6]),
    .QN(_26937_));
 DFF_X1 _60347_ (.D(\bp_fe_pc_gen_1.btb.N157 ),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.r_tag_r [7]),
    .QN(_26938_));
 DFF_X1 _60348_ (.D(\bp_fe_pc_gen_1.btb.N158 ),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.r_tag_r [8]),
    .QN(_26939_));
 DFF_X1 _60349_ (.D(\bp_fe_pc_gen_1.btb.N159 ),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.r_tag_r [9]),
    .QN(_26940_));
 DFF_X1 _60350_ (.D(\bp_fe_pc_gen_1.btb.N149 ),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.r_v_r ),
    .QN(_26941_));
 DFF_X1 _60351_ (.D(\bp_fe_pc_gen_1.btb.N160 ),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.r_idx_r [0]),
    .QN(_26942_));
 DFF_X1 _60352_ (.D(\bp_fe_pc_gen_1.btb.N161 ),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.r_idx_r [1]),
    .QN(_26943_));
 DFF_X1 _60353_ (.D(\bp_fe_pc_gen_1.btb.N162 ),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.r_idx_r [2]),
    .QN(_00071_));
 DFF_X1 _60354_ (.D(\bp_fe_pc_gen_1.btb.N163 ),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.r_idx_r [3]),
    .QN(_00070_));
 DFF_X1 _60355_ (.D(\bp_fe_pc_gen_1.btb.N164 ),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.r_idx_r [4]),
    .QN(_00069_));
 DFF_X1 _60356_ (.D(\bp_fe_pc_gen_1.btb.N165 ),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.r_idx_r [5]),
    .QN(_00072_));
 DFF_X1 _60357_ (.D(_00731_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [0]),
    .QN(_26944_));
 DFF_X1 _60358_ (.D(_00742_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [1]),
    .QN(_26945_));
 DFF_X1 _60359_ (.D(_00750_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [2]),
    .QN(_26946_));
 DFF_X1 _60360_ (.D(_00751_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [3]),
    .QN(_26947_));
 DFF_X1 _60361_ (.D(_00752_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [4]),
    .QN(_26948_));
 DFF_X1 _60362_ (.D(_00753_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [5]),
    .QN(_26949_));
 DFF_X1 _60363_ (.D(_00754_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [6]),
    .QN(_26950_));
 DFF_X1 _60364_ (.D(_00755_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [7]),
    .QN(_26951_));
 DFF_X1 _60365_ (.D(_00756_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [8]),
    .QN(_26952_));
 DFF_X1 _60366_ (.D(_00757_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [9]),
    .QN(_26953_));
 DFF_X1 _60367_ (.D(_00732_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [10]),
    .QN(_26954_));
 DFF_X1 _60368_ (.D(_00733_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [11]),
    .QN(_26955_));
 DFF_X1 _60369_ (.D(_00734_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [12]),
    .QN(_26956_));
 DFF_X1 _60370_ (.D(_00735_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [13]),
    .QN(_26957_));
 DFF_X1 _60371_ (.D(_00736_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [14]),
    .QN(_26958_));
 DFF_X1 _60372_ (.D(_00737_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [15]),
    .QN(_26959_));
 DFF_X1 _60373_ (.D(_00738_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [16]),
    .QN(_26960_));
 DFF_X1 _60374_ (.D(_00739_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [17]),
    .QN(_26961_));
 DFF_X1 _60375_ (.D(_00740_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [18]),
    .QN(_26962_));
 DFF_X1 _60376_ (.D(_00741_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [19]),
    .QN(_26963_));
 DFF_X1 _60377_ (.D(_00743_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [20]),
    .QN(_26964_));
 DFF_X1 _60378_ (.D(_00744_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [21]),
    .QN(_26965_));
 DFF_X1 _60379_ (.D(_00745_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [22]),
    .QN(_26966_));
 DFF_X1 _60380_ (.D(_00746_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [23]),
    .QN(_26967_));
 DFF_X1 _60381_ (.D(_00747_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [24]),
    .QN(_26968_));
 DFF_X1 _60382_ (.D(_00748_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [25]),
    .QN(_26969_));
 DFF_X1 _60383_ (.D(_00749_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_o [26]),
    .QN(_26970_));
 DFF_X1 _60384_ (.D(_06592_),
    .CK(clk_i),
    .Q(\icache.lce.lce_req_inst.tr_data_received_r ),
    .QN(_00602_));
 DFF_X1 _60385_ (.D(_05402_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.N0 ),
    .QN(_00597_));
 DFF_X1 _60386_ (.D(_05401_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.N10 ),
    .QN(_26971_));
 DFF_X1 _60387_ (.D(_05405_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.syn_ack_cnt_r ),
    .QN(_00600_));
 DFF_X1 _60388_ (.D(_04889_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [0]),
    .QN(_26972_));
 DFF_X1 _60389_ (.D(_05000_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [1]),
    .QN(_26973_));
 DFF_X1 _60390_ (.D(_05111_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [2]),
    .QN(_26974_));
 DFF_X1 _60391_ (.D(_05222_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [3]),
    .QN(_26975_));
 DFF_X1 _60392_ (.D(_05333_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [4]),
    .QN(_26976_));
 DFF_X1 _60393_ (.D(_05356_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [5]),
    .QN(_26977_));
 DFF_X1 _60394_ (.D(_05367_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [6]),
    .QN(_26978_));
 DFF_X1 _60395_ (.D(_05378_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [7]),
    .QN(_26979_));
 DFF_X1 _60396_ (.D(_05389_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [8]),
    .QN(_26980_));
 DFF_X1 _60397_ (.D(_05400_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [9]),
    .QN(_26981_));
 DFF_X1 _60398_ (.D(_04900_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [10]),
    .QN(_26982_));
 DFF_X1 _60399_ (.D(_04911_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [11]),
    .QN(_26983_));
 DFF_X1 _60400_ (.D(_04922_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [12]),
    .QN(_26984_));
 DFF_X1 _60401_ (.D(_04933_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [13]),
    .QN(_26985_));
 DFF_X1 _60402_ (.D(_04944_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [14]),
    .QN(_26986_));
 DFF_X1 _60403_ (.D(_04955_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [15]),
    .QN(_26987_));
 DFF_X1 _60404_ (.D(_04966_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [16]),
    .QN(_26988_));
 DFF_X1 _60405_ (.D(_04977_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [17]),
    .QN(_26989_));
 DFF_X1 _60406_ (.D(_04988_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [18]),
    .QN(_26990_));
 DFF_X1 _60407_ (.D(_04999_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [19]),
    .QN(_26991_));
 DFF_X1 _60408_ (.D(_05011_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [20]),
    .QN(_26992_));
 DFF_X1 _60409_ (.D(_05022_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [21]),
    .QN(_26993_));
 DFF_X1 _60410_ (.D(_05033_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [22]),
    .QN(_26994_));
 DFF_X1 _60411_ (.D(_05044_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [23]),
    .QN(_26995_));
 DFF_X1 _60412_ (.D(_05055_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [24]),
    .QN(_26996_));
 DFF_X1 _60413_ (.D(_05066_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [25]),
    .QN(_26997_));
 DFF_X1 _60414_ (.D(_05077_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [26]),
    .QN(_26998_));
 DFF_X1 _60415_ (.D(_05088_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [27]),
    .QN(_26999_));
 DFF_X1 _60416_ (.D(_05099_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [28]),
    .QN(_27000_));
 DFF_X1 _60417_ (.D(_05110_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [29]),
    .QN(_27001_));
 DFF_X1 _60418_ (.D(_05122_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [30]),
    .QN(_27002_));
 DFF_X1 _60419_ (.D(_05133_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [31]),
    .QN(_27003_));
 DFF_X1 _60420_ (.D(_05144_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [32]),
    .QN(_27004_));
 DFF_X1 _60421_ (.D(_05155_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [33]),
    .QN(_27005_));
 DFF_X1 _60422_ (.D(_05166_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [34]),
    .QN(_27006_));
 DFF_X1 _60423_ (.D(_05177_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [35]),
    .QN(_27007_));
 DFF_X1 _60424_ (.D(_05188_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [36]),
    .QN(_27008_));
 DFF_X1 _60425_ (.D(_05199_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [37]),
    .QN(_27009_));
 DFF_X1 _60426_ (.D(_05210_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [38]),
    .QN(_27010_));
 DFF_X1 _60427_ (.D(_05221_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [39]),
    .QN(_27011_));
 DFF_X1 _60428_ (.D(_05233_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [40]),
    .QN(_27012_));
 DFF_X1 _60429_ (.D(_05244_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [41]),
    .QN(_27013_));
 DFF_X1 _60430_ (.D(_05255_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [42]),
    .QN(_27014_));
 DFF_X1 _60431_ (.D(_05266_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [43]),
    .QN(_27015_));
 DFF_X1 _60432_ (.D(_05277_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [44]),
    .QN(_27016_));
 DFF_X1 _60433_ (.D(_05288_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [45]),
    .QN(_27017_));
 DFF_X1 _60434_ (.D(_05299_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [46]),
    .QN(_27018_));
 DFF_X1 _60435_ (.D(_05310_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [47]),
    .QN(_27019_));
 DFF_X1 _60436_ (.D(_05321_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [48]),
    .QN(_27020_));
 DFF_X1 _60437_ (.D(_05332_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [49]),
    .QN(_27021_));
 DFF_X1 _60438_ (.D(_05344_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [50]),
    .QN(_27022_));
 DFF_X1 _60439_ (.D(_05347_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [51]),
    .QN(_27023_));
 DFF_X1 _60440_ (.D(_05348_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [52]),
    .QN(_27024_));
 DFF_X1 _60441_ (.D(_05349_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [53]),
    .QN(_27025_));
 DFF_X1 _60442_ (.D(_05350_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [54]),
    .QN(_27026_));
 DFF_X1 _60443_ (.D(_05351_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [55]),
    .QN(_27027_));
 DFF_X1 _60444_ (.D(_05352_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [56]),
    .QN(_27028_));
 DFF_X1 _60445_ (.D(_05353_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [57]),
    .QN(_27029_));
 DFF_X1 _60446_ (.D(_05354_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [58]),
    .QN(_27030_));
 DFF_X1 _60447_ (.D(_05355_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [59]),
    .QN(_27031_));
 DFF_X1 _60448_ (.D(_05357_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [60]),
    .QN(_27032_));
 DFF_X1 _60449_ (.D(_05358_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [61]),
    .QN(_27033_));
 DFF_X1 _60450_ (.D(_05359_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [62]),
    .QN(_27034_));
 DFF_X1 _60451_ (.D(_05360_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [63]),
    .QN(_27035_));
 DFF_X1 _60452_ (.D(_05361_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [64]),
    .QN(_27036_));
 DFF_X1 _60453_ (.D(_05362_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [65]),
    .QN(_27037_));
 DFF_X1 _60454_ (.D(_05363_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [66]),
    .QN(_27038_));
 DFF_X1 _60455_ (.D(_05364_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [67]),
    .QN(_27039_));
 DFF_X1 _60456_ (.D(_05365_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [68]),
    .QN(_27040_));
 DFF_X1 _60457_ (.D(_05366_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [69]),
    .QN(_27041_));
 DFF_X1 _60458_ (.D(_05368_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [70]),
    .QN(_27042_));
 DFF_X1 _60459_ (.D(_05369_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [71]),
    .QN(_27043_));
 DFF_X1 _60460_ (.D(_05370_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [72]),
    .QN(_27044_));
 DFF_X1 _60461_ (.D(_05371_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [73]),
    .QN(_27045_));
 DFF_X1 _60462_ (.D(_05372_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [74]),
    .QN(_27046_));
 DFF_X1 _60463_ (.D(_05373_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [75]),
    .QN(_27047_));
 DFF_X1 _60464_ (.D(_05374_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [76]),
    .QN(_27048_));
 DFF_X1 _60465_ (.D(_05375_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [77]),
    .QN(_27049_));
 DFF_X1 _60466_ (.D(_05376_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [78]),
    .QN(_27050_));
 DFF_X1 _60467_ (.D(_05377_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [79]),
    .QN(_27051_));
 DFF_X1 _60468_ (.D(_05379_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [80]),
    .QN(_27052_));
 DFF_X1 _60469_ (.D(_05380_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [81]),
    .QN(_27053_));
 DFF_X1 _60470_ (.D(_05381_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [82]),
    .QN(_27054_));
 DFF_X1 _60471_ (.D(_05382_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [83]),
    .QN(_27055_));
 DFF_X1 _60472_ (.D(_05383_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [84]),
    .QN(_27056_));
 DFF_X1 _60473_ (.D(_05384_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [85]),
    .QN(_27057_));
 DFF_X1 _60474_ (.D(_05385_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [86]),
    .QN(_27058_));
 DFF_X1 _60475_ (.D(_05386_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [87]),
    .QN(_27059_));
 DFF_X1 _60476_ (.D(_05387_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [88]),
    .QN(_27060_));
 DFF_X1 _60477_ (.D(_05388_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [89]),
    .QN(_27061_));
 DFF_X1 _60478_ (.D(_05390_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [90]),
    .QN(_27062_));
 DFF_X1 _60479_ (.D(_05391_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [91]),
    .QN(_27063_));
 DFF_X1 _60480_ (.D(_05392_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [92]),
    .QN(_27064_));
 DFF_X1 _60481_ (.D(_05393_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [93]),
    .QN(_27065_));
 DFF_X1 _60482_ (.D(_05394_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [94]),
    .QN(_27066_));
 DFF_X1 _60483_ (.D(_05395_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [95]),
    .QN(_27067_));
 DFF_X1 _60484_ (.D(_05396_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [96]),
    .QN(_27068_));
 DFF_X1 _60485_ (.D(_05397_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [97]),
    .QN(_27069_));
 DFF_X1 _60486_ (.D(_05398_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [98]),
    .QN(_27070_));
 DFF_X1 _60487_ (.D(_05399_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [99]),
    .QN(_27071_));
 DFF_X1 _60488_ (.D(_04890_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [100]),
    .QN(_27072_));
 DFF_X1 _60489_ (.D(_04891_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [101]),
    .QN(_27073_));
 DFF_X1 _60490_ (.D(_04892_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [102]),
    .QN(_27074_));
 DFF_X1 _60491_ (.D(_04893_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [103]),
    .QN(_27075_));
 DFF_X1 _60492_ (.D(_04894_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [104]),
    .QN(_27076_));
 DFF_X1 _60493_ (.D(_04895_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [105]),
    .QN(_27077_));
 DFF_X1 _60494_ (.D(_04896_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [106]),
    .QN(_27078_));
 DFF_X1 _60495_ (.D(_04897_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [107]),
    .QN(_27079_));
 DFF_X1 _60496_ (.D(_04898_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [108]),
    .QN(_27080_));
 DFF_X1 _60497_ (.D(_04899_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [109]),
    .QN(_27081_));
 DFF_X1 _60498_ (.D(_04901_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [110]),
    .QN(_27082_));
 DFF_X1 _60499_ (.D(_04902_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [111]),
    .QN(_27083_));
 DFF_X1 _60500_ (.D(_04903_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [112]),
    .QN(_27084_));
 DFF_X1 _60501_ (.D(_04904_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [113]),
    .QN(_27085_));
 DFF_X1 _60502_ (.D(_04905_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [114]),
    .QN(_27086_));
 DFF_X1 _60503_ (.D(_04906_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [115]),
    .QN(_27087_));
 DFF_X1 _60504_ (.D(_04907_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [116]),
    .QN(_27088_));
 DFF_X1 _60505_ (.D(_04908_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [117]),
    .QN(_27089_));
 DFF_X1 _60506_ (.D(_04909_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [118]),
    .QN(_27090_));
 DFF_X1 _60507_ (.D(_04910_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [119]),
    .QN(_27091_));
 DFF_X1 _60508_ (.D(_04912_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [120]),
    .QN(_27092_));
 DFF_X1 _60509_ (.D(_04913_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [121]),
    .QN(_27093_));
 DFF_X1 _60510_ (.D(_04914_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [122]),
    .QN(_27094_));
 DFF_X1 _60511_ (.D(_04915_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [123]),
    .QN(_27095_));
 DFF_X1 _60512_ (.D(_04916_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [124]),
    .QN(_27096_));
 DFF_X1 _60513_ (.D(_04917_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [125]),
    .QN(_27097_));
 DFF_X1 _60514_ (.D(_04918_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [126]),
    .QN(_27098_));
 DFF_X1 _60515_ (.D(_04919_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [127]),
    .QN(_27099_));
 DFF_X1 _60516_ (.D(_04920_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [128]),
    .QN(_27100_));
 DFF_X1 _60517_ (.D(_04921_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [129]),
    .QN(_27101_));
 DFF_X1 _60518_ (.D(_04923_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [130]),
    .QN(_27102_));
 DFF_X1 _60519_ (.D(_04924_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [131]),
    .QN(_27103_));
 DFF_X1 _60520_ (.D(_04925_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [132]),
    .QN(_27104_));
 DFF_X1 _60521_ (.D(_04926_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [133]),
    .QN(_27105_));
 DFF_X1 _60522_ (.D(_04927_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [134]),
    .QN(_27106_));
 DFF_X1 _60523_ (.D(_04928_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [135]),
    .QN(_27107_));
 DFF_X1 _60524_ (.D(_04929_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [136]),
    .QN(_27108_));
 DFF_X1 _60525_ (.D(_04930_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [137]),
    .QN(_27109_));
 DFF_X1 _60526_ (.D(_04931_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [138]),
    .QN(_27110_));
 DFF_X1 _60527_ (.D(_04932_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [139]),
    .QN(_27111_));
 DFF_X1 _60528_ (.D(_04934_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [140]),
    .QN(_27112_));
 DFF_X1 _60529_ (.D(_04935_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [141]),
    .QN(_27113_));
 DFF_X1 _60530_ (.D(_04936_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [142]),
    .QN(_27114_));
 DFF_X1 _60531_ (.D(_04937_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [143]),
    .QN(_27115_));
 DFF_X1 _60532_ (.D(_04938_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [144]),
    .QN(_27116_));
 DFF_X1 _60533_ (.D(_04939_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [145]),
    .QN(_27117_));
 DFF_X1 _60534_ (.D(_04940_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [146]),
    .QN(_27118_));
 DFF_X1 _60535_ (.D(_04941_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [147]),
    .QN(_27119_));
 DFF_X1 _60536_ (.D(_04942_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [148]),
    .QN(_27120_));
 DFF_X1 _60537_ (.D(_04943_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [149]),
    .QN(_27121_));
 DFF_X1 _60538_ (.D(_04945_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [150]),
    .QN(_27122_));
 DFF_X1 _60539_ (.D(_04946_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [151]),
    .QN(_27123_));
 DFF_X1 _60540_ (.D(_04947_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [152]),
    .QN(_27124_));
 DFF_X1 _60541_ (.D(_04948_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [153]),
    .QN(_27125_));
 DFF_X1 _60542_ (.D(_04949_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [154]),
    .QN(_27126_));
 DFF_X1 _60543_ (.D(_04950_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [155]),
    .QN(_27127_));
 DFF_X1 _60544_ (.D(_04951_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [156]),
    .QN(_27128_));
 DFF_X1 _60545_ (.D(_04952_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [157]),
    .QN(_27129_));
 DFF_X1 _60546_ (.D(_04953_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [158]),
    .QN(_27130_));
 DFF_X1 _60547_ (.D(_04954_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [159]),
    .QN(_27131_));
 DFF_X1 _60548_ (.D(_04956_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [160]),
    .QN(_27132_));
 DFF_X1 _60549_ (.D(_04957_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [161]),
    .QN(_27133_));
 DFF_X1 _60550_ (.D(_04958_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [162]),
    .QN(_27134_));
 DFF_X1 _60551_ (.D(_04959_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [163]),
    .QN(_27135_));
 DFF_X1 _60552_ (.D(_04960_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [164]),
    .QN(_27136_));
 DFF_X1 _60553_ (.D(_04961_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [165]),
    .QN(_27137_));
 DFF_X1 _60554_ (.D(_04962_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [166]),
    .QN(_27138_));
 DFF_X1 _60555_ (.D(_04963_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [167]),
    .QN(_27139_));
 DFF_X1 _60556_ (.D(_04964_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [168]),
    .QN(_27140_));
 DFF_X1 _60557_ (.D(_04965_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [169]),
    .QN(_27141_));
 DFF_X1 _60558_ (.D(_04967_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [170]),
    .QN(_27142_));
 DFF_X1 _60559_ (.D(_04968_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [171]),
    .QN(_27143_));
 DFF_X1 _60560_ (.D(_04969_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [172]),
    .QN(_27144_));
 DFF_X1 _60561_ (.D(_04970_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [173]),
    .QN(_27145_));
 DFF_X1 _60562_ (.D(_04971_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [174]),
    .QN(_27146_));
 DFF_X1 _60563_ (.D(_04972_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [175]),
    .QN(_27147_));
 DFF_X1 _60564_ (.D(_04973_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [176]),
    .QN(_27148_));
 DFF_X1 _60565_ (.D(_04974_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [177]),
    .QN(_27149_));
 DFF_X1 _60566_ (.D(_04975_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [178]),
    .QN(_27150_));
 DFF_X1 _60567_ (.D(_04976_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [179]),
    .QN(_27151_));
 DFF_X1 _60568_ (.D(_04978_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [180]),
    .QN(_27152_));
 DFF_X1 _60569_ (.D(_04979_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [181]),
    .QN(_27153_));
 DFF_X1 _60570_ (.D(_04980_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [182]),
    .QN(_27154_));
 DFF_X1 _60571_ (.D(_04981_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [183]),
    .QN(_27155_));
 DFF_X1 _60572_ (.D(_04982_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [184]),
    .QN(_27156_));
 DFF_X1 _60573_ (.D(_04983_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [185]),
    .QN(_27157_));
 DFF_X1 _60574_ (.D(_04984_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [186]),
    .QN(_27158_));
 DFF_X1 _60575_ (.D(_04985_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [187]),
    .QN(_27159_));
 DFF_X1 _60576_ (.D(_04986_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [188]),
    .QN(_27160_));
 DFF_X1 _60577_ (.D(_04987_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [189]),
    .QN(_27161_));
 DFF_X1 _60578_ (.D(_04989_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [190]),
    .QN(_27162_));
 DFF_X1 _60579_ (.D(_04990_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [191]),
    .QN(_27163_));
 DFF_X1 _60580_ (.D(_04991_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [192]),
    .QN(_27164_));
 DFF_X1 _60581_ (.D(_04992_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [193]),
    .QN(_27165_));
 DFF_X1 _60582_ (.D(_04993_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [194]),
    .QN(_27166_));
 DFF_X1 _60583_ (.D(_04994_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [195]),
    .QN(_27167_));
 DFF_X1 _60584_ (.D(_04995_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [196]),
    .QN(_27168_));
 DFF_X1 _60585_ (.D(_04996_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [197]),
    .QN(_27169_));
 DFF_X1 _60586_ (.D(_04997_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [198]),
    .QN(_27170_));
 DFF_X1 _60587_ (.D(_04998_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [199]),
    .QN(_27171_));
 DFF_X1 _60588_ (.D(_05001_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [200]),
    .QN(_27172_));
 DFF_X1 _60589_ (.D(_05002_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [201]),
    .QN(_27173_));
 DFF_X1 _60590_ (.D(_05003_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [202]),
    .QN(_27174_));
 DFF_X1 _60591_ (.D(_05004_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [203]),
    .QN(_27175_));
 DFF_X1 _60592_ (.D(_05005_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [204]),
    .QN(_27176_));
 DFF_X1 _60593_ (.D(_05006_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [205]),
    .QN(_27177_));
 DFF_X1 _60594_ (.D(_05007_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [206]),
    .QN(_27178_));
 DFF_X1 _60595_ (.D(_05008_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [207]),
    .QN(_27179_));
 DFF_X1 _60596_ (.D(_05009_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [208]),
    .QN(_27180_));
 DFF_X1 _60597_ (.D(_05010_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [209]),
    .QN(_27181_));
 DFF_X1 _60598_ (.D(_05012_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [210]),
    .QN(_27182_));
 DFF_X1 _60599_ (.D(_05013_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [211]),
    .QN(_27183_));
 DFF_X1 _60600_ (.D(_05014_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [212]),
    .QN(_27184_));
 DFF_X1 _60601_ (.D(_05015_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [213]),
    .QN(_27185_));
 DFF_X1 _60602_ (.D(_05016_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [214]),
    .QN(_27186_));
 DFF_X1 _60603_ (.D(_05017_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [215]),
    .QN(_27187_));
 DFF_X1 _60604_ (.D(_05018_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [216]),
    .QN(_27188_));
 DFF_X1 _60605_ (.D(_05019_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [217]),
    .QN(_27189_));
 DFF_X1 _60606_ (.D(_05020_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [218]),
    .QN(_27190_));
 DFF_X1 _60607_ (.D(_05021_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [219]),
    .QN(_27191_));
 DFF_X1 _60608_ (.D(_05023_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [220]),
    .QN(_27192_));
 DFF_X1 _60609_ (.D(_05024_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [221]),
    .QN(_27193_));
 DFF_X1 _60610_ (.D(_05025_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [222]),
    .QN(_27194_));
 DFF_X1 _60611_ (.D(_05026_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [223]),
    .QN(_27195_));
 DFF_X1 _60612_ (.D(_05027_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [224]),
    .QN(_27196_));
 DFF_X1 _60613_ (.D(_05028_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [225]),
    .QN(_27197_));
 DFF_X1 _60614_ (.D(_05029_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [226]),
    .QN(_27198_));
 DFF_X1 _60615_ (.D(_05030_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [227]),
    .QN(_27199_));
 DFF_X1 _60616_ (.D(_05031_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [228]),
    .QN(_27200_));
 DFF_X1 _60617_ (.D(_05032_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [229]),
    .QN(_27201_));
 DFF_X1 _60618_ (.D(_05034_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [230]),
    .QN(_27202_));
 DFF_X1 _60619_ (.D(_05035_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [231]),
    .QN(_27203_));
 DFF_X1 _60620_ (.D(_05036_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [232]),
    .QN(_27204_));
 DFF_X1 _60621_ (.D(_05037_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [233]),
    .QN(_27205_));
 DFF_X1 _60622_ (.D(_05038_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [234]),
    .QN(_27206_));
 DFF_X1 _60623_ (.D(_05039_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [235]),
    .QN(_27207_));
 DFF_X1 _60624_ (.D(_05040_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [236]),
    .QN(_27208_));
 DFF_X1 _60625_ (.D(_05041_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [237]),
    .QN(_27209_));
 DFF_X1 _60626_ (.D(_05042_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [238]),
    .QN(_27210_));
 DFF_X1 _60627_ (.D(_05043_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [239]),
    .QN(_27211_));
 DFF_X1 _60628_ (.D(_05045_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [240]),
    .QN(_27212_));
 DFF_X1 _60629_ (.D(_05046_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [241]),
    .QN(_27213_));
 DFF_X1 _60630_ (.D(_05047_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [242]),
    .QN(_27214_));
 DFF_X1 _60631_ (.D(_05048_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [243]),
    .QN(_27215_));
 DFF_X1 _60632_ (.D(_05049_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [244]),
    .QN(_27216_));
 DFF_X1 _60633_ (.D(_05050_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [245]),
    .QN(_27217_));
 DFF_X1 _60634_ (.D(_05051_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [246]),
    .QN(_27218_));
 DFF_X1 _60635_ (.D(_05052_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [247]),
    .QN(_27219_));
 DFF_X1 _60636_ (.D(_05053_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [248]),
    .QN(_27220_));
 DFF_X1 _60637_ (.D(_05054_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [249]),
    .QN(_27221_));
 DFF_X1 _60638_ (.D(_05056_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [250]),
    .QN(_27222_));
 DFF_X1 _60639_ (.D(_05057_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [251]),
    .QN(_27223_));
 DFF_X1 _60640_ (.D(_05058_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [252]),
    .QN(_27224_));
 DFF_X1 _60641_ (.D(_05059_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [253]),
    .QN(_27225_));
 DFF_X1 _60642_ (.D(_05060_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [254]),
    .QN(_27226_));
 DFF_X1 _60643_ (.D(_05061_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [255]),
    .QN(_27227_));
 DFF_X1 _60644_ (.D(_05062_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [256]),
    .QN(_27228_));
 DFF_X1 _60645_ (.D(_05063_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [257]),
    .QN(_27229_));
 DFF_X1 _60646_ (.D(_05064_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [258]),
    .QN(_27230_));
 DFF_X1 _60647_ (.D(_05065_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [259]),
    .QN(_27231_));
 DFF_X1 _60648_ (.D(_05067_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [260]),
    .QN(_27232_));
 DFF_X1 _60649_ (.D(_05068_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [261]),
    .QN(_27233_));
 DFF_X1 _60650_ (.D(_05069_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [262]),
    .QN(_27234_));
 DFF_X1 _60651_ (.D(_05070_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [263]),
    .QN(_27235_));
 DFF_X1 _60652_ (.D(_05071_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [264]),
    .QN(_27236_));
 DFF_X1 _60653_ (.D(_05072_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [265]),
    .QN(_27237_));
 DFF_X1 _60654_ (.D(_05073_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [266]),
    .QN(_27238_));
 DFF_X1 _60655_ (.D(_05074_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [267]),
    .QN(_27239_));
 DFF_X1 _60656_ (.D(_05075_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [268]),
    .QN(_27240_));
 DFF_X1 _60657_ (.D(_05076_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [269]),
    .QN(_27241_));
 DFF_X1 _60658_ (.D(_05078_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [270]),
    .QN(_27242_));
 DFF_X1 _60659_ (.D(_05079_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [271]),
    .QN(_27243_));
 DFF_X1 _60660_ (.D(_05080_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [272]),
    .QN(_27244_));
 DFF_X1 _60661_ (.D(_05081_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [273]),
    .QN(_27245_));
 DFF_X1 _60662_ (.D(_05082_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [274]),
    .QN(_27246_));
 DFF_X1 _60663_ (.D(_05083_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [275]),
    .QN(_27247_));
 DFF_X1 _60664_ (.D(_05084_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [276]),
    .QN(_27248_));
 DFF_X1 _60665_ (.D(_05085_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [277]),
    .QN(_27249_));
 DFF_X1 _60666_ (.D(_05086_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [278]),
    .QN(_27250_));
 DFF_X1 _60667_ (.D(_05087_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [279]),
    .QN(_27251_));
 DFF_X1 _60668_ (.D(_05089_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [280]),
    .QN(_27252_));
 DFF_X1 _60669_ (.D(_05090_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [281]),
    .QN(_27253_));
 DFF_X1 _60670_ (.D(_05091_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [282]),
    .QN(_27254_));
 DFF_X1 _60671_ (.D(_05092_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [283]),
    .QN(_27255_));
 DFF_X1 _60672_ (.D(_05093_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [284]),
    .QN(_27256_));
 DFF_X1 _60673_ (.D(_05094_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [285]),
    .QN(_27257_));
 DFF_X1 _60674_ (.D(_05095_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [286]),
    .QN(_27258_));
 DFF_X1 _60675_ (.D(_05096_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [287]),
    .QN(_27259_));
 DFF_X1 _60676_ (.D(_05097_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [288]),
    .QN(_27260_));
 DFF_X1 _60677_ (.D(_05098_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [289]),
    .QN(_27261_));
 DFF_X1 _60678_ (.D(_05100_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [290]),
    .QN(_27262_));
 DFF_X1 _60679_ (.D(_05101_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [291]),
    .QN(_27263_));
 DFF_X1 _60680_ (.D(_05102_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [292]),
    .QN(_27264_));
 DFF_X1 _60681_ (.D(_05103_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [293]),
    .QN(_27265_));
 DFF_X1 _60682_ (.D(_05104_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [294]),
    .QN(_27266_));
 DFF_X1 _60683_ (.D(_05105_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [295]),
    .QN(_27267_));
 DFF_X1 _60684_ (.D(_05106_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [296]),
    .QN(_27268_));
 DFF_X1 _60685_ (.D(_05107_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [297]),
    .QN(_27269_));
 DFF_X1 _60686_ (.D(_05108_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [298]),
    .QN(_27270_));
 DFF_X1 _60687_ (.D(_05109_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [299]),
    .QN(_27271_));
 DFF_X1 _60688_ (.D(_05112_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [300]),
    .QN(_27272_));
 DFF_X1 _60689_ (.D(_05113_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [301]),
    .QN(_27273_));
 DFF_X1 _60690_ (.D(_05114_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [302]),
    .QN(_27274_));
 DFF_X1 _60691_ (.D(_05115_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [303]),
    .QN(_27275_));
 DFF_X1 _60692_ (.D(_05116_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [304]),
    .QN(_27276_));
 DFF_X1 _60693_ (.D(_05117_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [305]),
    .QN(_27277_));
 DFF_X1 _60694_ (.D(_05118_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [306]),
    .QN(_27278_));
 DFF_X1 _60695_ (.D(_05119_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [307]),
    .QN(_27279_));
 DFF_X1 _60696_ (.D(_05120_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [308]),
    .QN(_27280_));
 DFF_X1 _60697_ (.D(_05121_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [309]),
    .QN(_27281_));
 DFF_X1 _60698_ (.D(_05123_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [310]),
    .QN(_27282_));
 DFF_X1 _60699_ (.D(_05124_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [311]),
    .QN(_27283_));
 DFF_X1 _60700_ (.D(_05125_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [312]),
    .QN(_27284_));
 DFF_X1 _60701_ (.D(_05126_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [313]),
    .QN(_27285_));
 DFF_X1 _60702_ (.D(_05127_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [314]),
    .QN(_27286_));
 DFF_X1 _60703_ (.D(_05128_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [315]),
    .QN(_27287_));
 DFF_X1 _60704_ (.D(_05129_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [316]),
    .QN(_27288_));
 DFF_X1 _60705_ (.D(_05130_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [317]),
    .QN(_27289_));
 DFF_X1 _60706_ (.D(_05131_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [318]),
    .QN(_27290_));
 DFF_X1 _60707_ (.D(_05132_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [319]),
    .QN(_27291_));
 DFF_X1 _60708_ (.D(_05134_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [320]),
    .QN(_27292_));
 DFF_X1 _60709_ (.D(_05135_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [321]),
    .QN(_27293_));
 DFF_X1 _60710_ (.D(_05136_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [322]),
    .QN(_27294_));
 DFF_X1 _60711_ (.D(_05137_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [323]),
    .QN(_27295_));
 DFF_X1 _60712_ (.D(_05138_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [324]),
    .QN(_27296_));
 DFF_X1 _60713_ (.D(_05139_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [325]),
    .QN(_27297_));
 DFF_X1 _60714_ (.D(_05140_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [326]),
    .QN(_27298_));
 DFF_X1 _60715_ (.D(_05141_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [327]),
    .QN(_27299_));
 DFF_X1 _60716_ (.D(_05142_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [328]),
    .QN(_27300_));
 DFF_X1 _60717_ (.D(_05143_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [329]),
    .QN(_27301_));
 DFF_X1 _60718_ (.D(_05145_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [330]),
    .QN(_27302_));
 DFF_X1 _60719_ (.D(_05146_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [331]),
    .QN(_27303_));
 DFF_X1 _60720_ (.D(_05147_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [332]),
    .QN(_27304_));
 DFF_X1 _60721_ (.D(_05148_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [333]),
    .QN(_27305_));
 DFF_X1 _60722_ (.D(_05149_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [334]),
    .QN(_27306_));
 DFF_X1 _60723_ (.D(_05150_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [335]),
    .QN(_27307_));
 DFF_X1 _60724_ (.D(_05151_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [336]),
    .QN(_27308_));
 DFF_X1 _60725_ (.D(_05152_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [337]),
    .QN(_27309_));
 DFF_X1 _60726_ (.D(_05153_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [338]),
    .QN(_27310_));
 DFF_X1 _60727_ (.D(_05154_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [339]),
    .QN(_27311_));
 DFF_X1 _60728_ (.D(_05156_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [340]),
    .QN(_27312_));
 DFF_X1 _60729_ (.D(_05157_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [341]),
    .QN(_27313_));
 DFF_X1 _60730_ (.D(_05158_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [342]),
    .QN(_27314_));
 DFF_X1 _60731_ (.D(_05159_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [343]),
    .QN(_27315_));
 DFF_X1 _60732_ (.D(_05160_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [344]),
    .QN(_27316_));
 DFF_X1 _60733_ (.D(_05161_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [345]),
    .QN(_27317_));
 DFF_X1 _60734_ (.D(_05162_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [346]),
    .QN(_27318_));
 DFF_X1 _60735_ (.D(_05163_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [347]),
    .QN(_27319_));
 DFF_X1 _60736_ (.D(_05164_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [348]),
    .QN(_27320_));
 DFF_X1 _60737_ (.D(_05165_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [349]),
    .QN(_27321_));
 DFF_X1 _60738_ (.D(_05167_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [350]),
    .QN(_27322_));
 DFF_X1 _60739_ (.D(_05168_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [351]),
    .QN(_27323_));
 DFF_X1 _60740_ (.D(_05169_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [352]),
    .QN(_27324_));
 DFF_X1 _60741_ (.D(_05170_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [353]),
    .QN(_27325_));
 DFF_X1 _60742_ (.D(_05171_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [354]),
    .QN(_27326_));
 DFF_X1 _60743_ (.D(_05172_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [355]),
    .QN(_27327_));
 DFF_X1 _60744_ (.D(_05173_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [356]),
    .QN(_27328_));
 DFF_X1 _60745_ (.D(_05174_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [357]),
    .QN(_27329_));
 DFF_X1 _60746_ (.D(_05175_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [358]),
    .QN(_27330_));
 DFF_X1 _60747_ (.D(_05176_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [359]),
    .QN(_27331_));
 DFF_X1 _60748_ (.D(_05178_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [360]),
    .QN(_27332_));
 DFF_X1 _60749_ (.D(_05179_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [361]),
    .QN(_27333_));
 DFF_X1 _60750_ (.D(_05180_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [362]),
    .QN(_27334_));
 DFF_X1 _60751_ (.D(_05181_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [363]),
    .QN(_27335_));
 DFF_X1 _60752_ (.D(_05182_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [364]),
    .QN(_27336_));
 DFF_X1 _60753_ (.D(_05183_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [365]),
    .QN(_27337_));
 DFF_X1 _60754_ (.D(_05184_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [366]),
    .QN(_27338_));
 DFF_X1 _60755_ (.D(_05185_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [367]),
    .QN(_27339_));
 DFF_X1 _60756_ (.D(_05186_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [368]),
    .QN(_27340_));
 DFF_X1 _60757_ (.D(_05187_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [369]),
    .QN(_27341_));
 DFF_X1 _60758_ (.D(_05189_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [370]),
    .QN(_27342_));
 DFF_X1 _60759_ (.D(_05190_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [371]),
    .QN(_27343_));
 DFF_X1 _60760_ (.D(_05191_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [372]),
    .QN(_27344_));
 DFF_X1 _60761_ (.D(_05192_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [373]),
    .QN(_27345_));
 DFF_X1 _60762_ (.D(_05193_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [374]),
    .QN(_27346_));
 DFF_X1 _60763_ (.D(_05194_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [375]),
    .QN(_27347_));
 DFF_X1 _60764_ (.D(_05195_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [376]),
    .QN(_27348_));
 DFF_X1 _60765_ (.D(_05196_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [377]),
    .QN(_27349_));
 DFF_X1 _60766_ (.D(_05197_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [378]),
    .QN(_27350_));
 DFF_X1 _60767_ (.D(_05198_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [379]),
    .QN(_27351_));
 DFF_X1 _60768_ (.D(_05200_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [380]),
    .QN(_27352_));
 DFF_X1 _60769_ (.D(_05201_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [381]),
    .QN(_27353_));
 DFF_X1 _60770_ (.D(_05202_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [382]),
    .QN(_27354_));
 DFF_X1 _60771_ (.D(_05203_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [383]),
    .QN(_27355_));
 DFF_X1 _60772_ (.D(_05204_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [384]),
    .QN(_27356_));
 DFF_X1 _60773_ (.D(_05205_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [385]),
    .QN(_27357_));
 DFF_X1 _60774_ (.D(_05206_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [386]),
    .QN(_27358_));
 DFF_X1 _60775_ (.D(_05207_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [387]),
    .QN(_27359_));
 DFF_X1 _60776_ (.D(_05208_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [388]),
    .QN(_27360_));
 DFF_X1 _60777_ (.D(_05209_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [389]),
    .QN(_27361_));
 DFF_X1 _60778_ (.D(_05211_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [390]),
    .QN(_27362_));
 DFF_X1 _60779_ (.D(_05212_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [391]),
    .QN(_27363_));
 DFF_X1 _60780_ (.D(_05213_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [392]),
    .QN(_27364_));
 DFF_X1 _60781_ (.D(_05214_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [393]),
    .QN(_27365_));
 DFF_X1 _60782_ (.D(_05215_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [394]),
    .QN(_27366_));
 DFF_X1 _60783_ (.D(_05216_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [395]),
    .QN(_27367_));
 DFF_X1 _60784_ (.D(_05217_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [396]),
    .QN(_27368_));
 DFF_X1 _60785_ (.D(_05218_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [397]),
    .QN(_27369_));
 DFF_X1 _60786_ (.D(_05219_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [398]),
    .QN(_27370_));
 DFF_X1 _60787_ (.D(_05220_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [399]),
    .QN(_27371_));
 DFF_X1 _60788_ (.D(_05223_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [400]),
    .QN(_27372_));
 DFF_X1 _60789_ (.D(_05224_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [401]),
    .QN(_27373_));
 DFF_X1 _60790_ (.D(_05225_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [402]),
    .QN(_27374_));
 DFF_X1 _60791_ (.D(_05226_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [403]),
    .QN(_27375_));
 DFF_X1 _60792_ (.D(_05227_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [404]),
    .QN(_27376_));
 DFF_X1 _60793_ (.D(_05228_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [405]),
    .QN(_27377_));
 DFF_X1 _60794_ (.D(_05229_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [406]),
    .QN(_27378_));
 DFF_X1 _60795_ (.D(_05230_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [407]),
    .QN(_27379_));
 DFF_X1 _60796_ (.D(_05231_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [408]),
    .QN(_27380_));
 DFF_X1 _60797_ (.D(_05232_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [409]),
    .QN(_27381_));
 DFF_X1 _60798_ (.D(_05234_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [410]),
    .QN(_27382_));
 DFF_X1 _60799_ (.D(_05235_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [411]),
    .QN(_27383_));
 DFF_X1 _60800_ (.D(_05236_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [412]),
    .QN(_27384_));
 DFF_X1 _60801_ (.D(_05237_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [413]),
    .QN(_27385_));
 DFF_X1 _60802_ (.D(_05238_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [414]),
    .QN(_27386_));
 DFF_X1 _60803_ (.D(_05239_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [415]),
    .QN(_27387_));
 DFF_X1 _60804_ (.D(_05240_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [416]),
    .QN(_27388_));
 DFF_X1 _60805_ (.D(_05241_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [417]),
    .QN(_27389_));
 DFF_X1 _60806_ (.D(_05242_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [418]),
    .QN(_27390_));
 DFF_X1 _60807_ (.D(_05243_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [419]),
    .QN(_27391_));
 DFF_X1 _60808_ (.D(_05245_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [420]),
    .QN(_27392_));
 DFF_X1 _60809_ (.D(_05246_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [421]),
    .QN(_27393_));
 DFF_X1 _60810_ (.D(_05247_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [422]),
    .QN(_27394_));
 DFF_X1 _60811_ (.D(_05248_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [423]),
    .QN(_27395_));
 DFF_X1 _60812_ (.D(_05249_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [424]),
    .QN(_27396_));
 DFF_X1 _60813_ (.D(_05250_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [425]),
    .QN(_27397_));
 DFF_X1 _60814_ (.D(_05251_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [426]),
    .QN(_27398_));
 DFF_X1 _60815_ (.D(_05252_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [427]),
    .QN(_27399_));
 DFF_X1 _60816_ (.D(_05253_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [428]),
    .QN(_27400_));
 DFF_X1 _60817_ (.D(_05254_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [429]),
    .QN(_27401_));
 DFF_X1 _60818_ (.D(_05256_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [430]),
    .QN(_27402_));
 DFF_X1 _60819_ (.D(_05257_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [431]),
    .QN(_27403_));
 DFF_X1 _60820_ (.D(_05258_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [432]),
    .QN(_27404_));
 DFF_X1 _60821_ (.D(_05259_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [433]),
    .QN(_27405_));
 DFF_X1 _60822_ (.D(_05260_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [434]),
    .QN(_27406_));
 DFF_X1 _60823_ (.D(_05261_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [435]),
    .QN(_27407_));
 DFF_X1 _60824_ (.D(_05262_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [436]),
    .QN(_27408_));
 DFF_X1 _60825_ (.D(_05263_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [437]),
    .QN(_27409_));
 DFF_X1 _60826_ (.D(_05264_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [438]),
    .QN(_27410_));
 DFF_X1 _60827_ (.D(_05265_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [439]),
    .QN(_27411_));
 DFF_X1 _60828_ (.D(_05267_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [440]),
    .QN(_27412_));
 DFF_X1 _60829_ (.D(_05268_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [441]),
    .QN(_27413_));
 DFF_X1 _60830_ (.D(_05269_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [442]),
    .QN(_27414_));
 DFF_X1 _60831_ (.D(_05270_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [443]),
    .QN(_27415_));
 DFF_X1 _60832_ (.D(_05271_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [444]),
    .QN(_27416_));
 DFF_X1 _60833_ (.D(_05272_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [445]),
    .QN(_27417_));
 DFF_X1 _60834_ (.D(_05273_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [446]),
    .QN(_27418_));
 DFF_X1 _60835_ (.D(_05274_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [447]),
    .QN(_27419_));
 DFF_X1 _60836_ (.D(_05275_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [448]),
    .QN(_27420_));
 DFF_X1 _60837_ (.D(_05276_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [449]),
    .QN(_27421_));
 DFF_X1 _60838_ (.D(_05278_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [450]),
    .QN(_27422_));
 DFF_X1 _60839_ (.D(_05279_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [451]),
    .QN(_27423_));
 DFF_X1 _60840_ (.D(_05280_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [452]),
    .QN(_27424_));
 DFF_X1 _60841_ (.D(_05281_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [453]),
    .QN(_27425_));
 DFF_X1 _60842_ (.D(_05282_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [454]),
    .QN(_27426_));
 DFF_X1 _60843_ (.D(_05283_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [455]),
    .QN(_27427_));
 DFF_X1 _60844_ (.D(_05284_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [456]),
    .QN(_27428_));
 DFF_X1 _60845_ (.D(_05285_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [457]),
    .QN(_27429_));
 DFF_X1 _60846_ (.D(_05286_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [458]),
    .QN(_27430_));
 DFF_X1 _60847_ (.D(_05287_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [459]),
    .QN(_27431_));
 DFF_X1 _60848_ (.D(_05289_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [460]),
    .QN(_27432_));
 DFF_X1 _60849_ (.D(_05290_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [461]),
    .QN(_27433_));
 DFF_X1 _60850_ (.D(_05291_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [462]),
    .QN(_27434_));
 DFF_X1 _60851_ (.D(_05292_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [463]),
    .QN(_27435_));
 DFF_X1 _60852_ (.D(_05293_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [464]),
    .QN(_27436_));
 DFF_X1 _60853_ (.D(_05294_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [465]),
    .QN(_27437_));
 DFF_X1 _60854_ (.D(_05295_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [466]),
    .QN(_27438_));
 DFF_X1 _60855_ (.D(_05296_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [467]),
    .QN(_27439_));
 DFF_X1 _60856_ (.D(_05297_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [468]),
    .QN(_27440_));
 DFF_X1 _60857_ (.D(_05298_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [469]),
    .QN(_27441_));
 DFF_X1 _60858_ (.D(_05300_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [470]),
    .QN(_27442_));
 DFF_X1 _60859_ (.D(_05301_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [471]),
    .QN(_27443_));
 DFF_X1 _60860_ (.D(_05302_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [472]),
    .QN(_27444_));
 DFF_X1 _60861_ (.D(_05303_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [473]),
    .QN(_27445_));
 DFF_X1 _60862_ (.D(_05304_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [474]),
    .QN(_27446_));
 DFF_X1 _60863_ (.D(_05305_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [475]),
    .QN(_27447_));
 DFF_X1 _60864_ (.D(_05306_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [476]),
    .QN(_27448_));
 DFF_X1 _60865_ (.D(_05307_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [477]),
    .QN(_27449_));
 DFF_X1 _60866_ (.D(_05308_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [478]),
    .QN(_27450_));
 DFF_X1 _60867_ (.D(_05309_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [479]),
    .QN(_27451_));
 DFF_X1 _60868_ (.D(_05311_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [480]),
    .QN(_27452_));
 DFF_X1 _60869_ (.D(_05312_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [481]),
    .QN(_27453_));
 DFF_X1 _60870_ (.D(_05313_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [482]),
    .QN(_27454_));
 DFF_X1 _60871_ (.D(_05314_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [483]),
    .QN(_27455_));
 DFF_X1 _60872_ (.D(_05315_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [484]),
    .QN(_27456_));
 DFF_X1 _60873_ (.D(_05316_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [485]),
    .QN(_27457_));
 DFF_X1 _60874_ (.D(_05317_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [486]),
    .QN(_27458_));
 DFF_X1 _60875_ (.D(_05318_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [487]),
    .QN(_27459_));
 DFF_X1 _60876_ (.D(_05319_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [488]),
    .QN(_27460_));
 DFF_X1 _60877_ (.D(_05320_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [489]),
    .QN(_27461_));
 DFF_X1 _60878_ (.D(_05322_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [490]),
    .QN(_27462_));
 DFF_X1 _60879_ (.D(_05323_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [491]),
    .QN(_27463_));
 DFF_X1 _60880_ (.D(_05324_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [492]),
    .QN(_27464_));
 DFF_X1 _60881_ (.D(_05325_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [493]),
    .QN(_27465_));
 DFF_X1 _60882_ (.D(_05326_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [494]),
    .QN(_27466_));
 DFF_X1 _60883_ (.D(_05327_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [495]),
    .QN(_27467_));
 DFF_X1 _60884_ (.D(_05328_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [496]),
    .QN(_27468_));
 DFF_X1 _60885_ (.D(_05329_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [497]),
    .QN(_27469_));
 DFF_X1 _60886_ (.D(_05330_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [498]),
    .QN(_27470_));
 DFF_X1 _60887_ (.D(_05331_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [499]),
    .QN(_27471_));
 DFF_X1 _60888_ (.D(_05334_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [500]),
    .QN(_27472_));
 DFF_X1 _60889_ (.D(_05335_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [501]),
    .QN(_27473_));
 DFF_X1 _60890_ (.D(_05336_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [502]),
    .QN(_27474_));
 DFF_X1 _60891_ (.D(_05337_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [503]),
    .QN(_27475_));
 DFF_X1 _60892_ (.D(_05338_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [504]),
    .QN(_27476_));
 DFF_X1 _60893_ (.D(_05339_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [505]),
    .QN(_27477_));
 DFF_X1 _60894_ (.D(_05340_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [506]),
    .QN(_27478_));
 DFF_X1 _60895_ (.D(_05341_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [507]),
    .QN(_27479_));
 DFF_X1 _60896_ (.D(_05342_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [508]),
    .QN(_27480_));
 DFF_X1 _60897_ (.D(_05343_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [509]),
    .QN(_27481_));
 DFF_X1 _60898_ (.D(_05345_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [510]),
    .QN(_27482_));
 DFF_X1 _60899_ (.D(_05346_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.data_r [511]),
    .QN(_27483_));
 DFF_X1 _60900_ (.D(_05403_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.state_r [0]),
    .QN(_00599_));
 DFF_X1 _60901_ (.D(_05404_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.state_r [1]),
    .QN(_00598_));
 DFF_X1 _60902_ (.D(_06588_),
    .CK(clk_i),
    .Q(\icache.lce.lce_req_inst.set_tag_received_r ),
    .QN(_00601_));
 DFF_X1 _60903_ (.D(_06548_),
    .CK(clk_i),
    .Q(\icache.lce.lce_req_inst.cce_data_received_r ),
    .QN(_00603_));
 DFF_X1 _60904_ (.D(_06549_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.miss_addr_i [0]),
    .QN(_00606_));
 DFF_X1 _60905_ (.D(_06560_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.miss_addr_i [1]),
    .QN(_00607_));
 DFF_X1 _60906_ (.D(_06571_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.miss_addr_i [2]),
    .QN(_00608_));
 DFF_X1 _60907_ (.D(_06581_),
    .CK(clk_i),
    .Q(lce_req_o[10]),
    .QN(_27484_));
 DFF_X1 _60908_ (.D(_06582_),
    .CK(clk_i),
    .Q(lce_req_o[11]),
    .QN(_27485_));
 DFF_X1 _60909_ (.D(_06583_),
    .CK(clk_i),
    .Q(lce_req_o[12]),
    .QN(_27486_));
 DFF_X1 _60910_ (.D(_06584_),
    .CK(clk_i),
    .Q(lce_req_o[13]),
    .QN(_27487_));
 DFF_X1 _60911_ (.D(_06585_),
    .CK(clk_i),
    .Q(lce_req_o[14]),
    .QN(_27488_));
 DFF_X1 _60912_ (.D(_06586_),
    .CK(clk_i),
    .Q(lce_req_o[15]),
    .QN(_27489_));
 DFF_X1 _60913_ (.D(_06587_),
    .CK(clk_i),
    .Q(lce_req_o[16]),
    .QN(_27490_));
 DFF_X1 _60914_ (.D(_06550_),
    .CK(clk_i),
    .Q(lce_req_o[17]),
    .QN(_27491_));
 DFF_X1 _60915_ (.D(_06551_),
    .CK(clk_i),
    .Q(lce_req_o[18]),
    .QN(_27492_));
 DFF_X1 _60916_ (.D(_06552_),
    .CK(clk_i),
    .Q(lce_req_o[19]),
    .QN(_27493_));
 DFF_X1 _60917_ (.D(_06553_),
    .CK(clk_i),
    .Q(lce_req_o[20]),
    .QN(_27494_));
 DFF_X1 _60918_ (.D(_06554_),
    .CK(clk_i),
    .Q(lce_req_o[21]),
    .QN(_27495_));
 DFF_X1 _60919_ (.D(_06555_),
    .CK(clk_i),
    .Q(lce_req_o[22]),
    .QN(_27496_));
 DFF_X1 _60920_ (.D(_06556_),
    .CK(clk_i),
    .Q(lce_req_o[23]),
    .QN(_27497_));
 DFF_X1 _60921_ (.D(_06557_),
    .CK(clk_i),
    .Q(lce_req_o[24]),
    .QN(_27498_));
 DFF_X1 _60922_ (.D(_06558_),
    .CK(clk_i),
    .Q(lce_req_o[25]),
    .QN(_27499_));
 DFF_X1 _60923_ (.D(_06559_),
    .CK(clk_i),
    .Q(lce_req_o[26]),
    .QN(_27500_));
 DFF_X1 _60924_ (.D(_06561_),
    .CK(clk_i),
    .Q(lce_req_o[27]),
    .QN(_27501_));
 DFF_X1 _60925_ (.D(_06562_),
    .CK(clk_i),
    .Q(lce_req_o[28]),
    .QN(_27502_));
 DFF_X1 _60926_ (.D(_06563_),
    .CK(clk_i),
    .Q(lce_req_o[29]),
    .QN(_27503_));
 DFF_X1 _60927_ (.D(_06564_),
    .CK(clk_i),
    .Q(lce_req_o[30]),
    .QN(_27504_));
 DFF_X1 _60928_ (.D(_06565_),
    .CK(clk_i),
    .Q(lce_req_o[31]),
    .QN(_27505_));
 DFF_X1 _60929_ (.D(_06566_),
    .CK(clk_i),
    .Q(lce_req_o[32]),
    .QN(_27506_));
 DFF_X1 _60930_ (.D(_06567_),
    .CK(clk_i),
    .Q(lce_req_o[33]),
    .QN(_27507_));
 DFF_X1 _60931_ (.D(_06568_),
    .CK(clk_i),
    .Q(lce_req_o[34]),
    .QN(_27508_));
 DFF_X1 _60932_ (.D(_06569_),
    .CK(clk_i),
    .Q(lce_req_o[35]),
    .QN(_27509_));
 DFF_X1 _60933_ (.D(_06570_),
    .CK(clk_i),
    .Q(lce_req_o[36]),
    .QN(_27510_));
 DFF_X1 _60934_ (.D(_06572_),
    .CK(clk_i),
    .Q(lce_req_o[37]),
    .QN(_27511_));
 DFF_X1 _60935_ (.D(_06573_),
    .CK(clk_i),
    .Q(lce_req_o[38]),
    .QN(_27512_));
 DFF_X1 _60936_ (.D(_06574_),
    .CK(clk_i),
    .Q(lce_req_o[39]),
    .QN(_27513_));
 DFF_X1 _60937_ (.D(_06575_),
    .CK(clk_i),
    .Q(lce_req_o[40]),
    .QN(_27514_));
 DFF_X1 _60938_ (.D(_06576_),
    .CK(clk_i),
    .Q(lce_req_o[41]),
    .QN(_27515_));
 DFF_X1 _60939_ (.D(_06577_),
    .CK(clk_i),
    .Q(lce_req_o[42]),
    .QN(_27516_));
 DFF_X1 _60940_ (.D(_06578_),
    .CK(clk_i),
    .Q(lce_req_o[43]),
    .QN(_27517_));
 DFF_X1 _60941_ (.D(_06579_),
    .CK(clk_i),
    .Q(lce_req_o[44]),
    .QN(_27518_));
 DFF_X1 _60942_ (.D(_06580_),
    .CK(clk_i),
    .Q(lce_req_o[45]),
    .QN(_27519_));
 DFF_X1 _60943_ (.D(_06589_),
    .CK(clk_i),
    .Q(\icache.lce.lce_req_inst.state_r [0]),
    .QN(_00002_));
 DFF_X1 _60944_ (.D(_06590_),
    .CK(clk_i),
    .Q(\icache.lce.lce_req_inst.state_r [1]),
    .QN(_00604_));
 DFF_X1 _60945_ (.D(_06591_),
    .CK(clk_i),
    .Q(\icache.lce.lce_req_inst.state_r [2]),
    .QN(_00605_));
 DFF_X1 _60946_ (.D(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [0]),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.br_tgt_o [0]),
    .QN(_27520_));
 DFF_X1 _60947_ (.D(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [1]),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.br_tgt_o [1]),
    .QN(_27521_));
 DFF_X1 _60948_ (.D(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [2]),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.br_tgt_o [2]),
    .QN(_00082_));
 DFF_X1 _60949_ (.D(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [3]),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.br_tgt_o [3]),
    .QN(_00077_));
 DFF_X1 _60950_ (.D(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [4]),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.br_tgt_o [4]),
    .QN(_27522_));
 DFF_X1 _60951_ (.D(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [5]),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.br_tgt_o [5]),
    .QN(_27523_));
 DFF_X1 _60952_ (.D(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [6]),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.br_tgt_o [6]),
    .QN(_27524_));
 DFF_X1 _60953_ (.D(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [7]),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.br_tgt_o [7]),
    .QN(_27525_));
 DFF_X1 _60954_ (.D(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [8]),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.br_tgt_o [8]),
    .QN(_27526_));
 DFF_X1 _60955_ (.D(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [9]),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.br_tgt_o [9]),
    .QN(_27527_));
 DFF_X1 _60956_ (.D(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [10]),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.br_tgt_o [10]),
    .QN(_27528_));
 DFF_X1 _60957_ (.D(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [11]),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.br_tgt_o [11]),
    .QN(_27529_));
 DFF_X1 _60958_ (.D(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [12]),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.br_tgt_o [12]),
    .QN(_27530_));
 DFF_X1 _60959_ (.D(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [13]),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.br_tgt_o [13]),
    .QN(_27531_));
 DFF_X1 _60960_ (.D(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [14]),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.br_tgt_o [14]),
    .QN(_27532_));
 DFF_X1 _60961_ (.D(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [15]),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.br_tgt_o [15]),
    .QN(_27533_));
 DFF_X1 _60962_ (.D(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [16]),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.br_tgt_o [16]),
    .QN(_27534_));
 DFF_X1 _60963_ (.D(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [17]),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.br_tgt_o [17]),
    .QN(_27535_));
 DFF_X1 _60964_ (.D(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [18]),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.br_tgt_o [18]),
    .QN(_27536_));
 DFF_X1 _60965_ (.D(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [19]),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.br_tgt_o [19]),
    .QN(_27537_));
 DFF_X1 _60966_ (.D(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [20]),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.br_tgt_o [20]),
    .QN(_27538_));
 DFF_X1 _60967_ (.D(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [21]),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.br_tgt_o [21]),
    .QN(_27539_));
 DFF_X1 _60968_ (.D(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [22]),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.br_tgt_o [22]),
    .QN(_27540_));
 DFF_X1 _60969_ (.D(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [23]),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.br_tgt_o [23]),
    .QN(_27541_));
 DFF_X1 _60970_ (.D(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [24]),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.br_tgt_o [24]),
    .QN(_27542_));
 DFF_X1 _60971_ (.D(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [25]),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.br_tgt_o [25]),
    .QN(_27543_));
 DFF_X1 _60972_ (.D(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [26]),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.br_tgt_o [26]),
    .QN(_27544_));
 DFF_X1 _60973_ (.D(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [27]),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.br_tgt_o [27]),
    .QN(_27545_));
 DFF_X1 _60974_ (.D(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [28]),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.br_tgt_o [28]),
    .QN(_27546_));
 DFF_X1 _60975_ (.D(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [29]),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.br_tgt_o [29]),
    .QN(_27547_));
 DFF_X1 _60976_ (.D(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [30]),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.br_tgt_o [30]),
    .QN(_27548_));
 DFF_X1 _60977_ (.D(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [31]),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.br_tgt_o [31]),
    .QN(_27549_));
 DFF_X1 _60978_ (.D(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [32]),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.br_tgt_o [32]),
    .QN(_27550_));
 DFF_X1 _60979_ (.D(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [33]),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.br_tgt_o [33]),
    .QN(_27551_));
 DFF_X1 _60980_ (.D(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [34]),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.br_tgt_o [34]),
    .QN(_27552_));
 DFF_X1 _60981_ (.D(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [35]),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.br_tgt_o [35]),
    .QN(_27553_));
 DFF_X1 _60982_ (.D(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [36]),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.br_tgt_o [36]),
    .QN(_27554_));
 DFF_X1 _60983_ (.D(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [37]),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.br_tgt_o [37]),
    .QN(_27555_));
 DFF_X1 _60984_ (.D(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [38]),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.br_tgt_o [38]),
    .QN(_27556_));
 DFF_X1 _60985_ (.D(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [39]),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.data_o [39]),
    .QN(_27557_));
 DFF_X1 _60986_ (.D(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [40]),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.data_o [40]),
    .QN(_27558_));
 DFF_X1 _60987_ (.D(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [41]),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.data_o [41]),
    .QN(_27559_));
 DFF_X1 _60988_ (.D(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [42]),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.data_o [42]),
    .QN(_27560_));
 DFF_X1 _60989_ (.D(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [43]),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.data_o [43]),
    .QN(_27561_));
 DFF_X1 _60990_ (.D(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [44]),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.data_o [44]),
    .QN(_27562_));
 DFF_X1 _60991_ (.D(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [45]),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.data_o [45]),
    .QN(_27563_));
 DFF_X1 _60992_ (.D(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [46]),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.data_o [46]),
    .QN(_27564_));
 DFF_X1 _60993_ (.D(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [47]),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.data_o [47]),
    .QN(_27565_));
 DFF_X1 _60994_ (.D(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_data_lo [48]),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.data_o [48]),
    .QN(_27566_));
 DFF_X1 _60995_ (.D(_06593_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [0]),
    .QN(_27567_));
 DFF_X1 _60996_ (.D(_06785_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [6]),
    .QN(_27568_));
 DFF_X1 _60997_ (.D(_06794_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [7]),
    .QN(_27569_));
 DFF_X1 _60998_ (.D(_06805_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [8]),
    .QN(_27570_));
 DFF_X1 _60999_ (.D(_06816_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [9]),
    .QN(_27571_));
 DFF_X1 _61000_ (.D(_06599_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [10]),
    .QN(_27572_));
 DFF_X1 _61001_ (.D(_06610_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [11]),
    .QN(_27573_));
 DFF_X1 _61002_ (.D(_06621_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [12]),
    .QN(_27574_));
 DFF_X1 _61003_ (.D(_06627_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [13]),
    .QN(_27575_));
 DFF_X1 _61004_ (.D(_06638_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [14]),
    .QN(_27576_));
 DFF_X1 _61005_ (.D(_06649_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [15]),
    .QN(_27577_));
 DFF_X1 _61006_ (.D(_06656_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [16]),
    .QN(_27578_));
 DFF_X1 _61007_ (.D(_06666_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [17]),
    .QN(_27579_));
 DFF_X1 _61008_ (.D(_06677_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [18]),
    .QN(_27580_));
 DFF_X1 _61009_ (.D(_06687_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [19]),
    .QN(_27581_));
 DFF_X1 _61010_ (.D(_06694_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [20]),
    .QN(_27582_));
 DFF_X1 _61011_ (.D(_06705_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [21]),
    .QN(_27583_));
 DFF_X1 _61012_ (.D(_06716_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [22]),
    .QN(_27584_));
 DFF_X1 _61013_ (.D(_06722_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [23]),
    .QN(_27585_));
 DFF_X1 _61014_ (.D(_06733_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [24]),
    .QN(_27586_));
 DFF_X1 _61015_ (.D(_06744_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [25]),
    .QN(_27587_));
 DFF_X1 _61016_ (.D(_06749_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [26]),
    .QN(_27588_));
 DFF_X1 _61017_ (.D(_06750_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [27]),
    .QN(_27589_));
 DFF_X1 _61018_ (.D(_06751_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [28]),
    .QN(_27590_));
 DFF_X1 _61019_ (.D(_06752_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [29]),
    .QN(_27591_));
 DFF_X1 _61020_ (.D(_06753_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [30]),
    .QN(_27592_));
 DFF_X1 _61021_ (.D(_06754_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [31]),
    .QN(_27593_));
 DFF_X1 _61022_ (.D(_06755_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [32]),
    .QN(_27594_));
 DFF_X1 _61023_ (.D(_06756_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [33]),
    .QN(_27595_));
 DFF_X1 _61024_ (.D(_06757_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [39]),
    .QN(_27596_));
 DFF_X1 _61025_ (.D(_06758_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [40]),
    .QN(_27597_));
 DFF_X1 _61026_ (.D(_06759_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [41]),
    .QN(_27598_));
 DFF_X1 _61027_ (.D(_06760_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [42]),
    .QN(_27599_));
 DFF_X1 _61028_ (.D(_06761_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [43]),
    .QN(_27600_));
 DFF_X1 _61029_ (.D(_06762_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [44]),
    .QN(_27601_));
 DFF_X1 _61030_ (.D(_06763_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [45]),
    .QN(_27602_));
 DFF_X1 _61031_ (.D(_06764_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [46]),
    .QN(_27603_));
 DFF_X1 _61032_ (.D(_06765_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [47]),
    .QN(_27604_));
 DFF_X1 _61033_ (.D(_06766_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [48]),
    .QN(_27605_));
 DFF_X1 _61034_ (.D(_06767_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [49]),
    .QN(_27606_));
 DFF_X1 _61035_ (.D(_06768_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [50]),
    .QN(_27607_));
 DFF_X1 _61036_ (.D(_06769_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [51]),
    .QN(_27608_));
 DFF_X1 _61037_ (.D(_06770_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [52]),
    .QN(_27609_));
 DFF_X1 _61038_ (.D(_06771_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [53]),
    .QN(_27610_));
 DFF_X1 _61039_ (.D(_06772_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [54]),
    .QN(_27611_));
 DFF_X1 _61040_ (.D(_06773_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [55]),
    .QN(_27612_));
 DFF_X1 _61041_ (.D(_06774_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [56]),
    .QN(_27613_));
 DFF_X1 _61042_ (.D(_06775_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [57]),
    .QN(_27614_));
 DFF_X1 _61043_ (.D(_06776_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [58]),
    .QN(_27615_));
 DFF_X1 _61044_ (.D(_06777_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [59]),
    .QN(_27616_));
 DFF_X1 _61045_ (.D(_06778_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [60]),
    .QN(_27617_));
 DFF_X1 _61046_ (.D(_06779_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [61]),
    .QN(_27618_));
 DFF_X1 _61047_ (.D(_06780_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [62]),
    .QN(_27619_));
 DFF_X1 _61048_ (.D(_06781_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [63]),
    .QN(_27620_));
 DFF_X1 _61049_ (.D(_06782_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [64]),
    .QN(_27621_));
 DFF_X1 _61050_ (.D(_06783_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [65]),
    .QN(_27622_));
 DFF_X1 _61051_ (.D(_06784_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [66]),
    .QN(_27623_));
 DFF_X1 _61052_ (.D(_06786_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [72]),
    .QN(_27624_));
 DFF_X1 _61053_ (.D(_06787_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [73]),
    .QN(_27625_));
 DFF_X1 _61054_ (.D(_06788_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [74]),
    .QN(_27626_));
 DFF_X1 _61055_ (.D(_06789_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [75]),
    .QN(_27627_));
 DFF_X1 _61056_ (.D(_06790_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [76]),
    .QN(_27628_));
 DFF_X1 _61057_ (.D(_06791_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [77]),
    .QN(_27629_));
 DFF_X1 _61058_ (.D(_06792_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [78]),
    .QN(_27630_));
 DFF_X1 _61059_ (.D(_06793_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [79]),
    .QN(_27631_));
 DFF_X1 _61060_ (.D(_06795_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [80]),
    .QN(_27632_));
 DFF_X1 _61061_ (.D(_06796_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [81]),
    .QN(_27633_));
 DFF_X1 _61062_ (.D(_06797_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [82]),
    .QN(_27634_));
 DFF_X1 _61063_ (.D(_06798_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [83]),
    .QN(_27635_));
 DFF_X1 _61064_ (.D(_06799_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [84]),
    .QN(_27636_));
 DFF_X1 _61065_ (.D(_06800_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [85]),
    .QN(_27637_));
 DFF_X1 _61066_ (.D(_06801_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [86]),
    .QN(_27638_));
 DFF_X1 _61067_ (.D(_06802_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [87]),
    .QN(_27639_));
 DFF_X1 _61068_ (.D(_06803_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [88]),
    .QN(_27640_));
 DFF_X1 _61069_ (.D(_06804_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [89]),
    .QN(_27641_));
 DFF_X1 _61070_ (.D(_06806_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [90]),
    .QN(_27642_));
 DFF_X1 _61071_ (.D(_06807_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [91]),
    .QN(_27643_));
 DFF_X1 _61072_ (.D(_06808_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [92]),
    .QN(_27644_));
 DFF_X1 _61073_ (.D(_06809_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [93]),
    .QN(_27645_));
 DFF_X1 _61074_ (.D(_06810_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [94]),
    .QN(_27646_));
 DFF_X1 _61075_ (.D(_06811_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [95]),
    .QN(_27647_));
 DFF_X1 _61076_ (.D(_06812_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [96]),
    .QN(_27648_));
 DFF_X1 _61077_ (.D(_06813_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [97]),
    .QN(_27649_));
 DFF_X1 _61078_ (.D(_06814_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [98]),
    .QN(_27650_));
 DFF_X1 _61079_ (.D(_06815_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [99]),
    .QN(_27651_));
 DFF_X1 _61080_ (.D(_06594_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [105]),
    .QN(_27652_));
 DFF_X1 _61081_ (.D(_06595_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [106]),
    .QN(_27653_));
 DFF_X1 _61082_ (.D(_06596_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [107]),
    .QN(_27654_));
 DFF_X1 _61083_ (.D(_06597_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [108]),
    .QN(_27655_));
 DFF_X1 _61084_ (.D(_06598_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [109]),
    .QN(_27656_));
 DFF_X1 _61085_ (.D(_06600_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [110]),
    .QN(_27657_));
 DFF_X1 _61086_ (.D(_06601_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [111]),
    .QN(_27658_));
 DFF_X1 _61087_ (.D(_06602_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [112]),
    .QN(_27659_));
 DFF_X1 _61088_ (.D(_06603_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [113]),
    .QN(_27660_));
 DFF_X1 _61089_ (.D(_06604_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [114]),
    .QN(_27661_));
 DFF_X1 _61090_ (.D(_06605_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [115]),
    .QN(_27662_));
 DFF_X1 _61091_ (.D(_06606_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [116]),
    .QN(_27663_));
 DFF_X1 _61092_ (.D(_06607_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [117]),
    .QN(_27664_));
 DFF_X1 _61093_ (.D(_06608_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [118]),
    .QN(_27665_));
 DFF_X1 _61094_ (.D(_06609_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [119]),
    .QN(_27666_));
 DFF_X1 _61095_ (.D(_06611_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [120]),
    .QN(_27667_));
 DFF_X1 _61096_ (.D(_06612_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [121]),
    .QN(_27668_));
 DFF_X1 _61097_ (.D(_06613_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [122]),
    .QN(_27669_));
 DFF_X1 _61098_ (.D(_06614_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [123]),
    .QN(_27670_));
 DFF_X1 _61099_ (.D(_06615_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [124]),
    .QN(_27671_));
 DFF_X1 _61100_ (.D(_06616_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [125]),
    .QN(_27672_));
 DFF_X1 _61101_ (.D(_06617_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [126]),
    .QN(_27673_));
 DFF_X1 _61102_ (.D(_06618_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [127]),
    .QN(_27674_));
 DFF_X1 _61103_ (.D(_06619_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [128]),
    .QN(_27675_));
 DFF_X1 _61104_ (.D(_06620_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [129]),
    .QN(_27676_));
 DFF_X1 _61105_ (.D(_06622_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [130]),
    .QN(_27677_));
 DFF_X1 _61106_ (.D(_06623_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [131]),
    .QN(_27678_));
 DFF_X1 _61107_ (.D(_06624_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [132]),
    .QN(_27679_));
 DFF_X1 _61108_ (.D(_06625_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [138]),
    .QN(_27680_));
 DFF_X1 _61109_ (.D(_06626_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [139]),
    .QN(_27681_));
 DFF_X1 _61110_ (.D(_06628_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [140]),
    .QN(_27682_));
 DFF_X1 _61111_ (.D(_06629_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [141]),
    .QN(_27683_));
 DFF_X1 _61112_ (.D(_06630_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [142]),
    .QN(_27684_));
 DFF_X1 _61113_ (.D(_06631_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [143]),
    .QN(_27685_));
 DFF_X1 _61114_ (.D(_06632_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [144]),
    .QN(_27686_));
 DFF_X1 _61115_ (.D(_06633_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [145]),
    .QN(_27687_));
 DFF_X1 _61116_ (.D(_06634_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [146]),
    .QN(_27688_));
 DFF_X1 _61117_ (.D(_06635_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [147]),
    .QN(_27689_));
 DFF_X1 _61118_ (.D(_06636_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [148]),
    .QN(_27690_));
 DFF_X1 _61119_ (.D(_06637_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [149]),
    .QN(_27691_));
 DFF_X1 _61120_ (.D(_06639_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [150]),
    .QN(_27692_));
 DFF_X1 _61121_ (.D(_06640_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [151]),
    .QN(_27693_));
 DFF_X1 _61122_ (.D(_06641_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [152]),
    .QN(_27694_));
 DFF_X1 _61123_ (.D(_06642_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [153]),
    .QN(_27695_));
 DFF_X1 _61124_ (.D(_06643_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [154]),
    .QN(_27696_));
 DFF_X1 _61125_ (.D(_06644_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [155]),
    .QN(_27697_));
 DFF_X1 _61126_ (.D(_06645_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [156]),
    .QN(_27698_));
 DFF_X1 _61127_ (.D(_06646_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [157]),
    .QN(_27699_));
 DFF_X1 _61128_ (.D(_06647_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [158]),
    .QN(_27700_));
 DFF_X1 _61129_ (.D(_06648_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [159]),
    .QN(_27701_));
 DFF_X1 _61130_ (.D(_06650_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [160]),
    .QN(_27702_));
 DFF_X1 _61131_ (.D(_06651_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [161]),
    .QN(_27703_));
 DFF_X1 _61132_ (.D(_06652_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [162]),
    .QN(_27704_));
 DFF_X1 _61133_ (.D(_06653_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [163]),
    .QN(_27705_));
 DFF_X1 _61134_ (.D(_06654_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [164]),
    .QN(_27706_));
 DFF_X1 _61135_ (.D(_06655_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [165]),
    .QN(_27707_));
 DFF_X1 _61136_ (.D(_06657_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [171]),
    .QN(_27708_));
 DFF_X1 _61137_ (.D(_06658_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [172]),
    .QN(_27709_));
 DFF_X1 _61138_ (.D(_06659_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [173]),
    .QN(_27710_));
 DFF_X1 _61139_ (.D(_06660_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [174]),
    .QN(_27711_));
 DFF_X1 _61140_ (.D(_06661_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [175]),
    .QN(_27712_));
 DFF_X1 _61141_ (.D(_06662_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [176]),
    .QN(_27713_));
 DFF_X1 _61142_ (.D(_06663_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [177]),
    .QN(_27714_));
 DFF_X1 _61143_ (.D(_06664_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [178]),
    .QN(_27715_));
 DFF_X1 _61144_ (.D(_06665_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [179]),
    .QN(_27716_));
 DFF_X1 _61145_ (.D(_06667_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [180]),
    .QN(_27717_));
 DFF_X1 _61146_ (.D(_06668_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [181]),
    .QN(_27718_));
 DFF_X1 _61147_ (.D(_06669_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [182]),
    .QN(_27719_));
 DFF_X1 _61148_ (.D(_06670_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [183]),
    .QN(_27720_));
 DFF_X1 _61149_ (.D(_06671_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [184]),
    .QN(_27721_));
 DFF_X1 _61150_ (.D(_06672_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [185]),
    .QN(_27722_));
 DFF_X1 _61151_ (.D(_06673_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [186]),
    .QN(_27723_));
 DFF_X1 _61152_ (.D(_06674_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [187]),
    .QN(_27724_));
 DFF_X1 _61153_ (.D(_06675_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [188]),
    .QN(_27725_));
 DFF_X1 _61154_ (.D(_06676_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [189]),
    .QN(_27726_));
 DFF_X1 _61155_ (.D(_06678_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [190]),
    .QN(_27727_));
 DFF_X1 _61156_ (.D(_06679_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [191]),
    .QN(_27728_));
 DFF_X1 _61157_ (.D(_06680_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [192]),
    .QN(_27729_));
 DFF_X1 _61158_ (.D(_06681_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [193]),
    .QN(_27730_));
 DFF_X1 _61159_ (.D(_06682_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [194]),
    .QN(_27731_));
 DFF_X1 _61160_ (.D(_06683_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [195]),
    .QN(_27732_));
 DFF_X1 _61161_ (.D(_06684_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [196]),
    .QN(_27733_));
 DFF_X1 _61162_ (.D(_06685_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [197]),
    .QN(_27734_));
 DFF_X1 _61163_ (.D(_06686_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [198]),
    .QN(_27735_));
 DFF_X1 _61164_ (.D(_06688_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [204]),
    .QN(_27736_));
 DFF_X1 _61165_ (.D(_06689_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [205]),
    .QN(_27737_));
 DFF_X1 _61166_ (.D(_06690_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [206]),
    .QN(_27738_));
 DFF_X1 _61167_ (.D(_06691_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [207]),
    .QN(_27739_));
 DFF_X1 _61168_ (.D(_06692_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [208]),
    .QN(_27740_));
 DFF_X1 _61169_ (.D(_06693_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [209]),
    .QN(_27741_));
 DFF_X1 _61170_ (.D(_06695_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [210]),
    .QN(_27742_));
 DFF_X1 _61171_ (.D(_06696_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [211]),
    .QN(_27743_));
 DFF_X1 _61172_ (.D(_06697_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [212]),
    .QN(_27744_));
 DFF_X1 _61173_ (.D(_06698_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [213]),
    .QN(_27745_));
 DFF_X1 _61174_ (.D(_06699_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [214]),
    .QN(_27746_));
 DFF_X1 _61175_ (.D(_06700_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [215]),
    .QN(_27747_));
 DFF_X1 _61176_ (.D(_06701_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [216]),
    .QN(_27748_));
 DFF_X1 _61177_ (.D(_06702_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [217]),
    .QN(_27749_));
 DFF_X1 _61178_ (.D(_06703_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [218]),
    .QN(_27750_));
 DFF_X1 _61179_ (.D(_06704_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [219]),
    .QN(_27751_));
 DFF_X1 _61180_ (.D(_06706_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [220]),
    .QN(_27752_));
 DFF_X1 _61181_ (.D(_06707_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [221]),
    .QN(_27753_));
 DFF_X1 _61182_ (.D(_06708_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [222]),
    .QN(_27754_));
 DFF_X1 _61183_ (.D(_06709_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [223]),
    .QN(_27755_));
 DFF_X1 _61184_ (.D(_06710_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [224]),
    .QN(_27756_));
 DFF_X1 _61185_ (.D(_06711_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [225]),
    .QN(_27757_));
 DFF_X1 _61186_ (.D(_06712_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [226]),
    .QN(_27758_));
 DFF_X1 _61187_ (.D(_06713_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [227]),
    .QN(_27759_));
 DFF_X1 _61188_ (.D(_06714_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [228]),
    .QN(_27760_));
 DFF_X1 _61189_ (.D(_06715_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [229]),
    .QN(_27761_));
 DFF_X1 _61190_ (.D(_06717_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [230]),
    .QN(_27762_));
 DFF_X1 _61191_ (.D(_06718_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [231]),
    .QN(_27763_));
 DFF_X1 _61192_ (.D(_06719_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [237]),
    .QN(_27764_));
 DFF_X1 _61193_ (.D(_06720_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [238]),
    .QN(_27765_));
 DFF_X1 _61194_ (.D(_06721_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [239]),
    .QN(_27766_));
 DFF_X1 _61195_ (.D(_06723_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [240]),
    .QN(_27767_));
 DFF_X1 _61196_ (.D(_06724_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [241]),
    .QN(_27768_));
 DFF_X1 _61197_ (.D(_06725_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [242]),
    .QN(_27769_));
 DFF_X1 _61198_ (.D(_06726_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [243]),
    .QN(_27770_));
 DFF_X1 _61199_ (.D(_06727_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [244]),
    .QN(_27771_));
 DFF_X1 _61200_ (.D(_06728_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [245]),
    .QN(_27772_));
 DFF_X1 _61201_ (.D(_06729_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [246]),
    .QN(_27773_));
 DFF_X1 _61202_ (.D(_06730_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [247]),
    .QN(_27774_));
 DFF_X1 _61203_ (.D(_06731_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [248]),
    .QN(_27775_));
 DFF_X1 _61204_ (.D(_06732_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [249]),
    .QN(_27776_));
 DFF_X1 _61205_ (.D(_06734_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [250]),
    .QN(_27777_));
 DFF_X1 _61206_ (.D(_06735_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [251]),
    .QN(_27778_));
 DFF_X1 _61207_ (.D(_06736_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [252]),
    .QN(_27779_));
 DFF_X1 _61208_ (.D(_06737_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [253]),
    .QN(_27780_));
 DFF_X1 _61209_ (.D(_06738_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [254]),
    .QN(_27781_));
 DFF_X1 _61210_ (.D(_06739_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [255]),
    .QN(_27782_));
 DFF_X1 _61211_ (.D(_06740_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [256]),
    .QN(_27783_));
 DFF_X1 _61212_ (.D(_06741_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [257]),
    .QN(_27784_));
 DFF_X1 _61213_ (.D(_06742_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [258]),
    .QN(_27785_));
 DFF_X1 _61214_ (.D(_06743_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [259]),
    .QN(_27786_));
 DFF_X1 _61215_ (.D(_06745_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [260]),
    .QN(_27787_));
 DFF_X1 _61216_ (.D(_06746_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [261]),
    .QN(_27788_));
 DFF_X1 _61217_ (.D(_06747_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [262]),
    .QN(_27789_));
 DFF_X1 _61218_ (.D(_06748_),
    .CK(clk_i),
    .Q(\itlb.entry_ram.z_s1r1w_mem.synth.mem [263]),
    .QN(_27790_));
 DFF_X1 _61219_ (.D(\icache.lce.lce_cmd_inst.rv_adapter.N14 ),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.full_r ),
    .QN(lce_cmd_ready_o));
 DFF_X1 _61220_ (.D(\icache.lce.lce_cmd_inst.rv_adapter.N13 ),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.empty_r ),
    .QN(_00001_));
 DFF_X1 _61221_ (.D(_05406_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.head_r ),
    .QN(_27791_));
 DFF_X1 _61222_ (.D(_05407_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.w_addr_i ),
    .QN(_27792_));
 DFF_X1 _61223_ (.D(\icache.lce.lce_data_cmd.rv_adapter.N14 ),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.full_r ),
    .QN(lce_data_cmd_ready_o));
 DFF_X1 _61224_ (.D(\icache.lce.lce_data_cmd.rv_adapter.N13 ),
    .CK(clk_i),
    .Q(\icache.lce.N14 ),
    .QN(_00075_));
 DFF_X1 _61225_ (.D(_05512_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.head_r ),
    .QN(_27793_));
 DFF_X1 _61226_ (.D(_05513_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.w_addr_i ),
    .QN(_27794_));
 DFF_X1 _61227_ (.D(_00822_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [0]),
    .QN(_27795_));
 DFF_X1 _61228_ (.D(_01933_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1]),
    .QN(_27796_));
 DFF_X1 _61229_ (.D(_03044_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2]),
    .QN(_27797_));
 DFF_X1 _61230_ (.D(_03291_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3]),
    .QN(_27798_));
 DFF_X1 _61231_ (.D(_03402_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [4]),
    .QN(_27799_));
 DFF_X1 _61232_ (.D(_03513_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [5]),
    .QN(_27800_));
 DFF_X1 _61233_ (.D(_03624_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [6]),
    .QN(_27801_));
 DFF_X1 _61234_ (.D(_03735_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [7]),
    .QN(_27802_));
 DFF_X1 _61235_ (.D(_03846_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [8]),
    .QN(_27803_));
 DFF_X1 _61236_ (.D(_03957_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [9]),
    .QN(_27804_));
 DFF_X1 _61237_ (.D(_00933_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [10]),
    .QN(_27805_));
 DFF_X1 _61238_ (.D(_01044_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [11]),
    .QN(_27806_));
 DFF_X1 _61239_ (.D(_01155_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [12]),
    .QN(_27807_));
 DFF_X1 _61240_ (.D(_01266_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [13]),
    .QN(_27808_));
 DFF_X1 _61241_ (.D(_01377_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [14]),
    .QN(_27809_));
 DFF_X1 _61242_ (.D(_01488_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [15]),
    .QN(_27810_));
 DFF_X1 _61243_ (.D(_01599_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [16]),
    .QN(_27811_));
 DFF_X1 _61244_ (.D(_01710_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [17]),
    .QN(_27812_));
 DFF_X1 _61245_ (.D(_01821_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [18]),
    .QN(_27813_));
 DFF_X1 _61246_ (.D(_01932_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [19]),
    .QN(_27814_));
 DFF_X1 _61247_ (.D(_02044_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [20]),
    .QN(_27815_));
 DFF_X1 _61248_ (.D(_02155_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [21]),
    .QN(_27816_));
 DFF_X1 _61249_ (.D(_02266_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [22]),
    .QN(_27817_));
 DFF_X1 _61250_ (.D(_02377_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [23]),
    .QN(_27818_));
 DFF_X1 _61251_ (.D(_02488_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [24]),
    .QN(_27819_));
 DFF_X1 _61252_ (.D(_02599_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [25]),
    .QN(_27820_));
 DFF_X1 _61253_ (.D(_02710_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [26]),
    .QN(_27821_));
 DFF_X1 _61254_ (.D(_02821_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [27]),
    .QN(_27822_));
 DFF_X1 _61255_ (.D(_02932_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [28]),
    .QN(_27823_));
 DFF_X1 _61256_ (.D(_03043_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [29]),
    .QN(_27824_));
 DFF_X1 _61257_ (.D(_03155_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [30]),
    .QN(_27825_));
 DFF_X1 _61258_ (.D(_03202_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [31]),
    .QN(_27826_));
 DFF_X1 _61259_ (.D(_03213_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [32]),
    .QN(_27827_));
 DFF_X1 _61260_ (.D(_03224_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [33]),
    .QN(_27828_));
 DFF_X1 _61261_ (.D(_03235_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [34]),
    .QN(_27829_));
 DFF_X1 _61262_ (.D(_03246_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [35]),
    .QN(_27830_));
 DFF_X1 _61263_ (.D(_03257_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [36]),
    .QN(_27831_));
 DFF_X1 _61264_ (.D(_03268_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [37]),
    .QN(_27832_));
 DFF_X1 _61265_ (.D(_03279_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [38]),
    .QN(_27833_));
 DFF_X1 _61266_ (.D(_03290_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [39]),
    .QN(_27834_));
 DFF_X1 _61267_ (.D(_03302_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [40]),
    .QN(_27835_));
 DFF_X1 _61268_ (.D(_03313_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [41]),
    .QN(_27836_));
 DFF_X1 _61269_ (.D(_03324_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [42]),
    .QN(_27837_));
 DFF_X1 _61270_ (.D(_03335_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [43]),
    .QN(_27838_));
 DFF_X1 _61271_ (.D(_03346_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [44]),
    .QN(_27839_));
 DFF_X1 _61272_ (.D(_03357_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [45]),
    .QN(_27840_));
 DFF_X1 _61273_ (.D(_03368_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [46]),
    .QN(_27841_));
 DFF_X1 _61274_ (.D(_03379_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [47]),
    .QN(_27842_));
 DFF_X1 _61275_ (.D(_03390_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [48]),
    .QN(_27843_));
 DFF_X1 _61276_ (.D(_03401_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [49]),
    .QN(_27844_));
 DFF_X1 _61277_ (.D(_03413_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [50]),
    .QN(_27845_));
 DFF_X1 _61278_ (.D(_03424_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [51]),
    .QN(_27846_));
 DFF_X1 _61279_ (.D(_03435_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [52]),
    .QN(_27847_));
 DFF_X1 _61280_ (.D(_03446_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [53]),
    .QN(_27848_));
 DFF_X1 _61281_ (.D(_03457_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [54]),
    .QN(_27849_));
 DFF_X1 _61282_ (.D(_03468_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [55]),
    .QN(_27850_));
 DFF_X1 _61283_ (.D(_03479_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [56]),
    .QN(_27851_));
 DFF_X1 _61284_ (.D(_03490_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [57]),
    .QN(_27852_));
 DFF_X1 _61285_ (.D(_03501_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [58]),
    .QN(_27853_));
 DFF_X1 _61286_ (.D(_03512_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [59]),
    .QN(_27854_));
 DFF_X1 _61287_ (.D(_03524_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [60]),
    .QN(_27855_));
 DFF_X1 _61288_ (.D(_03535_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [61]),
    .QN(_27856_));
 DFF_X1 _61289_ (.D(_03546_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [62]),
    .QN(_27857_));
 DFF_X1 _61290_ (.D(_03557_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [63]),
    .QN(_27858_));
 DFF_X1 _61291_ (.D(_03568_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [64]),
    .QN(_27859_));
 DFF_X1 _61292_ (.D(_03579_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [65]),
    .QN(_27860_));
 DFF_X1 _61293_ (.D(_03590_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [66]),
    .QN(_27861_));
 DFF_X1 _61294_ (.D(_03601_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [67]),
    .QN(_27862_));
 DFF_X1 _61295_ (.D(_03612_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [68]),
    .QN(_27863_));
 DFF_X1 _61296_ (.D(_03623_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [69]),
    .QN(_27864_));
 DFF_X1 _61297_ (.D(_03635_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [70]),
    .QN(_27865_));
 DFF_X1 _61298_ (.D(_03646_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [71]),
    .QN(_27866_));
 DFF_X1 _61299_ (.D(_03657_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [72]),
    .QN(_27867_));
 DFF_X1 _61300_ (.D(_03668_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [73]),
    .QN(_27868_));
 DFF_X1 _61301_ (.D(_03679_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [74]),
    .QN(_27869_));
 DFF_X1 _61302_ (.D(_03690_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [75]),
    .QN(_27870_));
 DFF_X1 _61303_ (.D(_03701_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [76]),
    .QN(_27871_));
 DFF_X1 _61304_ (.D(_03712_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [77]),
    .QN(_27872_));
 DFF_X1 _61305_ (.D(_03723_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [78]),
    .QN(_27873_));
 DFF_X1 _61306_ (.D(_03734_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [79]),
    .QN(_27874_));
 DFF_X1 _61307_ (.D(_03746_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [80]),
    .QN(_27875_));
 DFF_X1 _61308_ (.D(_03757_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [81]),
    .QN(_27876_));
 DFF_X1 _61309_ (.D(_03768_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [82]),
    .QN(_27877_));
 DFF_X1 _61310_ (.D(_03779_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [83]),
    .QN(_27878_));
 DFF_X1 _61311_ (.D(_03790_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [84]),
    .QN(_27879_));
 DFF_X1 _61312_ (.D(_03801_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [85]),
    .QN(_27880_));
 DFF_X1 _61313_ (.D(_03812_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [86]),
    .QN(_27881_));
 DFF_X1 _61314_ (.D(_03823_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [87]),
    .QN(_27882_));
 DFF_X1 _61315_ (.D(_03834_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [88]),
    .QN(_27883_));
 DFF_X1 _61316_ (.D(_03845_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [89]),
    .QN(_27884_));
 DFF_X1 _61317_ (.D(_03857_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [90]),
    .QN(_27885_));
 DFF_X1 _61318_ (.D(_03868_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [91]),
    .QN(_27886_));
 DFF_X1 _61319_ (.D(_03879_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [92]),
    .QN(_27887_));
 DFF_X1 _61320_ (.D(_03890_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [93]),
    .QN(_27888_));
 DFF_X1 _61321_ (.D(_03901_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [94]),
    .QN(_27889_));
 DFF_X1 _61322_ (.D(_03912_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [95]),
    .QN(_27890_));
 DFF_X1 _61323_ (.D(_03923_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [96]),
    .QN(_27891_));
 DFF_X1 _61324_ (.D(_03934_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [97]),
    .QN(_27892_));
 DFF_X1 _61325_ (.D(_03945_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [98]),
    .QN(_27893_));
 DFF_X1 _61326_ (.D(_03956_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [99]),
    .QN(_27894_));
 DFF_X1 _61327_ (.D(_00833_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [100]),
    .QN(_27895_));
 DFF_X1 _61328_ (.D(_00844_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [101]),
    .QN(_27896_));
 DFF_X1 _61329_ (.D(_00855_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [102]),
    .QN(_27897_));
 DFF_X1 _61330_ (.D(_00866_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [103]),
    .QN(_27898_));
 DFF_X1 _61331_ (.D(_00877_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [104]),
    .QN(_27899_));
 DFF_X1 _61332_ (.D(_00888_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [105]),
    .QN(_27900_));
 DFF_X1 _61333_ (.D(_00899_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [106]),
    .QN(_27901_));
 DFF_X1 _61334_ (.D(_00910_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [107]),
    .QN(_27902_));
 DFF_X1 _61335_ (.D(_00921_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [108]),
    .QN(_27903_));
 DFF_X1 _61336_ (.D(_00932_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [109]),
    .QN(_27904_));
 DFF_X1 _61337_ (.D(_00944_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [110]),
    .QN(_27905_));
 DFF_X1 _61338_ (.D(_00955_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [111]),
    .QN(_27906_));
 DFF_X1 _61339_ (.D(_00966_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [112]),
    .QN(_27907_));
 DFF_X1 _61340_ (.D(_00977_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [113]),
    .QN(_27908_));
 DFF_X1 _61341_ (.D(_00988_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [114]),
    .QN(_27909_));
 DFF_X1 _61342_ (.D(_00999_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [115]),
    .QN(_27910_));
 DFF_X1 _61343_ (.D(_01010_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [116]),
    .QN(_27911_));
 DFF_X1 _61344_ (.D(_01021_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [117]),
    .QN(_27912_));
 DFF_X1 _61345_ (.D(_01032_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [118]),
    .QN(_27913_));
 DFF_X1 _61346_ (.D(_01043_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [119]),
    .QN(_27914_));
 DFF_X1 _61347_ (.D(_01055_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [120]),
    .QN(_27915_));
 DFF_X1 _61348_ (.D(_01066_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [121]),
    .QN(_27916_));
 DFF_X1 _61349_ (.D(_01077_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [122]),
    .QN(_27917_));
 DFF_X1 _61350_ (.D(_01088_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [123]),
    .QN(_27918_));
 DFF_X1 _61351_ (.D(_01099_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [124]),
    .QN(_27919_));
 DFF_X1 _61352_ (.D(_01110_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [125]),
    .QN(_27920_));
 DFF_X1 _61353_ (.D(_01121_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [126]),
    .QN(_27921_));
 DFF_X1 _61354_ (.D(_01132_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [127]),
    .QN(_27922_));
 DFF_X1 _61355_ (.D(_01143_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [128]),
    .QN(_27923_));
 DFF_X1 _61356_ (.D(_01154_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [129]),
    .QN(_27924_));
 DFF_X1 _61357_ (.D(_01166_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [130]),
    .QN(_27925_));
 DFF_X1 _61358_ (.D(_01177_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [131]),
    .QN(_27926_));
 DFF_X1 _61359_ (.D(_01188_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [132]),
    .QN(_27927_));
 DFF_X1 _61360_ (.D(_01199_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [133]),
    .QN(_27928_));
 DFF_X1 _61361_ (.D(_01210_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [134]),
    .QN(_27929_));
 DFF_X1 _61362_ (.D(_01221_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [135]),
    .QN(_27930_));
 DFF_X1 _61363_ (.D(_01232_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [136]),
    .QN(_27931_));
 DFF_X1 _61364_ (.D(_01243_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [137]),
    .QN(_27932_));
 DFF_X1 _61365_ (.D(_01254_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [138]),
    .QN(_27933_));
 DFF_X1 _61366_ (.D(_01265_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [139]),
    .QN(_27934_));
 DFF_X1 _61367_ (.D(_01277_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [140]),
    .QN(_27935_));
 DFF_X1 _61368_ (.D(_01288_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [141]),
    .QN(_27936_));
 DFF_X1 _61369_ (.D(_01299_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [142]),
    .QN(_27937_));
 DFF_X1 _61370_ (.D(_01310_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [143]),
    .QN(_27938_));
 DFF_X1 _61371_ (.D(_01321_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [144]),
    .QN(_27939_));
 DFF_X1 _61372_ (.D(_01332_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [145]),
    .QN(_27940_));
 DFF_X1 _61373_ (.D(_01343_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [146]),
    .QN(_27941_));
 DFF_X1 _61374_ (.D(_01354_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [147]),
    .QN(_27942_));
 DFF_X1 _61375_ (.D(_01365_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [148]),
    .QN(_27943_));
 DFF_X1 _61376_ (.D(_01376_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [149]),
    .QN(_27944_));
 DFF_X1 _61377_ (.D(_01388_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [150]),
    .QN(_27945_));
 DFF_X1 _61378_ (.D(_01399_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [151]),
    .QN(_27946_));
 DFF_X1 _61379_ (.D(_01410_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [152]),
    .QN(_27947_));
 DFF_X1 _61380_ (.D(_01421_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [153]),
    .QN(_27948_));
 DFF_X1 _61381_ (.D(_01432_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [154]),
    .QN(_27949_));
 DFF_X1 _61382_ (.D(_01443_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [155]),
    .QN(_27950_));
 DFF_X1 _61383_ (.D(_01454_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [156]),
    .QN(_27951_));
 DFF_X1 _61384_ (.D(_01465_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [157]),
    .QN(_27952_));
 DFF_X1 _61385_ (.D(_01476_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [158]),
    .QN(_27953_));
 DFF_X1 _61386_ (.D(_01487_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [159]),
    .QN(_27954_));
 DFF_X1 _61387_ (.D(_01499_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [160]),
    .QN(_27955_));
 DFF_X1 _61388_ (.D(_01510_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [161]),
    .QN(_27956_));
 DFF_X1 _61389_ (.D(_01521_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [162]),
    .QN(_27957_));
 DFF_X1 _61390_ (.D(_01532_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [163]),
    .QN(_27958_));
 DFF_X1 _61391_ (.D(_01543_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [164]),
    .QN(_27959_));
 DFF_X1 _61392_ (.D(_01554_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [165]),
    .QN(_27960_));
 DFF_X1 _61393_ (.D(_01565_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [166]),
    .QN(_27961_));
 DFF_X1 _61394_ (.D(_01576_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [167]),
    .QN(_27962_));
 DFF_X1 _61395_ (.D(_01587_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [168]),
    .QN(_27963_));
 DFF_X1 _61396_ (.D(_01598_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [169]),
    .QN(_27964_));
 DFF_X1 _61397_ (.D(_01610_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [170]),
    .QN(_27965_));
 DFF_X1 _61398_ (.D(_01621_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [171]),
    .QN(_27966_));
 DFF_X1 _61399_ (.D(_01632_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [172]),
    .QN(_27967_));
 DFF_X1 _61400_ (.D(_01643_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [173]),
    .QN(_27968_));
 DFF_X1 _61401_ (.D(_01654_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [174]),
    .QN(_27969_));
 DFF_X1 _61402_ (.D(_01665_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [175]),
    .QN(_27970_));
 DFF_X1 _61403_ (.D(_01676_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [176]),
    .QN(_27971_));
 DFF_X1 _61404_ (.D(_01687_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [177]),
    .QN(_27972_));
 DFF_X1 _61405_ (.D(_01698_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [178]),
    .QN(_27973_));
 DFF_X1 _61406_ (.D(_01709_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [179]),
    .QN(_27974_));
 DFF_X1 _61407_ (.D(_01721_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [180]),
    .QN(_27975_));
 DFF_X1 _61408_ (.D(_01732_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [181]),
    .QN(_27976_));
 DFF_X1 _61409_ (.D(_01743_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [182]),
    .QN(_27977_));
 DFF_X1 _61410_ (.D(_01754_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [183]),
    .QN(_27978_));
 DFF_X1 _61411_ (.D(_01765_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [184]),
    .QN(_27979_));
 DFF_X1 _61412_ (.D(_01776_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [185]),
    .QN(_27980_));
 DFF_X1 _61413_ (.D(_01787_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [186]),
    .QN(_27981_));
 DFF_X1 _61414_ (.D(_01798_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [187]),
    .QN(_27982_));
 DFF_X1 _61415_ (.D(_01809_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [188]),
    .QN(_27983_));
 DFF_X1 _61416_ (.D(_01820_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [189]),
    .QN(_27984_));
 DFF_X1 _61417_ (.D(_01832_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [190]),
    .QN(_27985_));
 DFF_X1 _61418_ (.D(_01843_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [191]),
    .QN(_27986_));
 DFF_X1 _61419_ (.D(_01854_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [192]),
    .QN(_27987_));
 DFF_X1 _61420_ (.D(_01865_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [193]),
    .QN(_27988_));
 DFF_X1 _61421_ (.D(_01876_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [194]),
    .QN(_27989_));
 DFF_X1 _61422_ (.D(_01887_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [195]),
    .QN(_27990_));
 DFF_X1 _61423_ (.D(_01898_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [196]),
    .QN(_27991_));
 DFF_X1 _61424_ (.D(_01909_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [197]),
    .QN(_27992_));
 DFF_X1 _61425_ (.D(_01920_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [198]),
    .QN(_27993_));
 DFF_X1 _61426_ (.D(_01931_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [199]),
    .QN(_27994_));
 DFF_X1 _61427_ (.D(_01944_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [200]),
    .QN(_27995_));
 DFF_X1 _61428_ (.D(_01955_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [201]),
    .QN(_27996_));
 DFF_X1 _61429_ (.D(_01966_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [202]),
    .QN(_27997_));
 DFF_X1 _61430_ (.D(_01977_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [203]),
    .QN(_27998_));
 DFF_X1 _61431_ (.D(_01988_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [204]),
    .QN(_27999_));
 DFF_X1 _61432_ (.D(_01999_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [205]),
    .QN(_28000_));
 DFF_X1 _61433_ (.D(_02010_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [206]),
    .QN(_28001_));
 DFF_X1 _61434_ (.D(_02021_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [207]),
    .QN(_28002_));
 DFF_X1 _61435_ (.D(_02032_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [208]),
    .QN(_28003_));
 DFF_X1 _61436_ (.D(_02043_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [209]),
    .QN(_28004_));
 DFF_X1 _61437_ (.D(_02055_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [210]),
    .QN(_28005_));
 DFF_X1 _61438_ (.D(_02066_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [211]),
    .QN(_28006_));
 DFF_X1 _61439_ (.D(_02077_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [212]),
    .QN(_28007_));
 DFF_X1 _61440_ (.D(_02088_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [213]),
    .QN(_28008_));
 DFF_X1 _61441_ (.D(_02099_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [214]),
    .QN(_28009_));
 DFF_X1 _61442_ (.D(_02110_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [215]),
    .QN(_28010_));
 DFF_X1 _61443_ (.D(_02121_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [216]),
    .QN(_28011_));
 DFF_X1 _61444_ (.D(_02132_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [217]),
    .QN(_28012_));
 DFF_X1 _61445_ (.D(_02143_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [218]),
    .QN(_28013_));
 DFF_X1 _61446_ (.D(_02154_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [219]),
    .QN(_28014_));
 DFF_X1 _61447_ (.D(_02166_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [220]),
    .QN(_28015_));
 DFF_X1 _61448_ (.D(_02177_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [221]),
    .QN(_28016_));
 DFF_X1 _61449_ (.D(_02188_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [222]),
    .QN(_28017_));
 DFF_X1 _61450_ (.D(_02199_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [223]),
    .QN(_28018_));
 DFF_X1 _61451_ (.D(_02210_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [224]),
    .QN(_28019_));
 DFF_X1 _61452_ (.D(_02221_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [225]),
    .QN(_28020_));
 DFF_X1 _61453_ (.D(_02232_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [226]),
    .QN(_28021_));
 DFF_X1 _61454_ (.D(_02243_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [227]),
    .QN(_28022_));
 DFF_X1 _61455_ (.D(_02254_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [228]),
    .QN(_28023_));
 DFF_X1 _61456_ (.D(_02265_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [229]),
    .QN(_28024_));
 DFF_X1 _61457_ (.D(_02277_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [230]),
    .QN(_28025_));
 DFF_X1 _61458_ (.D(_02288_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [231]),
    .QN(_28026_));
 DFF_X1 _61459_ (.D(_02299_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [232]),
    .QN(_28027_));
 DFF_X1 _61460_ (.D(_02310_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [233]),
    .QN(_28028_));
 DFF_X1 _61461_ (.D(_02321_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [234]),
    .QN(_28029_));
 DFF_X1 _61462_ (.D(_02332_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [235]),
    .QN(_28030_));
 DFF_X1 _61463_ (.D(_02343_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [236]),
    .QN(_28031_));
 DFF_X1 _61464_ (.D(_02354_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [237]),
    .QN(_28032_));
 DFF_X1 _61465_ (.D(_02365_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [238]),
    .QN(_28033_));
 DFF_X1 _61466_ (.D(_02376_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [239]),
    .QN(_28034_));
 DFF_X1 _61467_ (.D(_02388_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [240]),
    .QN(_28035_));
 DFF_X1 _61468_ (.D(_02399_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [241]),
    .QN(_28036_));
 DFF_X1 _61469_ (.D(_02410_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [242]),
    .QN(_28037_));
 DFF_X1 _61470_ (.D(_02421_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [243]),
    .QN(_28038_));
 DFF_X1 _61471_ (.D(_02432_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [244]),
    .QN(_28039_));
 DFF_X1 _61472_ (.D(_02443_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [245]),
    .QN(_28040_));
 DFF_X1 _61473_ (.D(_02454_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [246]),
    .QN(_28041_));
 DFF_X1 _61474_ (.D(_02465_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [247]),
    .QN(_28042_));
 DFF_X1 _61475_ (.D(_02476_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [248]),
    .QN(_28043_));
 DFF_X1 _61476_ (.D(_02487_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [249]),
    .QN(_28044_));
 DFF_X1 _61477_ (.D(_02499_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [250]),
    .QN(_28045_));
 DFF_X1 _61478_ (.D(_02510_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [251]),
    .QN(_28046_));
 DFF_X1 _61479_ (.D(_02521_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [252]),
    .QN(_28047_));
 DFF_X1 _61480_ (.D(_02532_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [253]),
    .QN(_28048_));
 DFF_X1 _61481_ (.D(_02543_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [254]),
    .QN(_28049_));
 DFF_X1 _61482_ (.D(_02554_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [255]),
    .QN(_28050_));
 DFF_X1 _61483_ (.D(_02565_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [256]),
    .QN(_28051_));
 DFF_X1 _61484_ (.D(_02576_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [257]),
    .QN(_28052_));
 DFF_X1 _61485_ (.D(_02587_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [258]),
    .QN(_28053_));
 DFF_X1 _61486_ (.D(_02598_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [259]),
    .QN(_28054_));
 DFF_X1 _61487_ (.D(_02610_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [260]),
    .QN(_28055_));
 DFF_X1 _61488_ (.D(_02621_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [261]),
    .QN(_28056_));
 DFF_X1 _61489_ (.D(_02632_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [262]),
    .QN(_28057_));
 DFF_X1 _61490_ (.D(_02643_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [263]),
    .QN(_28058_));
 DFF_X1 _61491_ (.D(_02654_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [264]),
    .QN(_28059_));
 DFF_X1 _61492_ (.D(_02665_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [265]),
    .QN(_28060_));
 DFF_X1 _61493_ (.D(_02676_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [266]),
    .QN(_28061_));
 DFF_X1 _61494_ (.D(_02687_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [267]),
    .QN(_28062_));
 DFF_X1 _61495_ (.D(_02698_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [268]),
    .QN(_28063_));
 DFF_X1 _61496_ (.D(_02709_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [269]),
    .QN(_28064_));
 DFF_X1 _61497_ (.D(_02721_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [270]),
    .QN(_28065_));
 DFF_X1 _61498_ (.D(_02732_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [271]),
    .QN(_28066_));
 DFF_X1 _61499_ (.D(_02743_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [272]),
    .QN(_28067_));
 DFF_X1 _61500_ (.D(_02754_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [273]),
    .QN(_28068_));
 DFF_X1 _61501_ (.D(_02765_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [274]),
    .QN(_28069_));
 DFF_X1 _61502_ (.D(_02776_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [275]),
    .QN(_28070_));
 DFF_X1 _61503_ (.D(_02787_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [276]),
    .QN(_28071_));
 DFF_X1 _61504_ (.D(_02798_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [277]),
    .QN(_28072_));
 DFF_X1 _61505_ (.D(_02809_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [278]),
    .QN(_28073_));
 DFF_X1 _61506_ (.D(_02820_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [279]),
    .QN(_28074_));
 DFF_X1 _61507_ (.D(_02832_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [280]),
    .QN(_28075_));
 DFF_X1 _61508_ (.D(_02843_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [281]),
    .QN(_28076_));
 DFF_X1 _61509_ (.D(_02854_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [282]),
    .QN(_28077_));
 DFF_X1 _61510_ (.D(_02865_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [283]),
    .QN(_28078_));
 DFF_X1 _61511_ (.D(_02876_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [284]),
    .QN(_28079_));
 DFF_X1 _61512_ (.D(_02887_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [285]),
    .QN(_28080_));
 DFF_X1 _61513_ (.D(_02898_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [286]),
    .QN(_28081_));
 DFF_X1 _61514_ (.D(_02909_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [287]),
    .QN(_28082_));
 DFF_X1 _61515_ (.D(_02920_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [288]),
    .QN(_28083_));
 DFF_X1 _61516_ (.D(_02931_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [289]),
    .QN(_28084_));
 DFF_X1 _61517_ (.D(_02943_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [290]),
    .QN(_28085_));
 DFF_X1 _61518_ (.D(_02954_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [291]),
    .QN(_28086_));
 DFF_X1 _61519_ (.D(_02965_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [292]),
    .QN(_28087_));
 DFF_X1 _61520_ (.D(_02976_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [293]),
    .QN(_28088_));
 DFF_X1 _61521_ (.D(_02987_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [294]),
    .QN(_28089_));
 DFF_X1 _61522_ (.D(_02998_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [295]),
    .QN(_28090_));
 DFF_X1 _61523_ (.D(_03009_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [296]),
    .QN(_28091_));
 DFF_X1 _61524_ (.D(_03020_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [297]),
    .QN(_28092_));
 DFF_X1 _61525_ (.D(_03031_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [298]),
    .QN(_28093_));
 DFF_X1 _61526_ (.D(_03042_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [299]),
    .QN(_28094_));
 DFF_X1 _61527_ (.D(_03055_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [300]),
    .QN(_28095_));
 DFF_X1 _61528_ (.D(_03066_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [301]),
    .QN(_28096_));
 DFF_X1 _61529_ (.D(_03077_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [302]),
    .QN(_28097_));
 DFF_X1 _61530_ (.D(_03088_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [303]),
    .QN(_28098_));
 DFF_X1 _61531_ (.D(_03099_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [304]),
    .QN(_28099_));
 DFF_X1 _61532_ (.D(_03110_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [305]),
    .QN(_28100_));
 DFF_X1 _61533_ (.D(_03121_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [306]),
    .QN(_28101_));
 DFF_X1 _61534_ (.D(_03132_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [307]),
    .QN(_28102_));
 DFF_X1 _61535_ (.D(_03143_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [308]),
    .QN(_28103_));
 DFF_X1 _61536_ (.D(_03154_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [309]),
    .QN(_28104_));
 DFF_X1 _61537_ (.D(_03166_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [310]),
    .QN(_28105_));
 DFF_X1 _61538_ (.D(_03177_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [311]),
    .QN(_28106_));
 DFF_X1 _61539_ (.D(_03188_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [312]),
    .QN(_28107_));
 DFF_X1 _61540_ (.D(_03195_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [313]),
    .QN(_28108_));
 DFF_X1 _61541_ (.D(_03196_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [314]),
    .QN(_28109_));
 DFF_X1 _61542_ (.D(_03197_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [315]),
    .QN(_28110_));
 DFF_X1 _61543_ (.D(_03198_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [316]),
    .QN(_28111_));
 DFF_X1 _61544_ (.D(_03199_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [317]),
    .QN(_28112_));
 DFF_X1 _61545_ (.D(_03200_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [318]),
    .QN(_28113_));
 DFF_X1 _61546_ (.D(_03201_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [319]),
    .QN(_28114_));
 DFF_X1 _61547_ (.D(_03203_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [320]),
    .QN(_28115_));
 DFF_X1 _61548_ (.D(_03204_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [321]),
    .QN(_28116_));
 DFF_X1 _61549_ (.D(_03205_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [322]),
    .QN(_28117_));
 DFF_X1 _61550_ (.D(_03206_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [323]),
    .QN(_28118_));
 DFF_X1 _61551_ (.D(_03207_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [324]),
    .QN(_28119_));
 DFF_X1 _61552_ (.D(_03208_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [325]),
    .QN(_28120_));
 DFF_X1 _61553_ (.D(_03209_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [326]),
    .QN(_28121_));
 DFF_X1 _61554_ (.D(_03210_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [327]),
    .QN(_28122_));
 DFF_X1 _61555_ (.D(_03211_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [328]),
    .QN(_28123_));
 DFF_X1 _61556_ (.D(_03212_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [329]),
    .QN(_28124_));
 DFF_X1 _61557_ (.D(_03214_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [330]),
    .QN(_28125_));
 DFF_X1 _61558_ (.D(_03215_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [331]),
    .QN(_28126_));
 DFF_X1 _61559_ (.D(_03216_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [332]),
    .QN(_28127_));
 DFF_X1 _61560_ (.D(_03217_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [333]),
    .QN(_28128_));
 DFF_X1 _61561_ (.D(_03218_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [334]),
    .QN(_28129_));
 DFF_X1 _61562_ (.D(_03219_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [335]),
    .QN(_28130_));
 DFF_X1 _61563_ (.D(_03220_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [336]),
    .QN(_28131_));
 DFF_X1 _61564_ (.D(_03221_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [337]),
    .QN(_28132_));
 DFF_X1 _61565_ (.D(_03222_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [338]),
    .QN(_28133_));
 DFF_X1 _61566_ (.D(_03223_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [339]),
    .QN(_28134_));
 DFF_X1 _61567_ (.D(_03225_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [340]),
    .QN(_28135_));
 DFF_X1 _61568_ (.D(_03226_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [341]),
    .QN(_28136_));
 DFF_X1 _61569_ (.D(_03227_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [342]),
    .QN(_28137_));
 DFF_X1 _61570_ (.D(_03228_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [343]),
    .QN(_28138_));
 DFF_X1 _61571_ (.D(_03229_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [344]),
    .QN(_28139_));
 DFF_X1 _61572_ (.D(_03230_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [345]),
    .QN(_28140_));
 DFF_X1 _61573_ (.D(_03231_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [346]),
    .QN(_28141_));
 DFF_X1 _61574_ (.D(_03232_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [347]),
    .QN(_28142_));
 DFF_X1 _61575_ (.D(_03233_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [348]),
    .QN(_28143_));
 DFF_X1 _61576_ (.D(_03234_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [349]),
    .QN(_28144_));
 DFF_X1 _61577_ (.D(_03236_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [350]),
    .QN(_28145_));
 DFF_X1 _61578_ (.D(_03237_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [351]),
    .QN(_28146_));
 DFF_X1 _61579_ (.D(_03238_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [352]),
    .QN(_28147_));
 DFF_X1 _61580_ (.D(_03239_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [353]),
    .QN(_28148_));
 DFF_X1 _61581_ (.D(_03240_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [354]),
    .QN(_28149_));
 DFF_X1 _61582_ (.D(_03241_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [355]),
    .QN(_28150_));
 DFF_X1 _61583_ (.D(_03242_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [356]),
    .QN(_28151_));
 DFF_X1 _61584_ (.D(_03243_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [357]),
    .QN(_28152_));
 DFF_X1 _61585_ (.D(_03244_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [358]),
    .QN(_28153_));
 DFF_X1 _61586_ (.D(_03245_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [359]),
    .QN(_28154_));
 DFF_X1 _61587_ (.D(_03247_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [360]),
    .QN(_28155_));
 DFF_X1 _61588_ (.D(_03248_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [361]),
    .QN(_28156_));
 DFF_X1 _61589_ (.D(_03249_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [362]),
    .QN(_28157_));
 DFF_X1 _61590_ (.D(_03250_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [363]),
    .QN(_28158_));
 DFF_X1 _61591_ (.D(_03251_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [364]),
    .QN(_28159_));
 DFF_X1 _61592_ (.D(_03252_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [365]),
    .QN(_28160_));
 DFF_X1 _61593_ (.D(_03253_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [366]),
    .QN(_28161_));
 DFF_X1 _61594_ (.D(_03254_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [367]),
    .QN(_28162_));
 DFF_X1 _61595_ (.D(_03255_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [368]),
    .QN(_28163_));
 DFF_X1 _61596_ (.D(_03256_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [369]),
    .QN(_28164_));
 DFF_X1 _61597_ (.D(_03258_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [370]),
    .QN(_28165_));
 DFF_X1 _61598_ (.D(_03259_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [371]),
    .QN(_28166_));
 DFF_X1 _61599_ (.D(_03260_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [372]),
    .QN(_28167_));
 DFF_X1 _61600_ (.D(_03261_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [373]),
    .QN(_28168_));
 DFF_X1 _61601_ (.D(_03262_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [374]),
    .QN(_28169_));
 DFF_X1 _61602_ (.D(_03263_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [375]),
    .QN(_28170_));
 DFF_X1 _61603_ (.D(_03264_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [376]),
    .QN(_28171_));
 DFF_X1 _61604_ (.D(_03265_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [377]),
    .QN(_28172_));
 DFF_X1 _61605_ (.D(_03266_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [378]),
    .QN(_28173_));
 DFF_X1 _61606_ (.D(_03267_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [379]),
    .QN(_28174_));
 DFF_X1 _61607_ (.D(_03269_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [380]),
    .QN(_28175_));
 DFF_X1 _61608_ (.D(_03270_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [381]),
    .QN(_28176_));
 DFF_X1 _61609_ (.D(_03271_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [382]),
    .QN(_28177_));
 DFF_X1 _61610_ (.D(_03272_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [383]),
    .QN(_28178_));
 DFF_X1 _61611_ (.D(_03273_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [384]),
    .QN(_28179_));
 DFF_X1 _61612_ (.D(_03274_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [385]),
    .QN(_28180_));
 DFF_X1 _61613_ (.D(_03275_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [386]),
    .QN(_28181_));
 DFF_X1 _61614_ (.D(_03276_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [387]),
    .QN(_28182_));
 DFF_X1 _61615_ (.D(_03277_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [388]),
    .QN(_28183_));
 DFF_X1 _61616_ (.D(_03278_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [389]),
    .QN(_28184_));
 DFF_X1 _61617_ (.D(_03280_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [390]),
    .QN(_28185_));
 DFF_X1 _61618_ (.D(_03281_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [391]),
    .QN(_28186_));
 DFF_X1 _61619_ (.D(_03282_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [392]),
    .QN(_28187_));
 DFF_X1 _61620_ (.D(_03283_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [393]),
    .QN(_28188_));
 DFF_X1 _61621_ (.D(_03284_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [394]),
    .QN(_28189_));
 DFF_X1 _61622_ (.D(_03285_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [395]),
    .QN(_28190_));
 DFF_X1 _61623_ (.D(_03286_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [396]),
    .QN(_28191_));
 DFF_X1 _61624_ (.D(_03287_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [397]),
    .QN(_28192_));
 DFF_X1 _61625_ (.D(_03288_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [398]),
    .QN(_28193_));
 DFF_X1 _61626_ (.D(_03289_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [399]),
    .QN(_28194_));
 DFF_X1 _61627_ (.D(_03292_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [400]),
    .QN(_28195_));
 DFF_X1 _61628_ (.D(_03293_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [401]),
    .QN(_28196_));
 DFF_X1 _61629_ (.D(_03294_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [402]),
    .QN(_28197_));
 DFF_X1 _61630_ (.D(_03295_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [403]),
    .QN(_28198_));
 DFF_X1 _61631_ (.D(_03296_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [404]),
    .QN(_28199_));
 DFF_X1 _61632_ (.D(_03297_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [405]),
    .QN(_28200_));
 DFF_X1 _61633_ (.D(_03298_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [406]),
    .QN(_28201_));
 DFF_X1 _61634_ (.D(_03299_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [407]),
    .QN(_28202_));
 DFF_X1 _61635_ (.D(_03300_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [408]),
    .QN(_28203_));
 DFF_X1 _61636_ (.D(_03301_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [409]),
    .QN(_28204_));
 DFF_X1 _61637_ (.D(_03303_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [410]),
    .QN(_28205_));
 DFF_X1 _61638_ (.D(_03304_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [411]),
    .QN(_28206_));
 DFF_X1 _61639_ (.D(_03305_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [412]),
    .QN(_28207_));
 DFF_X1 _61640_ (.D(_03306_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [413]),
    .QN(_28208_));
 DFF_X1 _61641_ (.D(_03307_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [414]),
    .QN(_28209_));
 DFF_X1 _61642_ (.D(_03308_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [415]),
    .QN(_28210_));
 DFF_X1 _61643_ (.D(_03309_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [416]),
    .QN(_28211_));
 DFF_X1 _61644_ (.D(_03310_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [417]),
    .QN(_28212_));
 DFF_X1 _61645_ (.D(_03311_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [418]),
    .QN(_28213_));
 DFF_X1 _61646_ (.D(_03312_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [419]),
    .QN(_28214_));
 DFF_X1 _61647_ (.D(_03314_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [420]),
    .QN(_28215_));
 DFF_X1 _61648_ (.D(_03315_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [421]),
    .QN(_28216_));
 DFF_X1 _61649_ (.D(_03316_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [422]),
    .QN(_28217_));
 DFF_X1 _61650_ (.D(_03317_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [423]),
    .QN(_28218_));
 DFF_X1 _61651_ (.D(_03318_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [424]),
    .QN(_28219_));
 DFF_X1 _61652_ (.D(_03319_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [425]),
    .QN(_28220_));
 DFF_X1 _61653_ (.D(_03320_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [426]),
    .QN(_28221_));
 DFF_X1 _61654_ (.D(_03321_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [427]),
    .QN(_28222_));
 DFF_X1 _61655_ (.D(_03322_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [428]),
    .QN(_28223_));
 DFF_X1 _61656_ (.D(_03323_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [429]),
    .QN(_28224_));
 DFF_X1 _61657_ (.D(_03325_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [430]),
    .QN(_28225_));
 DFF_X1 _61658_ (.D(_03326_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [431]),
    .QN(_28226_));
 DFF_X1 _61659_ (.D(_03327_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [432]),
    .QN(_28227_));
 DFF_X1 _61660_ (.D(_03328_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [433]),
    .QN(_28228_));
 DFF_X1 _61661_ (.D(_03329_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [434]),
    .QN(_28229_));
 DFF_X1 _61662_ (.D(_03330_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [435]),
    .QN(_28230_));
 DFF_X1 _61663_ (.D(_03331_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [436]),
    .QN(_28231_));
 DFF_X1 _61664_ (.D(_03332_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [437]),
    .QN(_28232_));
 DFF_X1 _61665_ (.D(_03333_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [438]),
    .QN(_28233_));
 DFF_X1 _61666_ (.D(_03334_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [439]),
    .QN(_28234_));
 DFF_X1 _61667_ (.D(_03336_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [440]),
    .QN(_28235_));
 DFF_X1 _61668_ (.D(_03337_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [441]),
    .QN(_28236_));
 DFF_X1 _61669_ (.D(_03338_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [442]),
    .QN(_28237_));
 DFF_X1 _61670_ (.D(_03339_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [443]),
    .QN(_28238_));
 DFF_X1 _61671_ (.D(_03340_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [444]),
    .QN(_28239_));
 DFF_X1 _61672_ (.D(_03341_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [445]),
    .QN(_28240_));
 DFF_X1 _61673_ (.D(_03342_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [446]),
    .QN(_28241_));
 DFF_X1 _61674_ (.D(_03343_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [447]),
    .QN(_28242_));
 DFF_X1 _61675_ (.D(_03344_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [448]),
    .QN(_28243_));
 DFF_X1 _61676_ (.D(_03345_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [449]),
    .QN(_28244_));
 DFF_X1 _61677_ (.D(_03347_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [450]),
    .QN(_28245_));
 DFF_X1 _61678_ (.D(_03348_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [451]),
    .QN(_28246_));
 DFF_X1 _61679_ (.D(_03349_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [452]),
    .QN(_28247_));
 DFF_X1 _61680_ (.D(_03350_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [453]),
    .QN(_28248_));
 DFF_X1 _61681_ (.D(_03351_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [454]),
    .QN(_28249_));
 DFF_X1 _61682_ (.D(_03352_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [455]),
    .QN(_28250_));
 DFF_X1 _61683_ (.D(_03353_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [456]),
    .QN(_28251_));
 DFF_X1 _61684_ (.D(_03354_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [457]),
    .QN(_28252_));
 DFF_X1 _61685_ (.D(_03355_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [458]),
    .QN(_28253_));
 DFF_X1 _61686_ (.D(_03356_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [459]),
    .QN(_28254_));
 DFF_X1 _61687_ (.D(_03358_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [460]),
    .QN(_28255_));
 DFF_X1 _61688_ (.D(_03359_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [461]),
    .QN(_28256_));
 DFF_X1 _61689_ (.D(_03360_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [462]),
    .QN(_28257_));
 DFF_X1 _61690_ (.D(_03361_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [463]),
    .QN(_28258_));
 DFF_X1 _61691_ (.D(_03362_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [464]),
    .QN(_28259_));
 DFF_X1 _61692_ (.D(_03363_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [465]),
    .QN(_28260_));
 DFF_X1 _61693_ (.D(_03364_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [466]),
    .QN(_28261_));
 DFF_X1 _61694_ (.D(_03365_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [467]),
    .QN(_28262_));
 DFF_X1 _61695_ (.D(_03366_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [468]),
    .QN(_28263_));
 DFF_X1 _61696_ (.D(_03367_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [469]),
    .QN(_28264_));
 DFF_X1 _61697_ (.D(_03369_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [470]),
    .QN(_28265_));
 DFF_X1 _61698_ (.D(_03370_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [471]),
    .QN(_28266_));
 DFF_X1 _61699_ (.D(_03371_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [472]),
    .QN(_28267_));
 DFF_X1 _61700_ (.D(_03372_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [473]),
    .QN(_28268_));
 DFF_X1 _61701_ (.D(_03373_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [474]),
    .QN(_28269_));
 DFF_X1 _61702_ (.D(_03374_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [475]),
    .QN(_28270_));
 DFF_X1 _61703_ (.D(_03375_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [476]),
    .QN(_28271_));
 DFF_X1 _61704_ (.D(_03376_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [477]),
    .QN(_28272_));
 DFF_X1 _61705_ (.D(_03377_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [478]),
    .QN(_28273_));
 DFF_X1 _61706_ (.D(_03378_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [479]),
    .QN(_28274_));
 DFF_X1 _61707_ (.D(_03380_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [480]),
    .QN(_28275_));
 DFF_X1 _61708_ (.D(_03381_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [481]),
    .QN(_28276_));
 DFF_X1 _61709_ (.D(_03382_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [482]),
    .QN(_28277_));
 DFF_X1 _61710_ (.D(_03383_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [483]),
    .QN(_28278_));
 DFF_X1 _61711_ (.D(_03384_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [484]),
    .QN(_28279_));
 DFF_X1 _61712_ (.D(_03385_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [485]),
    .QN(_28280_));
 DFF_X1 _61713_ (.D(_03386_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [486]),
    .QN(_28281_));
 DFF_X1 _61714_ (.D(_03387_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [487]),
    .QN(_28282_));
 DFF_X1 _61715_ (.D(_03388_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [488]),
    .QN(_28283_));
 DFF_X1 _61716_ (.D(_03389_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [489]),
    .QN(_28284_));
 DFF_X1 _61717_ (.D(_03391_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [490]),
    .QN(_28285_));
 DFF_X1 _61718_ (.D(_03392_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [491]),
    .QN(_28286_));
 DFF_X1 _61719_ (.D(_03393_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [492]),
    .QN(_28287_));
 DFF_X1 _61720_ (.D(_03394_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [493]),
    .QN(_28288_));
 DFF_X1 _61721_ (.D(_03395_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [494]),
    .QN(_28289_));
 DFF_X1 _61722_ (.D(_03396_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [495]),
    .QN(_28290_));
 DFF_X1 _61723_ (.D(_03397_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [496]),
    .QN(_28291_));
 DFF_X1 _61724_ (.D(_03398_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [497]),
    .QN(_28292_));
 DFF_X1 _61725_ (.D(_03399_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [498]),
    .QN(_28293_));
 DFF_X1 _61726_ (.D(_03400_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [499]),
    .QN(_28294_));
 DFF_X1 _61727_ (.D(_03403_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [500]),
    .QN(_28295_));
 DFF_X1 _61728_ (.D(_03404_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [501]),
    .QN(_28296_));
 DFF_X1 _61729_ (.D(_03405_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [502]),
    .QN(_28297_));
 DFF_X1 _61730_ (.D(_03406_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [503]),
    .QN(_28298_));
 DFF_X1 _61731_ (.D(_03407_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [504]),
    .QN(_28299_));
 DFF_X1 _61732_ (.D(_03408_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [505]),
    .QN(_28300_));
 DFF_X1 _61733_ (.D(_03409_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [506]),
    .QN(_28301_));
 DFF_X1 _61734_ (.D(_03410_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [507]),
    .QN(_28302_));
 DFF_X1 _61735_ (.D(_03411_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [508]),
    .QN(_28303_));
 DFF_X1 _61736_ (.D(_03412_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [509]),
    .QN(_28304_));
 DFF_X1 _61737_ (.D(_03414_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [510]),
    .QN(_28305_));
 DFF_X1 _61738_ (.D(_03415_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [511]),
    .QN(_28306_));
 DFF_X1 _61739_ (.D(_03416_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [512]),
    .QN(_28307_));
 DFF_X1 _61740_ (.D(_03417_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [513]),
    .QN(_28308_));
 DFF_X1 _61741_ (.D(_03418_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [514]),
    .QN(_28309_));
 DFF_X1 _61742_ (.D(_03419_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [515]),
    .QN(_28310_));
 DFF_X1 _61743_ (.D(_03420_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [516]),
    .QN(_28311_));
 DFF_X1 _61744_ (.D(_03421_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [517]),
    .QN(_28312_));
 DFF_X1 _61745_ (.D(_03422_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [518]),
    .QN(_28313_));
 DFF_X1 _61746_ (.D(_03423_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [519]),
    .QN(_28314_));
 DFF_X1 _61747_ (.D(_03425_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [520]),
    .QN(_28315_));
 DFF_X1 _61748_ (.D(_03426_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [521]),
    .QN(_28316_));
 DFF_X1 _61749_ (.D(_03427_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [522]),
    .QN(_28317_));
 DFF_X1 _61750_ (.D(_03428_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [523]),
    .QN(_28318_));
 DFF_X1 _61751_ (.D(_03429_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [524]),
    .QN(_28319_));
 DFF_X1 _61752_ (.D(_03430_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [525]),
    .QN(_28320_));
 DFF_X1 _61753_ (.D(_03431_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [526]),
    .QN(_28321_));
 DFF_X1 _61754_ (.D(_03432_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [527]),
    .QN(_28322_));
 DFF_X1 _61755_ (.D(_03433_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [528]),
    .QN(_28323_));
 DFF_X1 _61756_ (.D(_03434_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [529]),
    .QN(_28324_));
 DFF_X1 _61757_ (.D(_03436_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [530]),
    .QN(_28325_));
 DFF_X1 _61758_ (.D(_03437_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [531]),
    .QN(_28326_));
 DFF_X1 _61759_ (.D(_03438_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [532]),
    .QN(_28327_));
 DFF_X1 _61760_ (.D(_03439_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [533]),
    .QN(_28328_));
 DFF_X1 _61761_ (.D(_03440_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [534]),
    .QN(_28329_));
 DFF_X1 _61762_ (.D(_03441_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [535]),
    .QN(_28330_));
 DFF_X1 _61763_ (.D(_03442_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [536]),
    .QN(_28331_));
 DFF_X1 _61764_ (.D(_03443_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [537]),
    .QN(_28332_));
 DFF_X1 _61765_ (.D(_03444_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [538]),
    .QN(_28333_));
 DFF_X1 _61766_ (.D(_03445_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [539]),
    .QN(_28334_));
 DFF_X1 _61767_ (.D(_03447_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [540]),
    .QN(_28335_));
 DFF_X1 _61768_ (.D(_03448_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [541]),
    .QN(_28336_));
 DFF_X1 _61769_ (.D(_03449_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [542]),
    .QN(_28337_));
 DFF_X1 _61770_ (.D(_03450_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [543]),
    .QN(_28338_));
 DFF_X1 _61771_ (.D(_03451_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [544]),
    .QN(_28339_));
 DFF_X1 _61772_ (.D(_03452_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [545]),
    .QN(_28340_));
 DFF_X1 _61773_ (.D(_03453_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [546]),
    .QN(_28341_));
 DFF_X1 _61774_ (.D(_03454_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [547]),
    .QN(_28342_));
 DFF_X1 _61775_ (.D(_03455_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [548]),
    .QN(_28343_));
 DFF_X1 _61776_ (.D(_03456_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [549]),
    .QN(_28344_));
 DFF_X1 _61777_ (.D(_03458_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [550]),
    .QN(_28345_));
 DFF_X1 _61778_ (.D(_03459_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [551]),
    .QN(_28346_));
 DFF_X1 _61779_ (.D(_03460_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [552]),
    .QN(_28347_));
 DFF_X1 _61780_ (.D(_03461_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [553]),
    .QN(_28348_));
 DFF_X1 _61781_ (.D(_03462_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [554]),
    .QN(_28349_));
 DFF_X1 _61782_ (.D(_03463_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [555]),
    .QN(_28350_));
 DFF_X1 _61783_ (.D(_03464_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [556]),
    .QN(_28351_));
 DFF_X1 _61784_ (.D(_03465_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [557]),
    .QN(_28352_));
 DFF_X1 _61785_ (.D(_03466_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [558]),
    .QN(_28353_));
 DFF_X1 _61786_ (.D(_03467_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [559]),
    .QN(_28354_));
 DFF_X1 _61787_ (.D(_03469_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [560]),
    .QN(_28355_));
 DFF_X1 _61788_ (.D(_03470_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [561]),
    .QN(_28356_));
 DFF_X1 _61789_ (.D(_03471_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [562]),
    .QN(_28357_));
 DFF_X1 _61790_ (.D(_03472_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [563]),
    .QN(_28358_));
 DFF_X1 _61791_ (.D(_03473_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [564]),
    .QN(_28359_));
 DFF_X1 _61792_ (.D(_03474_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [565]),
    .QN(_28360_));
 DFF_X1 _61793_ (.D(_03475_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [566]),
    .QN(_28361_));
 DFF_X1 _61794_ (.D(_03476_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [567]),
    .QN(_28362_));
 DFF_X1 _61795_ (.D(_03477_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [568]),
    .QN(_28363_));
 DFF_X1 _61796_ (.D(_03478_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [569]),
    .QN(_28364_));
 DFF_X1 _61797_ (.D(_03480_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [570]),
    .QN(_28365_));
 DFF_X1 _61798_ (.D(_03481_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [571]),
    .QN(_28366_));
 DFF_X1 _61799_ (.D(_03482_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [572]),
    .QN(_28367_));
 DFF_X1 _61800_ (.D(_03483_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [573]),
    .QN(_28368_));
 DFF_X1 _61801_ (.D(_03484_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [574]),
    .QN(_28369_));
 DFF_X1 _61802_ (.D(_03485_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [575]),
    .QN(_28370_));
 DFF_X1 _61803_ (.D(_03486_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [576]),
    .QN(_28371_));
 DFF_X1 _61804_ (.D(_03487_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [577]),
    .QN(_28372_));
 DFF_X1 _61805_ (.D(_03488_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [578]),
    .QN(_28373_));
 DFF_X1 _61806_ (.D(_03489_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [579]),
    .QN(_28374_));
 DFF_X1 _61807_ (.D(_03491_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [580]),
    .QN(_28375_));
 DFF_X1 _61808_ (.D(_03492_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [581]),
    .QN(_28376_));
 DFF_X1 _61809_ (.D(_03493_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [582]),
    .QN(_28377_));
 DFF_X1 _61810_ (.D(_03494_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [583]),
    .QN(_28378_));
 DFF_X1 _61811_ (.D(_03495_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [584]),
    .QN(_28379_));
 DFF_X1 _61812_ (.D(_03496_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [585]),
    .QN(_28380_));
 DFF_X1 _61813_ (.D(_03497_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [586]),
    .QN(_28381_));
 DFF_X1 _61814_ (.D(_03498_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [587]),
    .QN(_28382_));
 DFF_X1 _61815_ (.D(_03499_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [588]),
    .QN(_28383_));
 DFF_X1 _61816_ (.D(_03500_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [589]),
    .QN(_28384_));
 DFF_X1 _61817_ (.D(_03502_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [590]),
    .QN(_28385_));
 DFF_X1 _61818_ (.D(_03503_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [591]),
    .QN(_28386_));
 DFF_X1 _61819_ (.D(_03504_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [592]),
    .QN(_28387_));
 DFF_X1 _61820_ (.D(_03505_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [593]),
    .QN(_28388_));
 DFF_X1 _61821_ (.D(_03506_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [594]),
    .QN(_28389_));
 DFF_X1 _61822_ (.D(_03507_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [595]),
    .QN(_28390_));
 DFF_X1 _61823_ (.D(_03508_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [596]),
    .QN(_28391_));
 DFF_X1 _61824_ (.D(_03509_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [597]),
    .QN(_28392_));
 DFF_X1 _61825_ (.D(_03510_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [598]),
    .QN(_28393_));
 DFF_X1 _61826_ (.D(_03511_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [599]),
    .QN(_28394_));
 DFF_X1 _61827_ (.D(_03514_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [600]),
    .QN(_28395_));
 DFF_X1 _61828_ (.D(_03515_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [601]),
    .QN(_28396_));
 DFF_X1 _61829_ (.D(_03516_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [602]),
    .QN(_28397_));
 DFF_X1 _61830_ (.D(_03517_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [603]),
    .QN(_28398_));
 DFF_X1 _61831_ (.D(_03518_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [604]),
    .QN(_28399_));
 DFF_X1 _61832_ (.D(_03519_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [605]),
    .QN(_28400_));
 DFF_X1 _61833_ (.D(_03520_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [606]),
    .QN(_28401_));
 DFF_X1 _61834_ (.D(_03521_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [607]),
    .QN(_28402_));
 DFF_X1 _61835_ (.D(_03522_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [608]),
    .QN(_28403_));
 DFF_X1 _61836_ (.D(_03523_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [609]),
    .QN(_28404_));
 DFF_X1 _61837_ (.D(_03525_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [610]),
    .QN(_28405_));
 DFF_X1 _61838_ (.D(_03526_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [611]),
    .QN(_28406_));
 DFF_X1 _61839_ (.D(_03527_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [612]),
    .QN(_28407_));
 DFF_X1 _61840_ (.D(_03528_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [613]),
    .QN(_28408_));
 DFF_X1 _61841_ (.D(_03529_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [614]),
    .QN(_28409_));
 DFF_X1 _61842_ (.D(_03530_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [615]),
    .QN(_28410_));
 DFF_X1 _61843_ (.D(_03531_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [616]),
    .QN(_28411_));
 DFF_X1 _61844_ (.D(_03532_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [617]),
    .QN(_28412_));
 DFF_X1 _61845_ (.D(_03533_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [618]),
    .QN(_28413_));
 DFF_X1 _61846_ (.D(_03534_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [619]),
    .QN(_28414_));
 DFF_X1 _61847_ (.D(_03536_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [620]),
    .QN(_28415_));
 DFF_X1 _61848_ (.D(_03537_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [621]),
    .QN(_28416_));
 DFF_X1 _61849_ (.D(_03538_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [622]),
    .QN(_28417_));
 DFF_X1 _61850_ (.D(_03539_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [623]),
    .QN(_28418_));
 DFF_X1 _61851_ (.D(_03540_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [624]),
    .QN(_28419_));
 DFF_X1 _61852_ (.D(_03541_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [625]),
    .QN(_28420_));
 DFF_X1 _61853_ (.D(_03542_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [626]),
    .QN(_28421_));
 DFF_X1 _61854_ (.D(_03543_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [627]),
    .QN(_28422_));
 DFF_X1 _61855_ (.D(_03544_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [628]),
    .QN(_28423_));
 DFF_X1 _61856_ (.D(_03545_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [629]),
    .QN(_28424_));
 DFF_X1 _61857_ (.D(_03547_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [630]),
    .QN(_28425_));
 DFF_X1 _61858_ (.D(_03548_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [631]),
    .QN(_28426_));
 DFF_X1 _61859_ (.D(_03549_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [632]),
    .QN(_28427_));
 DFF_X1 _61860_ (.D(_03550_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [633]),
    .QN(_28428_));
 DFF_X1 _61861_ (.D(_03551_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [634]),
    .QN(_28429_));
 DFF_X1 _61862_ (.D(_03552_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [635]),
    .QN(_28430_));
 DFF_X1 _61863_ (.D(_03553_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [636]),
    .QN(_28431_));
 DFF_X1 _61864_ (.D(_03554_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [637]),
    .QN(_28432_));
 DFF_X1 _61865_ (.D(_03555_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [638]),
    .QN(_28433_));
 DFF_X1 _61866_ (.D(_03556_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [639]),
    .QN(_28434_));
 DFF_X1 _61867_ (.D(_03558_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [640]),
    .QN(_28435_));
 DFF_X1 _61868_ (.D(_03559_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [641]),
    .QN(_28436_));
 DFF_X1 _61869_ (.D(_03560_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [642]),
    .QN(_28437_));
 DFF_X1 _61870_ (.D(_03561_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [643]),
    .QN(_28438_));
 DFF_X1 _61871_ (.D(_03562_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [644]),
    .QN(_28439_));
 DFF_X1 _61872_ (.D(_03563_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [645]),
    .QN(_28440_));
 DFF_X1 _61873_ (.D(_03564_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [646]),
    .QN(_28441_));
 DFF_X1 _61874_ (.D(_03565_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [647]),
    .QN(_28442_));
 DFF_X1 _61875_ (.D(_03566_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [648]),
    .QN(_28443_));
 DFF_X1 _61876_ (.D(_03567_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [649]),
    .QN(_28444_));
 DFF_X1 _61877_ (.D(_03569_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [650]),
    .QN(_28445_));
 DFF_X1 _61878_ (.D(_03570_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [651]),
    .QN(_28446_));
 DFF_X1 _61879_ (.D(_03571_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [652]),
    .QN(_28447_));
 DFF_X1 _61880_ (.D(_03572_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [653]),
    .QN(_28448_));
 DFF_X1 _61881_ (.D(_03573_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [654]),
    .QN(_28449_));
 DFF_X1 _61882_ (.D(_03574_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [655]),
    .QN(_28450_));
 DFF_X1 _61883_ (.D(_03575_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [656]),
    .QN(_28451_));
 DFF_X1 _61884_ (.D(_03576_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [657]),
    .QN(_28452_));
 DFF_X1 _61885_ (.D(_03577_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [658]),
    .QN(_28453_));
 DFF_X1 _61886_ (.D(_03578_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [659]),
    .QN(_28454_));
 DFF_X1 _61887_ (.D(_03580_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [660]),
    .QN(_28455_));
 DFF_X1 _61888_ (.D(_03581_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [661]),
    .QN(_28456_));
 DFF_X1 _61889_ (.D(_03582_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [662]),
    .QN(_28457_));
 DFF_X1 _61890_ (.D(_03583_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [663]),
    .QN(_28458_));
 DFF_X1 _61891_ (.D(_03584_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [664]),
    .QN(_28459_));
 DFF_X1 _61892_ (.D(_03585_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [665]),
    .QN(_28460_));
 DFF_X1 _61893_ (.D(_03586_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [666]),
    .QN(_28461_));
 DFF_X1 _61894_ (.D(_03587_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [667]),
    .QN(_28462_));
 DFF_X1 _61895_ (.D(_03588_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [668]),
    .QN(_28463_));
 DFF_X1 _61896_ (.D(_03589_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [669]),
    .QN(_28464_));
 DFF_X1 _61897_ (.D(_03591_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [670]),
    .QN(_28465_));
 DFF_X1 _61898_ (.D(_03592_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [671]),
    .QN(_28466_));
 DFF_X1 _61899_ (.D(_03593_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [672]),
    .QN(_28467_));
 DFF_X1 _61900_ (.D(_03594_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [673]),
    .QN(_28468_));
 DFF_X1 _61901_ (.D(_03595_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [674]),
    .QN(_28469_));
 DFF_X1 _61902_ (.D(_03596_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [675]),
    .QN(_28470_));
 DFF_X1 _61903_ (.D(_03597_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [676]),
    .QN(_28471_));
 DFF_X1 _61904_ (.D(_03598_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [677]),
    .QN(_28472_));
 DFF_X1 _61905_ (.D(_03599_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [678]),
    .QN(_28473_));
 DFF_X1 _61906_ (.D(_03600_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [679]),
    .QN(_28474_));
 DFF_X1 _61907_ (.D(_03602_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [680]),
    .QN(_28475_));
 DFF_X1 _61908_ (.D(_03603_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [681]),
    .QN(_28476_));
 DFF_X1 _61909_ (.D(_03604_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [682]),
    .QN(_28477_));
 DFF_X1 _61910_ (.D(_03605_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [683]),
    .QN(_28478_));
 DFF_X1 _61911_ (.D(_03606_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [684]),
    .QN(_28479_));
 DFF_X1 _61912_ (.D(_03607_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [685]),
    .QN(_28480_));
 DFF_X1 _61913_ (.D(_03608_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [686]),
    .QN(_28481_));
 DFF_X1 _61914_ (.D(_03609_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [687]),
    .QN(_28482_));
 DFF_X1 _61915_ (.D(_03610_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [688]),
    .QN(_28483_));
 DFF_X1 _61916_ (.D(_03611_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [689]),
    .QN(_28484_));
 DFF_X1 _61917_ (.D(_03613_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [690]),
    .QN(_28485_));
 DFF_X1 _61918_ (.D(_03614_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [691]),
    .QN(_28486_));
 DFF_X1 _61919_ (.D(_03615_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [692]),
    .QN(_28487_));
 DFF_X1 _61920_ (.D(_03616_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [693]),
    .QN(_28488_));
 DFF_X1 _61921_ (.D(_03617_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [694]),
    .QN(_28489_));
 DFF_X1 _61922_ (.D(_03618_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [695]),
    .QN(_28490_));
 DFF_X1 _61923_ (.D(_03619_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [696]),
    .QN(_28491_));
 DFF_X1 _61924_ (.D(_03620_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [697]),
    .QN(_28492_));
 DFF_X1 _61925_ (.D(_03621_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [698]),
    .QN(_28493_));
 DFF_X1 _61926_ (.D(_03622_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [699]),
    .QN(_28494_));
 DFF_X1 _61927_ (.D(_03625_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [700]),
    .QN(_28495_));
 DFF_X1 _61928_ (.D(_03626_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [701]),
    .QN(_28496_));
 DFF_X1 _61929_ (.D(_03627_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [702]),
    .QN(_28497_));
 DFF_X1 _61930_ (.D(_03628_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [703]),
    .QN(_28498_));
 DFF_X1 _61931_ (.D(_03629_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [704]),
    .QN(_28499_));
 DFF_X1 _61932_ (.D(_03630_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [705]),
    .QN(_28500_));
 DFF_X1 _61933_ (.D(_03631_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [706]),
    .QN(_28501_));
 DFF_X1 _61934_ (.D(_03632_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [707]),
    .QN(_28502_));
 DFF_X1 _61935_ (.D(_03633_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [708]),
    .QN(_28503_));
 DFF_X1 _61936_ (.D(_03634_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [709]),
    .QN(_28504_));
 DFF_X1 _61937_ (.D(_03636_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [710]),
    .QN(_28505_));
 DFF_X1 _61938_ (.D(_03637_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [711]),
    .QN(_28506_));
 DFF_X1 _61939_ (.D(_03638_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [712]),
    .QN(_28507_));
 DFF_X1 _61940_ (.D(_03639_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [713]),
    .QN(_28508_));
 DFF_X1 _61941_ (.D(_03640_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [714]),
    .QN(_28509_));
 DFF_X1 _61942_ (.D(_03641_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [715]),
    .QN(_28510_));
 DFF_X1 _61943_ (.D(_03642_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [716]),
    .QN(_28511_));
 DFF_X1 _61944_ (.D(_03643_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [717]),
    .QN(_28512_));
 DFF_X1 _61945_ (.D(_03644_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [718]),
    .QN(_28513_));
 DFF_X1 _61946_ (.D(_03645_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [719]),
    .QN(_28514_));
 DFF_X1 _61947_ (.D(_03647_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [720]),
    .QN(_28515_));
 DFF_X1 _61948_ (.D(_03648_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [721]),
    .QN(_28516_));
 DFF_X1 _61949_ (.D(_03649_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [722]),
    .QN(_28517_));
 DFF_X1 _61950_ (.D(_03650_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [723]),
    .QN(_28518_));
 DFF_X1 _61951_ (.D(_03651_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [724]),
    .QN(_28519_));
 DFF_X1 _61952_ (.D(_03652_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [725]),
    .QN(_28520_));
 DFF_X1 _61953_ (.D(_03653_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [726]),
    .QN(_28521_));
 DFF_X1 _61954_ (.D(_03654_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [727]),
    .QN(_28522_));
 DFF_X1 _61955_ (.D(_03655_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [728]),
    .QN(_28523_));
 DFF_X1 _61956_ (.D(_03656_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [729]),
    .QN(_28524_));
 DFF_X1 _61957_ (.D(_03658_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [730]),
    .QN(_28525_));
 DFF_X1 _61958_ (.D(_03659_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [731]),
    .QN(_28526_));
 DFF_X1 _61959_ (.D(_03660_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [732]),
    .QN(_28527_));
 DFF_X1 _61960_ (.D(_03661_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [733]),
    .QN(_28528_));
 DFF_X1 _61961_ (.D(_03662_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [734]),
    .QN(_28529_));
 DFF_X1 _61962_ (.D(_03663_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [735]),
    .QN(_28530_));
 DFF_X1 _61963_ (.D(_03664_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [736]),
    .QN(_28531_));
 DFF_X1 _61964_ (.D(_03665_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [737]),
    .QN(_28532_));
 DFF_X1 _61965_ (.D(_03666_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [738]),
    .QN(_28533_));
 DFF_X1 _61966_ (.D(_03667_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [739]),
    .QN(_28534_));
 DFF_X1 _61967_ (.D(_03669_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [740]),
    .QN(_28535_));
 DFF_X1 _61968_ (.D(_03670_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [741]),
    .QN(_28536_));
 DFF_X1 _61969_ (.D(_03671_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [742]),
    .QN(_28537_));
 DFF_X1 _61970_ (.D(_03672_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [743]),
    .QN(_28538_));
 DFF_X1 _61971_ (.D(_03673_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [744]),
    .QN(_28539_));
 DFF_X1 _61972_ (.D(_03674_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [745]),
    .QN(_28540_));
 DFF_X1 _61973_ (.D(_03675_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [746]),
    .QN(_28541_));
 DFF_X1 _61974_ (.D(_03676_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [747]),
    .QN(_28542_));
 DFF_X1 _61975_ (.D(_03677_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [748]),
    .QN(_28543_));
 DFF_X1 _61976_ (.D(_03678_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [749]),
    .QN(_28544_));
 DFF_X1 _61977_ (.D(_03680_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [750]),
    .QN(_28545_));
 DFF_X1 _61978_ (.D(_03681_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [751]),
    .QN(_28546_));
 DFF_X1 _61979_ (.D(_03682_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [752]),
    .QN(_28547_));
 DFF_X1 _61980_ (.D(_03683_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [753]),
    .QN(_28548_));
 DFF_X1 _61981_ (.D(_03684_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [754]),
    .QN(_28549_));
 DFF_X1 _61982_ (.D(_03685_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [755]),
    .QN(_28550_));
 DFF_X1 _61983_ (.D(_03686_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [756]),
    .QN(_28551_));
 DFF_X1 _61984_ (.D(_03687_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [757]),
    .QN(_28552_));
 DFF_X1 _61985_ (.D(_03688_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [758]),
    .QN(_28553_));
 DFF_X1 _61986_ (.D(_03689_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [759]),
    .QN(_28554_));
 DFF_X1 _61987_ (.D(_03691_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [760]),
    .QN(_28555_));
 DFF_X1 _61988_ (.D(_03692_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [761]),
    .QN(_28556_));
 DFF_X1 _61989_ (.D(_03693_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [762]),
    .QN(_28557_));
 DFF_X1 _61990_ (.D(_03694_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [763]),
    .QN(_28558_));
 DFF_X1 _61991_ (.D(_03695_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [764]),
    .QN(_28559_));
 DFF_X1 _61992_ (.D(_03696_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [765]),
    .QN(_28560_));
 DFF_X1 _61993_ (.D(_03697_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [766]),
    .QN(_28561_));
 DFF_X1 _61994_ (.D(_03698_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [767]),
    .QN(_28562_));
 DFF_X1 _61995_ (.D(_03699_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [768]),
    .QN(_28563_));
 DFF_X1 _61996_ (.D(_03700_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [769]),
    .QN(_28564_));
 DFF_X1 _61997_ (.D(_03702_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [770]),
    .QN(_28565_));
 DFF_X1 _61998_ (.D(_03703_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [771]),
    .QN(_28566_));
 DFF_X1 _61999_ (.D(_03704_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [772]),
    .QN(_28567_));
 DFF_X1 _62000_ (.D(_03705_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [773]),
    .QN(_28568_));
 DFF_X1 _62001_ (.D(_03706_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [774]),
    .QN(_28569_));
 DFF_X1 _62002_ (.D(_03707_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [775]),
    .QN(_28570_));
 DFF_X1 _62003_ (.D(_03708_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [776]),
    .QN(_28571_));
 DFF_X1 _62004_ (.D(_03709_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [777]),
    .QN(_28572_));
 DFF_X1 _62005_ (.D(_03710_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [778]),
    .QN(_28573_));
 DFF_X1 _62006_ (.D(_03711_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [779]),
    .QN(_28574_));
 DFF_X1 _62007_ (.D(_03713_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [780]),
    .QN(_28575_));
 DFF_X1 _62008_ (.D(_03714_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [781]),
    .QN(_28576_));
 DFF_X1 _62009_ (.D(_03715_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [782]),
    .QN(_28577_));
 DFF_X1 _62010_ (.D(_03716_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [783]),
    .QN(_28578_));
 DFF_X1 _62011_ (.D(_03717_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [784]),
    .QN(_28579_));
 DFF_X1 _62012_ (.D(_03718_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [785]),
    .QN(_28580_));
 DFF_X1 _62013_ (.D(_03719_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [786]),
    .QN(_28581_));
 DFF_X1 _62014_ (.D(_03720_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [787]),
    .QN(_28582_));
 DFF_X1 _62015_ (.D(_03721_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [788]),
    .QN(_28583_));
 DFF_X1 _62016_ (.D(_03722_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [789]),
    .QN(_28584_));
 DFF_X1 _62017_ (.D(_03724_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [790]),
    .QN(_28585_));
 DFF_X1 _62018_ (.D(_03725_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [791]),
    .QN(_28586_));
 DFF_X1 _62019_ (.D(_03726_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [792]),
    .QN(_28587_));
 DFF_X1 _62020_ (.D(_03727_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [793]),
    .QN(_28588_));
 DFF_X1 _62021_ (.D(_03728_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [794]),
    .QN(_28589_));
 DFF_X1 _62022_ (.D(_03729_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [795]),
    .QN(_28590_));
 DFF_X1 _62023_ (.D(_03730_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [796]),
    .QN(_28591_));
 DFF_X1 _62024_ (.D(_03731_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [797]),
    .QN(_28592_));
 DFF_X1 _62025_ (.D(_03732_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [798]),
    .QN(_28593_));
 DFF_X1 _62026_ (.D(_03733_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [799]),
    .QN(_28594_));
 DFF_X1 _62027_ (.D(_03736_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [800]),
    .QN(_28595_));
 DFF_X1 _62028_ (.D(_03737_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [801]),
    .QN(_28596_));
 DFF_X1 _62029_ (.D(_03738_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [802]),
    .QN(_28597_));
 DFF_X1 _62030_ (.D(_03739_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [803]),
    .QN(_28598_));
 DFF_X1 _62031_ (.D(_03740_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [804]),
    .QN(_28599_));
 DFF_X1 _62032_ (.D(_03741_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [805]),
    .QN(_28600_));
 DFF_X1 _62033_ (.D(_03742_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [806]),
    .QN(_28601_));
 DFF_X1 _62034_ (.D(_03743_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [807]),
    .QN(_28602_));
 DFF_X1 _62035_ (.D(_03744_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [808]),
    .QN(_28603_));
 DFF_X1 _62036_ (.D(_03745_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [809]),
    .QN(_28604_));
 DFF_X1 _62037_ (.D(_03747_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [810]),
    .QN(_28605_));
 DFF_X1 _62038_ (.D(_03748_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [811]),
    .QN(_28606_));
 DFF_X1 _62039_ (.D(_03749_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [812]),
    .QN(_28607_));
 DFF_X1 _62040_ (.D(_03750_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [813]),
    .QN(_28608_));
 DFF_X1 _62041_ (.D(_03751_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [814]),
    .QN(_28609_));
 DFF_X1 _62042_ (.D(_03752_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [815]),
    .QN(_28610_));
 DFF_X1 _62043_ (.D(_03753_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [816]),
    .QN(_28611_));
 DFF_X1 _62044_ (.D(_03754_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [817]),
    .QN(_28612_));
 DFF_X1 _62045_ (.D(_03755_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [818]),
    .QN(_28613_));
 DFF_X1 _62046_ (.D(_03756_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [819]),
    .QN(_28614_));
 DFF_X1 _62047_ (.D(_03758_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [820]),
    .QN(_28615_));
 DFF_X1 _62048_ (.D(_03759_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [821]),
    .QN(_28616_));
 DFF_X1 _62049_ (.D(_03760_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [822]),
    .QN(_28617_));
 DFF_X1 _62050_ (.D(_03761_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [823]),
    .QN(_28618_));
 DFF_X1 _62051_ (.D(_03762_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [824]),
    .QN(_28619_));
 DFF_X1 _62052_ (.D(_03763_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [825]),
    .QN(_28620_));
 DFF_X1 _62053_ (.D(_03764_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [826]),
    .QN(_28621_));
 DFF_X1 _62054_ (.D(_03765_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [827]),
    .QN(_28622_));
 DFF_X1 _62055_ (.D(_03766_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [828]),
    .QN(_28623_));
 DFF_X1 _62056_ (.D(_03767_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [829]),
    .QN(_28624_));
 DFF_X1 _62057_ (.D(_03769_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [830]),
    .QN(_28625_));
 DFF_X1 _62058_ (.D(_03770_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [831]),
    .QN(_28626_));
 DFF_X1 _62059_ (.D(_03771_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [832]),
    .QN(_28627_));
 DFF_X1 _62060_ (.D(_03772_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [833]),
    .QN(_28628_));
 DFF_X1 _62061_ (.D(_03773_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [834]),
    .QN(_28629_));
 DFF_X1 _62062_ (.D(_03774_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [835]),
    .QN(_28630_));
 DFF_X1 _62063_ (.D(_03775_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [836]),
    .QN(_28631_));
 DFF_X1 _62064_ (.D(_03776_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [837]),
    .QN(_28632_));
 DFF_X1 _62065_ (.D(_03777_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [838]),
    .QN(_28633_));
 DFF_X1 _62066_ (.D(_03778_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [839]),
    .QN(_28634_));
 DFF_X1 _62067_ (.D(_03780_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [840]),
    .QN(_28635_));
 DFF_X1 _62068_ (.D(_03781_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [841]),
    .QN(_28636_));
 DFF_X1 _62069_ (.D(_03782_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [842]),
    .QN(_28637_));
 DFF_X1 _62070_ (.D(_03783_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [843]),
    .QN(_28638_));
 DFF_X1 _62071_ (.D(_03784_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [844]),
    .QN(_28639_));
 DFF_X1 _62072_ (.D(_03785_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [845]),
    .QN(_28640_));
 DFF_X1 _62073_ (.D(_03786_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [846]),
    .QN(_28641_));
 DFF_X1 _62074_ (.D(_03787_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [847]),
    .QN(_28642_));
 DFF_X1 _62075_ (.D(_03788_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [848]),
    .QN(_28643_));
 DFF_X1 _62076_ (.D(_03789_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [849]),
    .QN(_28644_));
 DFF_X1 _62077_ (.D(_03791_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [850]),
    .QN(_28645_));
 DFF_X1 _62078_ (.D(_03792_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [851]),
    .QN(_28646_));
 DFF_X1 _62079_ (.D(_03793_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [852]),
    .QN(_28647_));
 DFF_X1 _62080_ (.D(_03794_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [853]),
    .QN(_28648_));
 DFF_X1 _62081_ (.D(_03795_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [854]),
    .QN(_28649_));
 DFF_X1 _62082_ (.D(_03796_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [855]),
    .QN(_28650_));
 DFF_X1 _62083_ (.D(_03797_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [856]),
    .QN(_28651_));
 DFF_X1 _62084_ (.D(_03798_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [857]),
    .QN(_28652_));
 DFF_X1 _62085_ (.D(_03799_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [858]),
    .QN(_28653_));
 DFF_X1 _62086_ (.D(_03800_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [859]),
    .QN(_28654_));
 DFF_X1 _62087_ (.D(_03802_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [860]),
    .QN(_28655_));
 DFF_X1 _62088_ (.D(_03803_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [861]),
    .QN(_28656_));
 DFF_X1 _62089_ (.D(_03804_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [862]),
    .QN(_28657_));
 DFF_X1 _62090_ (.D(_03805_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [863]),
    .QN(_28658_));
 DFF_X1 _62091_ (.D(_03806_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [864]),
    .QN(_28659_));
 DFF_X1 _62092_ (.D(_03807_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [865]),
    .QN(_28660_));
 DFF_X1 _62093_ (.D(_03808_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [866]),
    .QN(_28661_));
 DFF_X1 _62094_ (.D(_03809_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [867]),
    .QN(_28662_));
 DFF_X1 _62095_ (.D(_03810_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [868]),
    .QN(_28663_));
 DFF_X1 _62096_ (.D(_03811_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [869]),
    .QN(_28664_));
 DFF_X1 _62097_ (.D(_03813_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [870]),
    .QN(_28665_));
 DFF_X1 _62098_ (.D(_03814_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [871]),
    .QN(_28666_));
 DFF_X1 _62099_ (.D(_03815_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [872]),
    .QN(_28667_));
 DFF_X1 _62100_ (.D(_03816_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [873]),
    .QN(_28668_));
 DFF_X1 _62101_ (.D(_03817_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [874]),
    .QN(_28669_));
 DFF_X1 _62102_ (.D(_03818_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [875]),
    .QN(_28670_));
 DFF_X1 _62103_ (.D(_03819_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [876]),
    .QN(_28671_));
 DFF_X1 _62104_ (.D(_03820_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [877]),
    .QN(_28672_));
 DFF_X1 _62105_ (.D(_03821_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [878]),
    .QN(_28673_));
 DFF_X1 _62106_ (.D(_03822_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [879]),
    .QN(_28674_));
 DFF_X1 _62107_ (.D(_03824_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [880]),
    .QN(_28675_));
 DFF_X1 _62108_ (.D(_03825_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [881]),
    .QN(_28676_));
 DFF_X1 _62109_ (.D(_03826_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [882]),
    .QN(_28677_));
 DFF_X1 _62110_ (.D(_03827_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [883]),
    .QN(_28678_));
 DFF_X1 _62111_ (.D(_03828_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [884]),
    .QN(_28679_));
 DFF_X1 _62112_ (.D(_03829_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [885]),
    .QN(_28680_));
 DFF_X1 _62113_ (.D(_03830_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [886]),
    .QN(_28681_));
 DFF_X1 _62114_ (.D(_03831_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [887]),
    .QN(_28682_));
 DFF_X1 _62115_ (.D(_03832_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [888]),
    .QN(_28683_));
 DFF_X1 _62116_ (.D(_03833_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [889]),
    .QN(_28684_));
 DFF_X1 _62117_ (.D(_03835_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [890]),
    .QN(_28685_));
 DFF_X1 _62118_ (.D(_03836_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [891]),
    .QN(_28686_));
 DFF_X1 _62119_ (.D(_03837_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [892]),
    .QN(_28687_));
 DFF_X1 _62120_ (.D(_03838_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [893]),
    .QN(_28688_));
 DFF_X1 _62121_ (.D(_03839_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [894]),
    .QN(_28689_));
 DFF_X1 _62122_ (.D(_03840_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [895]),
    .QN(_28690_));
 DFF_X1 _62123_ (.D(_03841_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [896]),
    .QN(_28691_));
 DFF_X1 _62124_ (.D(_03842_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [897]),
    .QN(_28692_));
 DFF_X1 _62125_ (.D(_03843_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [898]),
    .QN(_28693_));
 DFF_X1 _62126_ (.D(_03844_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [899]),
    .QN(_28694_));
 DFF_X1 _62127_ (.D(_03847_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [900]),
    .QN(_28695_));
 DFF_X1 _62128_ (.D(_03848_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [901]),
    .QN(_28696_));
 DFF_X1 _62129_ (.D(_03849_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [902]),
    .QN(_28697_));
 DFF_X1 _62130_ (.D(_03850_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [903]),
    .QN(_28698_));
 DFF_X1 _62131_ (.D(_03851_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [904]),
    .QN(_28699_));
 DFF_X1 _62132_ (.D(_03852_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [905]),
    .QN(_28700_));
 DFF_X1 _62133_ (.D(_03853_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [906]),
    .QN(_28701_));
 DFF_X1 _62134_ (.D(_03854_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [907]),
    .QN(_28702_));
 DFF_X1 _62135_ (.D(_03855_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [908]),
    .QN(_28703_));
 DFF_X1 _62136_ (.D(_03856_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [909]),
    .QN(_28704_));
 DFF_X1 _62137_ (.D(_03858_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [910]),
    .QN(_28705_));
 DFF_X1 _62138_ (.D(_03859_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [911]),
    .QN(_28706_));
 DFF_X1 _62139_ (.D(_03860_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [912]),
    .QN(_28707_));
 DFF_X1 _62140_ (.D(_03861_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [913]),
    .QN(_28708_));
 DFF_X1 _62141_ (.D(_03862_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [914]),
    .QN(_28709_));
 DFF_X1 _62142_ (.D(_03863_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [915]),
    .QN(_28710_));
 DFF_X1 _62143_ (.D(_03864_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [916]),
    .QN(_28711_));
 DFF_X1 _62144_ (.D(_03865_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [917]),
    .QN(_28712_));
 DFF_X1 _62145_ (.D(_03866_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [918]),
    .QN(_28713_));
 DFF_X1 _62146_ (.D(_03867_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [919]),
    .QN(_28714_));
 DFF_X1 _62147_ (.D(_03869_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [920]),
    .QN(_28715_));
 DFF_X1 _62148_ (.D(_03870_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [921]),
    .QN(_28716_));
 DFF_X1 _62149_ (.D(_03871_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [922]),
    .QN(_28717_));
 DFF_X1 _62150_ (.D(_03872_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [923]),
    .QN(_28718_));
 DFF_X1 _62151_ (.D(_03873_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [924]),
    .QN(_28719_));
 DFF_X1 _62152_ (.D(_03874_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [925]),
    .QN(_28720_));
 DFF_X1 _62153_ (.D(_03875_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [926]),
    .QN(_28721_));
 DFF_X1 _62154_ (.D(_03876_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [927]),
    .QN(_28722_));
 DFF_X1 _62155_ (.D(_03877_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [928]),
    .QN(_28723_));
 DFF_X1 _62156_ (.D(_03878_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [929]),
    .QN(_28724_));
 DFF_X1 _62157_ (.D(_03880_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [930]),
    .QN(_28725_));
 DFF_X1 _62158_ (.D(_03881_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [931]),
    .QN(_28726_));
 DFF_X1 _62159_ (.D(_03882_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [932]),
    .QN(_28727_));
 DFF_X1 _62160_ (.D(_03883_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [933]),
    .QN(_28728_));
 DFF_X1 _62161_ (.D(_03884_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [934]),
    .QN(_28729_));
 DFF_X1 _62162_ (.D(_03885_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [935]),
    .QN(_28730_));
 DFF_X1 _62163_ (.D(_03886_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [936]),
    .QN(_28731_));
 DFF_X1 _62164_ (.D(_03887_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [937]),
    .QN(_28732_));
 DFF_X1 _62165_ (.D(_03888_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [938]),
    .QN(_28733_));
 DFF_X1 _62166_ (.D(_03889_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [939]),
    .QN(_28734_));
 DFF_X1 _62167_ (.D(_03891_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [940]),
    .QN(_28735_));
 DFF_X1 _62168_ (.D(_03892_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [941]),
    .QN(_28736_));
 DFF_X1 _62169_ (.D(_03893_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [942]),
    .QN(_28737_));
 DFF_X1 _62170_ (.D(_03894_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [943]),
    .QN(_28738_));
 DFF_X1 _62171_ (.D(_03895_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [944]),
    .QN(_28739_));
 DFF_X1 _62172_ (.D(_03896_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [945]),
    .QN(_28740_));
 DFF_X1 _62173_ (.D(_03897_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [946]),
    .QN(_28741_));
 DFF_X1 _62174_ (.D(_03898_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [947]),
    .QN(_28742_));
 DFF_X1 _62175_ (.D(_03899_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [948]),
    .QN(_28743_));
 DFF_X1 _62176_ (.D(_03900_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [949]),
    .QN(_28744_));
 DFF_X1 _62177_ (.D(_03902_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [950]),
    .QN(_28745_));
 DFF_X1 _62178_ (.D(_03903_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [951]),
    .QN(_28746_));
 DFF_X1 _62179_ (.D(_03904_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [952]),
    .QN(_28747_));
 DFF_X1 _62180_ (.D(_03905_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [953]),
    .QN(_28748_));
 DFF_X1 _62181_ (.D(_03906_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [954]),
    .QN(_28749_));
 DFF_X1 _62182_ (.D(_03907_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [955]),
    .QN(_28750_));
 DFF_X1 _62183_ (.D(_03908_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [956]),
    .QN(_28751_));
 DFF_X1 _62184_ (.D(_03909_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [957]),
    .QN(_28752_));
 DFF_X1 _62185_ (.D(_03910_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [958]),
    .QN(_28753_));
 DFF_X1 _62186_ (.D(_03911_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [959]),
    .QN(_28754_));
 DFF_X1 _62187_ (.D(_03913_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [960]),
    .QN(_28755_));
 DFF_X1 _62188_ (.D(_03914_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [961]),
    .QN(_28756_));
 DFF_X1 _62189_ (.D(_03915_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [962]),
    .QN(_28757_));
 DFF_X1 _62190_ (.D(_03916_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [963]),
    .QN(_28758_));
 DFF_X1 _62191_ (.D(_03917_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [964]),
    .QN(_28759_));
 DFF_X1 _62192_ (.D(_03918_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [965]),
    .QN(_28760_));
 DFF_X1 _62193_ (.D(_03919_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [966]),
    .QN(_28761_));
 DFF_X1 _62194_ (.D(_03920_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [967]),
    .QN(_28762_));
 DFF_X1 _62195_ (.D(_03921_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [968]),
    .QN(_28763_));
 DFF_X1 _62196_ (.D(_03922_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [969]),
    .QN(_28764_));
 DFF_X1 _62197_ (.D(_03924_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [970]),
    .QN(_28765_));
 DFF_X1 _62198_ (.D(_03925_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [971]),
    .QN(_28766_));
 DFF_X1 _62199_ (.D(_03926_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [972]),
    .QN(_28767_));
 DFF_X1 _62200_ (.D(_03927_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [973]),
    .QN(_28768_));
 DFF_X1 _62201_ (.D(_03928_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [974]),
    .QN(_28769_));
 DFF_X1 _62202_ (.D(_03929_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [975]),
    .QN(_28770_));
 DFF_X1 _62203_ (.D(_03930_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [976]),
    .QN(_28771_));
 DFF_X1 _62204_ (.D(_03931_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [977]),
    .QN(_28772_));
 DFF_X1 _62205_ (.D(_03932_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [978]),
    .QN(_28773_));
 DFF_X1 _62206_ (.D(_03933_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [979]),
    .QN(_28774_));
 DFF_X1 _62207_ (.D(_03935_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [980]),
    .QN(_28775_));
 DFF_X1 _62208_ (.D(_03936_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [981]),
    .QN(_28776_));
 DFF_X1 _62209_ (.D(_03937_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [982]),
    .QN(_28777_));
 DFF_X1 _62210_ (.D(_03938_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [983]),
    .QN(_28778_));
 DFF_X1 _62211_ (.D(_03939_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [984]),
    .QN(_28779_));
 DFF_X1 _62212_ (.D(_03940_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [985]),
    .QN(_28780_));
 DFF_X1 _62213_ (.D(_03941_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [986]),
    .QN(_28781_));
 DFF_X1 _62214_ (.D(_03942_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [987]),
    .QN(_28782_));
 DFF_X1 _62215_ (.D(_03943_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [988]),
    .QN(_28783_));
 DFF_X1 _62216_ (.D(_03944_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [989]),
    .QN(_28784_));
 DFF_X1 _62217_ (.D(_03946_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [990]),
    .QN(_28785_));
 DFF_X1 _62218_ (.D(_03947_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [991]),
    .QN(_28786_));
 DFF_X1 _62219_ (.D(_03948_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [992]),
    .QN(_28787_));
 DFF_X1 _62220_ (.D(_03949_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [993]),
    .QN(_28788_));
 DFF_X1 _62221_ (.D(_03950_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [994]),
    .QN(_28789_));
 DFF_X1 _62222_ (.D(_03951_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [995]),
    .QN(_28790_));
 DFF_X1 _62223_ (.D(_03952_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [996]),
    .QN(_28791_));
 DFF_X1 _62224_ (.D(_03953_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [997]),
    .QN(_28792_));
 DFF_X1 _62225_ (.D(_03954_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [998]),
    .QN(_28793_));
 DFF_X1 _62226_ (.D(_03955_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [999]),
    .QN(_28794_));
 DFF_X1 _62227_ (.D(_00823_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1000]),
    .QN(_28795_));
 DFF_X1 _62228_ (.D(_00824_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1001]),
    .QN(_28796_));
 DFF_X1 _62229_ (.D(_00825_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1002]),
    .QN(_28797_));
 DFF_X1 _62230_ (.D(_00826_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1003]),
    .QN(_28798_));
 DFF_X1 _62231_ (.D(_00827_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1004]),
    .QN(_28799_));
 DFF_X1 _62232_ (.D(_00828_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1005]),
    .QN(_28800_));
 DFF_X1 _62233_ (.D(_00829_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1006]),
    .QN(_28801_));
 DFF_X1 _62234_ (.D(_00830_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1007]),
    .QN(_28802_));
 DFF_X1 _62235_ (.D(_00831_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1008]),
    .QN(_28803_));
 DFF_X1 _62236_ (.D(_00832_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1009]),
    .QN(_28804_));
 DFF_X1 _62237_ (.D(_00834_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1010]),
    .QN(_28805_));
 DFF_X1 _62238_ (.D(_00835_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1011]),
    .QN(_28806_));
 DFF_X1 _62239_ (.D(_00836_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1012]),
    .QN(_28807_));
 DFF_X1 _62240_ (.D(_00837_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1013]),
    .QN(_28808_));
 DFF_X1 _62241_ (.D(_00838_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1014]),
    .QN(_28809_));
 DFF_X1 _62242_ (.D(_00839_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1015]),
    .QN(_28810_));
 DFF_X1 _62243_ (.D(_00840_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1016]),
    .QN(_28811_));
 DFF_X1 _62244_ (.D(_00841_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1017]),
    .QN(_28812_));
 DFF_X1 _62245_ (.D(_00842_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1018]),
    .QN(_28813_));
 DFF_X1 _62246_ (.D(_00843_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1019]),
    .QN(_28814_));
 DFF_X1 _62247_ (.D(_00845_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1020]),
    .QN(_28815_));
 DFF_X1 _62248_ (.D(_00846_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1021]),
    .QN(_28816_));
 DFF_X1 _62249_ (.D(_00847_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1022]),
    .QN(_28817_));
 DFF_X1 _62250_ (.D(_00848_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1023]),
    .QN(_28818_));
 DFF_X1 _62251_ (.D(_00849_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1024]),
    .QN(_28819_));
 DFF_X1 _62252_ (.D(_00850_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1025]),
    .QN(_28820_));
 DFF_X1 _62253_ (.D(_00851_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1026]),
    .QN(_28821_));
 DFF_X1 _62254_ (.D(_00852_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1027]),
    .QN(_28822_));
 DFF_X1 _62255_ (.D(_00853_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1028]),
    .QN(_28823_));
 DFF_X1 _62256_ (.D(_00854_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1029]),
    .QN(_28824_));
 DFF_X1 _62257_ (.D(_00856_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1030]),
    .QN(_28825_));
 DFF_X1 _62258_ (.D(_00857_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1031]),
    .QN(_28826_));
 DFF_X1 _62259_ (.D(_00858_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1032]),
    .QN(_28827_));
 DFF_X1 _62260_ (.D(_00859_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1033]),
    .QN(_28828_));
 DFF_X1 _62261_ (.D(_00860_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1034]),
    .QN(_28829_));
 DFF_X1 _62262_ (.D(_00861_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1035]),
    .QN(_28830_));
 DFF_X1 _62263_ (.D(_00862_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1036]),
    .QN(_28831_));
 DFF_X1 _62264_ (.D(_00863_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1037]),
    .QN(_28832_));
 DFF_X1 _62265_ (.D(_00864_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1038]),
    .QN(_28833_));
 DFF_X1 _62266_ (.D(_00865_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1039]),
    .QN(_28834_));
 DFF_X1 _62267_ (.D(_00867_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1040]),
    .QN(_28835_));
 DFF_X1 _62268_ (.D(_00868_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1041]),
    .QN(_28836_));
 DFF_X1 _62269_ (.D(_00869_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1042]),
    .QN(_28837_));
 DFF_X1 _62270_ (.D(_00870_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1043]),
    .QN(_28838_));
 DFF_X1 _62271_ (.D(_00871_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1044]),
    .QN(_28839_));
 DFF_X1 _62272_ (.D(_00872_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1045]),
    .QN(_28840_));
 DFF_X1 _62273_ (.D(_00873_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1046]),
    .QN(_28841_));
 DFF_X1 _62274_ (.D(_00874_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1047]),
    .QN(_28842_));
 DFF_X1 _62275_ (.D(_00875_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1048]),
    .QN(_28843_));
 DFF_X1 _62276_ (.D(_00876_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1049]),
    .QN(_28844_));
 DFF_X1 _62277_ (.D(_00878_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1050]),
    .QN(_28845_));
 DFF_X1 _62278_ (.D(_00879_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1051]),
    .QN(_28846_));
 DFF_X1 _62279_ (.D(_00880_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1052]),
    .QN(_28847_));
 DFF_X1 _62280_ (.D(_00881_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1053]),
    .QN(_28848_));
 DFF_X1 _62281_ (.D(_00882_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1054]),
    .QN(_28849_));
 DFF_X1 _62282_ (.D(_00883_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1055]),
    .QN(_28850_));
 DFF_X1 _62283_ (.D(_00884_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1056]),
    .QN(_28851_));
 DFF_X1 _62284_ (.D(_00885_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1057]),
    .QN(_28852_));
 DFF_X1 _62285_ (.D(_00886_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1058]),
    .QN(_28853_));
 DFF_X1 _62286_ (.D(_00887_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1059]),
    .QN(_28854_));
 DFF_X1 _62287_ (.D(_00889_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1060]),
    .QN(_28855_));
 DFF_X1 _62288_ (.D(_00890_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1061]),
    .QN(_28856_));
 DFF_X1 _62289_ (.D(_00891_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1062]),
    .QN(_28857_));
 DFF_X1 _62290_ (.D(_00892_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1063]),
    .QN(_28858_));
 DFF_X1 _62291_ (.D(_00893_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1064]),
    .QN(_28859_));
 DFF_X1 _62292_ (.D(_00894_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1065]),
    .QN(_28860_));
 DFF_X1 _62293_ (.D(_00895_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1066]),
    .QN(_28861_));
 DFF_X1 _62294_ (.D(_00896_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1067]),
    .QN(_28862_));
 DFF_X1 _62295_ (.D(_00897_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1068]),
    .QN(_28863_));
 DFF_X1 _62296_ (.D(_00898_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1069]),
    .QN(_28864_));
 DFF_X1 _62297_ (.D(_00900_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1070]),
    .QN(_28865_));
 DFF_X1 _62298_ (.D(_00901_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1071]),
    .QN(_28866_));
 DFF_X1 _62299_ (.D(_00902_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1072]),
    .QN(_28867_));
 DFF_X1 _62300_ (.D(_00903_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1073]),
    .QN(_28868_));
 DFF_X1 _62301_ (.D(_00904_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1074]),
    .QN(_28869_));
 DFF_X1 _62302_ (.D(_00905_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1075]),
    .QN(_28870_));
 DFF_X1 _62303_ (.D(_00906_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1076]),
    .QN(_28871_));
 DFF_X1 _62304_ (.D(_00907_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1077]),
    .QN(_28872_));
 DFF_X1 _62305_ (.D(_00908_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1078]),
    .QN(_28873_));
 DFF_X1 _62306_ (.D(_00909_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1079]),
    .QN(_28874_));
 DFF_X1 _62307_ (.D(_00911_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1080]),
    .QN(_28875_));
 DFF_X1 _62308_ (.D(_00912_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1081]),
    .QN(_28876_));
 DFF_X1 _62309_ (.D(_00913_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1082]),
    .QN(_28877_));
 DFF_X1 _62310_ (.D(_00914_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1083]),
    .QN(_28878_));
 DFF_X1 _62311_ (.D(_00915_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1084]),
    .QN(_28879_));
 DFF_X1 _62312_ (.D(_00916_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1085]),
    .QN(_28880_));
 DFF_X1 _62313_ (.D(_00917_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1086]),
    .QN(_28881_));
 DFF_X1 _62314_ (.D(_00918_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1087]),
    .QN(_28882_));
 DFF_X1 _62315_ (.D(_00919_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1088]),
    .QN(_28883_));
 DFF_X1 _62316_ (.D(_00920_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1089]),
    .QN(_28884_));
 DFF_X1 _62317_ (.D(_00922_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1090]),
    .QN(_28885_));
 DFF_X1 _62318_ (.D(_00923_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1091]),
    .QN(_28886_));
 DFF_X1 _62319_ (.D(_00924_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1092]),
    .QN(_28887_));
 DFF_X1 _62320_ (.D(_00925_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1093]),
    .QN(_28888_));
 DFF_X1 _62321_ (.D(_00926_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1094]),
    .QN(_28889_));
 DFF_X1 _62322_ (.D(_00927_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1095]),
    .QN(_28890_));
 DFF_X1 _62323_ (.D(_00928_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1096]),
    .QN(_28891_));
 DFF_X1 _62324_ (.D(_00929_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1097]),
    .QN(_28892_));
 DFF_X1 _62325_ (.D(_00930_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1098]),
    .QN(_28893_));
 DFF_X1 _62326_ (.D(_00931_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1099]),
    .QN(_28894_));
 DFF_X1 _62327_ (.D(_00934_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1100]),
    .QN(_28895_));
 DFF_X1 _62328_ (.D(_00935_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1101]),
    .QN(_28896_));
 DFF_X1 _62329_ (.D(_00936_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1102]),
    .QN(_28897_));
 DFF_X1 _62330_ (.D(_00937_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1103]),
    .QN(_28898_));
 DFF_X1 _62331_ (.D(_00938_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1104]),
    .QN(_28899_));
 DFF_X1 _62332_ (.D(_00939_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1105]),
    .QN(_28900_));
 DFF_X1 _62333_ (.D(_00940_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1106]),
    .QN(_28901_));
 DFF_X1 _62334_ (.D(_00941_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1107]),
    .QN(_28902_));
 DFF_X1 _62335_ (.D(_00942_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1108]),
    .QN(_28903_));
 DFF_X1 _62336_ (.D(_00943_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1109]),
    .QN(_28904_));
 DFF_X1 _62337_ (.D(_00945_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1110]),
    .QN(_28905_));
 DFF_X1 _62338_ (.D(_00946_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1111]),
    .QN(_28906_));
 DFF_X1 _62339_ (.D(_00947_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1112]),
    .QN(_28907_));
 DFF_X1 _62340_ (.D(_00948_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1113]),
    .QN(_28908_));
 DFF_X1 _62341_ (.D(_00949_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1114]),
    .QN(_28909_));
 DFF_X1 _62342_ (.D(_00950_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1115]),
    .QN(_28910_));
 DFF_X1 _62343_ (.D(_00951_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1116]),
    .QN(_28911_));
 DFF_X1 _62344_ (.D(_00952_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1117]),
    .QN(_28912_));
 DFF_X1 _62345_ (.D(_00953_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1118]),
    .QN(_28913_));
 DFF_X1 _62346_ (.D(_00954_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1119]),
    .QN(_28914_));
 DFF_X1 _62347_ (.D(_00956_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1120]),
    .QN(_28915_));
 DFF_X1 _62348_ (.D(_00957_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1121]),
    .QN(_28916_));
 DFF_X1 _62349_ (.D(_00958_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1122]),
    .QN(_28917_));
 DFF_X1 _62350_ (.D(_00959_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1123]),
    .QN(_28918_));
 DFF_X1 _62351_ (.D(_00960_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1124]),
    .QN(_28919_));
 DFF_X1 _62352_ (.D(_00961_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1125]),
    .QN(_28920_));
 DFF_X1 _62353_ (.D(_00962_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1126]),
    .QN(_28921_));
 DFF_X1 _62354_ (.D(_00963_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1127]),
    .QN(_28922_));
 DFF_X1 _62355_ (.D(_00964_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1128]),
    .QN(_28923_));
 DFF_X1 _62356_ (.D(_00965_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1129]),
    .QN(_28924_));
 DFF_X1 _62357_ (.D(_00967_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1130]),
    .QN(_28925_));
 DFF_X1 _62358_ (.D(_00968_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1131]),
    .QN(_28926_));
 DFF_X1 _62359_ (.D(_00969_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1132]),
    .QN(_28927_));
 DFF_X1 _62360_ (.D(_00970_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1133]),
    .QN(_28928_));
 DFF_X1 _62361_ (.D(_00971_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1134]),
    .QN(_28929_));
 DFF_X1 _62362_ (.D(_00972_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1135]),
    .QN(_28930_));
 DFF_X1 _62363_ (.D(_00973_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1136]),
    .QN(_28931_));
 DFF_X1 _62364_ (.D(_00974_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1137]),
    .QN(_28932_));
 DFF_X1 _62365_ (.D(_00975_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1138]),
    .QN(_28933_));
 DFF_X1 _62366_ (.D(_00976_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1139]),
    .QN(_28934_));
 DFF_X1 _62367_ (.D(_00978_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1140]),
    .QN(_28935_));
 DFF_X1 _62368_ (.D(_00979_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1141]),
    .QN(_28936_));
 DFF_X1 _62369_ (.D(_00980_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1142]),
    .QN(_28937_));
 DFF_X1 _62370_ (.D(_00981_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1143]),
    .QN(_28938_));
 DFF_X1 _62371_ (.D(_00982_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1144]),
    .QN(_28939_));
 DFF_X1 _62372_ (.D(_00983_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1145]),
    .QN(_28940_));
 DFF_X1 _62373_ (.D(_00984_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1146]),
    .QN(_28941_));
 DFF_X1 _62374_ (.D(_00985_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1147]),
    .QN(_28942_));
 DFF_X1 _62375_ (.D(_00986_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1148]),
    .QN(_28943_));
 DFF_X1 _62376_ (.D(_00987_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1149]),
    .QN(_28944_));
 DFF_X1 _62377_ (.D(_00989_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1150]),
    .QN(_28945_));
 DFF_X1 _62378_ (.D(_00990_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1151]),
    .QN(_28946_));
 DFF_X1 _62379_ (.D(_00991_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1152]),
    .QN(_28947_));
 DFF_X1 _62380_ (.D(_00992_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1153]),
    .QN(_28948_));
 DFF_X1 _62381_ (.D(_00993_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1154]),
    .QN(_28949_));
 DFF_X1 _62382_ (.D(_00994_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1155]),
    .QN(_28950_));
 DFF_X1 _62383_ (.D(_00995_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1156]),
    .QN(_28951_));
 DFF_X1 _62384_ (.D(_00996_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1157]),
    .QN(_28952_));
 DFF_X1 _62385_ (.D(_00997_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1158]),
    .QN(_28953_));
 DFF_X1 _62386_ (.D(_00998_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1159]),
    .QN(_28954_));
 DFF_X1 _62387_ (.D(_01000_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1160]),
    .QN(_28955_));
 DFF_X1 _62388_ (.D(_01001_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1161]),
    .QN(_28956_));
 DFF_X1 _62389_ (.D(_01002_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1162]),
    .QN(_28957_));
 DFF_X1 _62390_ (.D(_01003_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1163]),
    .QN(_28958_));
 DFF_X1 _62391_ (.D(_01004_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1164]),
    .QN(_28959_));
 DFF_X1 _62392_ (.D(_01005_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1165]),
    .QN(_28960_));
 DFF_X1 _62393_ (.D(_01006_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1166]),
    .QN(_28961_));
 DFF_X1 _62394_ (.D(_01007_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1167]),
    .QN(_28962_));
 DFF_X1 _62395_ (.D(_01008_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1168]),
    .QN(_28963_));
 DFF_X1 _62396_ (.D(_01009_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1169]),
    .QN(_28964_));
 DFF_X1 _62397_ (.D(_01011_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1170]),
    .QN(_28965_));
 DFF_X1 _62398_ (.D(_01012_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1171]),
    .QN(_28966_));
 DFF_X1 _62399_ (.D(_01013_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1172]),
    .QN(_28967_));
 DFF_X1 _62400_ (.D(_01014_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1173]),
    .QN(_28968_));
 DFF_X1 _62401_ (.D(_01015_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1174]),
    .QN(_28969_));
 DFF_X1 _62402_ (.D(_01016_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1175]),
    .QN(_28970_));
 DFF_X1 _62403_ (.D(_01017_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1176]),
    .QN(_28971_));
 DFF_X1 _62404_ (.D(_01018_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1177]),
    .QN(_28972_));
 DFF_X1 _62405_ (.D(_01019_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1178]),
    .QN(_28973_));
 DFF_X1 _62406_ (.D(_01020_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1179]),
    .QN(_28974_));
 DFF_X1 _62407_ (.D(_01022_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1180]),
    .QN(_28975_));
 DFF_X1 _62408_ (.D(_01023_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1181]),
    .QN(_28976_));
 DFF_X1 _62409_ (.D(_01024_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1182]),
    .QN(_28977_));
 DFF_X1 _62410_ (.D(_01025_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1183]),
    .QN(_28978_));
 DFF_X1 _62411_ (.D(_01026_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1184]),
    .QN(_28979_));
 DFF_X1 _62412_ (.D(_01027_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1185]),
    .QN(_28980_));
 DFF_X1 _62413_ (.D(_01028_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1186]),
    .QN(_28981_));
 DFF_X1 _62414_ (.D(_01029_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1187]),
    .QN(_28982_));
 DFF_X1 _62415_ (.D(_01030_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1188]),
    .QN(_28983_));
 DFF_X1 _62416_ (.D(_01031_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1189]),
    .QN(_28984_));
 DFF_X1 _62417_ (.D(_01033_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1190]),
    .QN(_28985_));
 DFF_X1 _62418_ (.D(_01034_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1191]),
    .QN(_28986_));
 DFF_X1 _62419_ (.D(_01035_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1192]),
    .QN(_28987_));
 DFF_X1 _62420_ (.D(_01036_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1193]),
    .QN(_28988_));
 DFF_X1 _62421_ (.D(_01037_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1194]),
    .QN(_28989_));
 DFF_X1 _62422_ (.D(_01038_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1195]),
    .QN(_28990_));
 DFF_X1 _62423_ (.D(_01039_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1196]),
    .QN(_28991_));
 DFF_X1 _62424_ (.D(_01040_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1197]),
    .QN(_28992_));
 DFF_X1 _62425_ (.D(_01041_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1198]),
    .QN(_28993_));
 DFF_X1 _62426_ (.D(_01042_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1199]),
    .QN(_28994_));
 DFF_X1 _62427_ (.D(_01045_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1200]),
    .QN(_28995_));
 DFF_X1 _62428_ (.D(_01046_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1201]),
    .QN(_28996_));
 DFF_X1 _62429_ (.D(_01047_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1202]),
    .QN(_28997_));
 DFF_X1 _62430_ (.D(_01048_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1203]),
    .QN(_28998_));
 DFF_X1 _62431_ (.D(_01049_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1204]),
    .QN(_28999_));
 DFF_X1 _62432_ (.D(_01050_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1205]),
    .QN(_29000_));
 DFF_X1 _62433_ (.D(_01051_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1206]),
    .QN(_29001_));
 DFF_X1 _62434_ (.D(_01052_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1207]),
    .QN(_29002_));
 DFF_X1 _62435_ (.D(_01053_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1208]),
    .QN(_29003_));
 DFF_X1 _62436_ (.D(_01054_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1209]),
    .QN(_29004_));
 DFF_X1 _62437_ (.D(_01056_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1210]),
    .QN(_29005_));
 DFF_X1 _62438_ (.D(_01057_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1211]),
    .QN(_29006_));
 DFF_X1 _62439_ (.D(_01058_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1212]),
    .QN(_29007_));
 DFF_X1 _62440_ (.D(_01059_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1213]),
    .QN(_29008_));
 DFF_X1 _62441_ (.D(_01060_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1214]),
    .QN(_29009_));
 DFF_X1 _62442_ (.D(_01061_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1215]),
    .QN(_29010_));
 DFF_X1 _62443_ (.D(_01062_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1216]),
    .QN(_29011_));
 DFF_X1 _62444_ (.D(_01063_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1217]),
    .QN(_29012_));
 DFF_X1 _62445_ (.D(_01064_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1218]),
    .QN(_29013_));
 DFF_X1 _62446_ (.D(_01065_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1219]),
    .QN(_29014_));
 DFF_X1 _62447_ (.D(_01067_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1220]),
    .QN(_29015_));
 DFF_X1 _62448_ (.D(_01068_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1221]),
    .QN(_29016_));
 DFF_X1 _62449_ (.D(_01069_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1222]),
    .QN(_29017_));
 DFF_X1 _62450_ (.D(_01070_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1223]),
    .QN(_29018_));
 DFF_X1 _62451_ (.D(_01071_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1224]),
    .QN(_29019_));
 DFF_X1 _62452_ (.D(_01072_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1225]),
    .QN(_29020_));
 DFF_X1 _62453_ (.D(_01073_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1226]),
    .QN(_29021_));
 DFF_X1 _62454_ (.D(_01074_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1227]),
    .QN(_29022_));
 DFF_X1 _62455_ (.D(_01075_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1228]),
    .QN(_29023_));
 DFF_X1 _62456_ (.D(_01076_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1229]),
    .QN(_29024_));
 DFF_X1 _62457_ (.D(_01078_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1230]),
    .QN(_29025_));
 DFF_X1 _62458_ (.D(_01079_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1231]),
    .QN(_29026_));
 DFF_X1 _62459_ (.D(_01080_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1232]),
    .QN(_29027_));
 DFF_X1 _62460_ (.D(_01081_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1233]),
    .QN(_29028_));
 DFF_X1 _62461_ (.D(_01082_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1234]),
    .QN(_29029_));
 DFF_X1 _62462_ (.D(_01083_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1235]),
    .QN(_29030_));
 DFF_X1 _62463_ (.D(_01084_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1236]),
    .QN(_29031_));
 DFF_X1 _62464_ (.D(_01085_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1237]),
    .QN(_29032_));
 DFF_X1 _62465_ (.D(_01086_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1238]),
    .QN(_29033_));
 DFF_X1 _62466_ (.D(_01087_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1239]),
    .QN(_29034_));
 DFF_X1 _62467_ (.D(_01089_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1240]),
    .QN(_29035_));
 DFF_X1 _62468_ (.D(_01090_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1241]),
    .QN(_29036_));
 DFF_X1 _62469_ (.D(_01091_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1242]),
    .QN(_29037_));
 DFF_X1 _62470_ (.D(_01092_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1243]),
    .QN(_29038_));
 DFF_X1 _62471_ (.D(_01093_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1244]),
    .QN(_29039_));
 DFF_X1 _62472_ (.D(_01094_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1245]),
    .QN(_29040_));
 DFF_X1 _62473_ (.D(_01095_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1246]),
    .QN(_29041_));
 DFF_X1 _62474_ (.D(_01096_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1247]),
    .QN(_29042_));
 DFF_X1 _62475_ (.D(_01097_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1248]),
    .QN(_29043_));
 DFF_X1 _62476_ (.D(_01098_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1249]),
    .QN(_29044_));
 DFF_X1 _62477_ (.D(_01100_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1250]),
    .QN(_29045_));
 DFF_X1 _62478_ (.D(_01101_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1251]),
    .QN(_29046_));
 DFF_X1 _62479_ (.D(_01102_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1252]),
    .QN(_29047_));
 DFF_X1 _62480_ (.D(_01103_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1253]),
    .QN(_29048_));
 DFF_X1 _62481_ (.D(_01104_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1254]),
    .QN(_29049_));
 DFF_X1 _62482_ (.D(_01105_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1255]),
    .QN(_29050_));
 DFF_X1 _62483_ (.D(_01106_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1256]),
    .QN(_29051_));
 DFF_X1 _62484_ (.D(_01107_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1257]),
    .QN(_29052_));
 DFF_X1 _62485_ (.D(_01108_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1258]),
    .QN(_29053_));
 DFF_X1 _62486_ (.D(_01109_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1259]),
    .QN(_29054_));
 DFF_X1 _62487_ (.D(_01111_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1260]),
    .QN(_29055_));
 DFF_X1 _62488_ (.D(_01112_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1261]),
    .QN(_29056_));
 DFF_X1 _62489_ (.D(_01113_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1262]),
    .QN(_29057_));
 DFF_X1 _62490_ (.D(_01114_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1263]),
    .QN(_29058_));
 DFF_X1 _62491_ (.D(_01115_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1264]),
    .QN(_29059_));
 DFF_X1 _62492_ (.D(_01116_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1265]),
    .QN(_29060_));
 DFF_X1 _62493_ (.D(_01117_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1266]),
    .QN(_29061_));
 DFF_X1 _62494_ (.D(_01118_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1267]),
    .QN(_29062_));
 DFF_X1 _62495_ (.D(_01119_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1268]),
    .QN(_29063_));
 DFF_X1 _62496_ (.D(_01120_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1269]),
    .QN(_29064_));
 DFF_X1 _62497_ (.D(_01122_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1270]),
    .QN(_29065_));
 DFF_X1 _62498_ (.D(_01123_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1271]),
    .QN(_29066_));
 DFF_X1 _62499_ (.D(_01124_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1272]),
    .QN(_29067_));
 DFF_X1 _62500_ (.D(_01125_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1273]),
    .QN(_29068_));
 DFF_X1 _62501_ (.D(_01126_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1274]),
    .QN(_29069_));
 DFF_X1 _62502_ (.D(_01127_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1275]),
    .QN(_29070_));
 DFF_X1 _62503_ (.D(_01128_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1276]),
    .QN(_29071_));
 DFF_X1 _62504_ (.D(_01129_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1277]),
    .QN(_29072_));
 DFF_X1 _62505_ (.D(_01130_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1278]),
    .QN(_29073_));
 DFF_X1 _62506_ (.D(_01131_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1279]),
    .QN(_29074_));
 DFF_X1 _62507_ (.D(_01133_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1280]),
    .QN(_29075_));
 DFF_X1 _62508_ (.D(_01134_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1281]),
    .QN(_29076_));
 DFF_X1 _62509_ (.D(_01135_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1282]),
    .QN(_29077_));
 DFF_X1 _62510_ (.D(_01136_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1283]),
    .QN(_29078_));
 DFF_X1 _62511_ (.D(_01137_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1284]),
    .QN(_29079_));
 DFF_X1 _62512_ (.D(_01138_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1285]),
    .QN(_29080_));
 DFF_X1 _62513_ (.D(_01139_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1286]),
    .QN(_29081_));
 DFF_X1 _62514_ (.D(_01140_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1287]),
    .QN(_29082_));
 DFF_X1 _62515_ (.D(_01141_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1288]),
    .QN(_29083_));
 DFF_X1 _62516_ (.D(_01142_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1289]),
    .QN(_29084_));
 DFF_X1 _62517_ (.D(_01144_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1290]),
    .QN(_29085_));
 DFF_X1 _62518_ (.D(_01145_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1291]),
    .QN(_29086_));
 DFF_X1 _62519_ (.D(_01146_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1292]),
    .QN(_29087_));
 DFF_X1 _62520_ (.D(_01147_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1293]),
    .QN(_29088_));
 DFF_X1 _62521_ (.D(_01148_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1294]),
    .QN(_29089_));
 DFF_X1 _62522_ (.D(_01149_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1295]),
    .QN(_29090_));
 DFF_X1 _62523_ (.D(_01150_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1296]),
    .QN(_29091_));
 DFF_X1 _62524_ (.D(_01151_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1297]),
    .QN(_29092_));
 DFF_X1 _62525_ (.D(_01152_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1298]),
    .QN(_29093_));
 DFF_X1 _62526_ (.D(_01153_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1299]),
    .QN(_29094_));
 DFF_X1 _62527_ (.D(_01156_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1300]),
    .QN(_29095_));
 DFF_X1 _62528_ (.D(_01157_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1301]),
    .QN(_29096_));
 DFF_X1 _62529_ (.D(_01158_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1302]),
    .QN(_29097_));
 DFF_X1 _62530_ (.D(_01159_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1303]),
    .QN(_29098_));
 DFF_X1 _62531_ (.D(_01160_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1304]),
    .QN(_29099_));
 DFF_X1 _62532_ (.D(_01161_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1305]),
    .QN(_29100_));
 DFF_X1 _62533_ (.D(_01162_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1306]),
    .QN(_29101_));
 DFF_X1 _62534_ (.D(_01163_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1307]),
    .QN(_29102_));
 DFF_X1 _62535_ (.D(_01164_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1308]),
    .QN(_29103_));
 DFF_X1 _62536_ (.D(_01165_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1309]),
    .QN(_29104_));
 DFF_X1 _62537_ (.D(_01167_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1310]),
    .QN(_29105_));
 DFF_X1 _62538_ (.D(_01168_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1311]),
    .QN(_29106_));
 DFF_X1 _62539_ (.D(_01169_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1312]),
    .QN(_29107_));
 DFF_X1 _62540_ (.D(_01170_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1313]),
    .QN(_29108_));
 DFF_X1 _62541_ (.D(_01171_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1314]),
    .QN(_29109_));
 DFF_X1 _62542_ (.D(_01172_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1315]),
    .QN(_29110_));
 DFF_X1 _62543_ (.D(_01173_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1316]),
    .QN(_29111_));
 DFF_X1 _62544_ (.D(_01174_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1317]),
    .QN(_29112_));
 DFF_X1 _62545_ (.D(_01175_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1318]),
    .QN(_29113_));
 DFF_X1 _62546_ (.D(_01176_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1319]),
    .QN(_29114_));
 DFF_X1 _62547_ (.D(_01178_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1320]),
    .QN(_29115_));
 DFF_X1 _62548_ (.D(_01179_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1321]),
    .QN(_29116_));
 DFF_X1 _62549_ (.D(_01180_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1322]),
    .QN(_29117_));
 DFF_X1 _62550_ (.D(_01181_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1323]),
    .QN(_29118_));
 DFF_X1 _62551_ (.D(_01182_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1324]),
    .QN(_29119_));
 DFF_X1 _62552_ (.D(_01183_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1325]),
    .QN(_29120_));
 DFF_X1 _62553_ (.D(_01184_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1326]),
    .QN(_29121_));
 DFF_X1 _62554_ (.D(_01185_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1327]),
    .QN(_29122_));
 DFF_X1 _62555_ (.D(_01186_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1328]),
    .QN(_29123_));
 DFF_X1 _62556_ (.D(_01187_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1329]),
    .QN(_29124_));
 DFF_X1 _62557_ (.D(_01189_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1330]),
    .QN(_29125_));
 DFF_X1 _62558_ (.D(_01190_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1331]),
    .QN(_29126_));
 DFF_X1 _62559_ (.D(_01191_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1332]),
    .QN(_29127_));
 DFF_X1 _62560_ (.D(_01192_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1333]),
    .QN(_29128_));
 DFF_X1 _62561_ (.D(_01193_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1334]),
    .QN(_29129_));
 DFF_X1 _62562_ (.D(_01194_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1335]),
    .QN(_29130_));
 DFF_X1 _62563_ (.D(_01195_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1336]),
    .QN(_29131_));
 DFF_X1 _62564_ (.D(_01196_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1337]),
    .QN(_29132_));
 DFF_X1 _62565_ (.D(_01197_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1338]),
    .QN(_29133_));
 DFF_X1 _62566_ (.D(_01198_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1339]),
    .QN(_29134_));
 DFF_X1 _62567_ (.D(_01200_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1340]),
    .QN(_29135_));
 DFF_X1 _62568_ (.D(_01201_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1341]),
    .QN(_29136_));
 DFF_X1 _62569_ (.D(_01202_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1342]),
    .QN(_29137_));
 DFF_X1 _62570_ (.D(_01203_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1343]),
    .QN(_29138_));
 DFF_X1 _62571_ (.D(_01204_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1344]),
    .QN(_29139_));
 DFF_X1 _62572_ (.D(_01205_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1345]),
    .QN(_29140_));
 DFF_X1 _62573_ (.D(_01206_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1346]),
    .QN(_29141_));
 DFF_X1 _62574_ (.D(_01207_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1347]),
    .QN(_29142_));
 DFF_X1 _62575_ (.D(_01208_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1348]),
    .QN(_29143_));
 DFF_X1 _62576_ (.D(_01209_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1349]),
    .QN(_29144_));
 DFF_X1 _62577_ (.D(_01211_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1350]),
    .QN(_29145_));
 DFF_X1 _62578_ (.D(_01212_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1351]),
    .QN(_29146_));
 DFF_X1 _62579_ (.D(_01213_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1352]),
    .QN(_29147_));
 DFF_X1 _62580_ (.D(_01214_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1353]),
    .QN(_29148_));
 DFF_X1 _62581_ (.D(_01215_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1354]),
    .QN(_29149_));
 DFF_X1 _62582_ (.D(_01216_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1355]),
    .QN(_29150_));
 DFF_X1 _62583_ (.D(_01217_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1356]),
    .QN(_29151_));
 DFF_X1 _62584_ (.D(_01218_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1357]),
    .QN(_29152_));
 DFF_X1 _62585_ (.D(_01219_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1358]),
    .QN(_29153_));
 DFF_X1 _62586_ (.D(_01220_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1359]),
    .QN(_29154_));
 DFF_X1 _62587_ (.D(_01222_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1360]),
    .QN(_29155_));
 DFF_X1 _62588_ (.D(_01223_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1361]),
    .QN(_29156_));
 DFF_X1 _62589_ (.D(_01224_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1362]),
    .QN(_29157_));
 DFF_X1 _62590_ (.D(_01225_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1363]),
    .QN(_29158_));
 DFF_X1 _62591_ (.D(_01226_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1364]),
    .QN(_29159_));
 DFF_X1 _62592_ (.D(_01227_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1365]),
    .QN(_29160_));
 DFF_X1 _62593_ (.D(_01228_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1366]),
    .QN(_29161_));
 DFF_X1 _62594_ (.D(_01229_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1367]),
    .QN(_29162_));
 DFF_X1 _62595_ (.D(_01230_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1368]),
    .QN(_29163_));
 DFF_X1 _62596_ (.D(_01231_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1369]),
    .QN(_29164_));
 DFF_X1 _62597_ (.D(_01233_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1370]),
    .QN(_29165_));
 DFF_X1 _62598_ (.D(_01234_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1371]),
    .QN(_29166_));
 DFF_X1 _62599_ (.D(_01235_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1372]),
    .QN(_29167_));
 DFF_X1 _62600_ (.D(_01236_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1373]),
    .QN(_29168_));
 DFF_X1 _62601_ (.D(_01237_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1374]),
    .QN(_29169_));
 DFF_X1 _62602_ (.D(_01238_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1375]),
    .QN(_29170_));
 DFF_X1 _62603_ (.D(_01239_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1376]),
    .QN(_29171_));
 DFF_X1 _62604_ (.D(_01240_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1377]),
    .QN(_29172_));
 DFF_X1 _62605_ (.D(_01241_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1378]),
    .QN(_29173_));
 DFF_X1 _62606_ (.D(_01242_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1379]),
    .QN(_29174_));
 DFF_X1 _62607_ (.D(_01244_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1380]),
    .QN(_29175_));
 DFF_X1 _62608_ (.D(_01245_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1381]),
    .QN(_29176_));
 DFF_X1 _62609_ (.D(_01246_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1382]),
    .QN(_29177_));
 DFF_X1 _62610_ (.D(_01247_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1383]),
    .QN(_29178_));
 DFF_X1 _62611_ (.D(_01248_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1384]),
    .QN(_29179_));
 DFF_X1 _62612_ (.D(_01249_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1385]),
    .QN(_29180_));
 DFF_X1 _62613_ (.D(_01250_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1386]),
    .QN(_29181_));
 DFF_X1 _62614_ (.D(_01251_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1387]),
    .QN(_29182_));
 DFF_X1 _62615_ (.D(_01252_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1388]),
    .QN(_29183_));
 DFF_X1 _62616_ (.D(_01253_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1389]),
    .QN(_29184_));
 DFF_X1 _62617_ (.D(_01255_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1390]),
    .QN(_29185_));
 DFF_X1 _62618_ (.D(_01256_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1391]),
    .QN(_29186_));
 DFF_X1 _62619_ (.D(_01257_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1392]),
    .QN(_29187_));
 DFF_X1 _62620_ (.D(_01258_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1393]),
    .QN(_29188_));
 DFF_X1 _62621_ (.D(_01259_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1394]),
    .QN(_29189_));
 DFF_X1 _62622_ (.D(_01260_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1395]),
    .QN(_29190_));
 DFF_X1 _62623_ (.D(_01261_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1396]),
    .QN(_29191_));
 DFF_X1 _62624_ (.D(_01262_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1397]),
    .QN(_29192_));
 DFF_X1 _62625_ (.D(_01263_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1398]),
    .QN(_29193_));
 DFF_X1 _62626_ (.D(_01264_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1399]),
    .QN(_29194_));
 DFF_X1 _62627_ (.D(_01267_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1400]),
    .QN(_29195_));
 DFF_X1 _62628_ (.D(_01268_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1401]),
    .QN(_29196_));
 DFF_X1 _62629_ (.D(_01269_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1402]),
    .QN(_29197_));
 DFF_X1 _62630_ (.D(_01270_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1403]),
    .QN(_29198_));
 DFF_X1 _62631_ (.D(_01271_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1404]),
    .QN(_29199_));
 DFF_X1 _62632_ (.D(_01272_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1405]),
    .QN(_29200_));
 DFF_X1 _62633_ (.D(_01273_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1406]),
    .QN(_29201_));
 DFF_X1 _62634_ (.D(_01274_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1407]),
    .QN(_29202_));
 DFF_X1 _62635_ (.D(_01275_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1408]),
    .QN(_29203_));
 DFF_X1 _62636_ (.D(_01276_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1409]),
    .QN(_29204_));
 DFF_X1 _62637_ (.D(_01278_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1410]),
    .QN(_29205_));
 DFF_X1 _62638_ (.D(_01279_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1411]),
    .QN(_29206_));
 DFF_X1 _62639_ (.D(_01280_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1412]),
    .QN(_29207_));
 DFF_X1 _62640_ (.D(_01281_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1413]),
    .QN(_29208_));
 DFF_X1 _62641_ (.D(_01282_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1414]),
    .QN(_29209_));
 DFF_X1 _62642_ (.D(_01283_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1415]),
    .QN(_29210_));
 DFF_X1 _62643_ (.D(_01284_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1416]),
    .QN(_29211_));
 DFF_X1 _62644_ (.D(_01285_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1417]),
    .QN(_29212_));
 DFF_X1 _62645_ (.D(_01286_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1418]),
    .QN(_29213_));
 DFF_X1 _62646_ (.D(_01287_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1419]),
    .QN(_29214_));
 DFF_X1 _62647_ (.D(_01289_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1420]),
    .QN(_29215_));
 DFF_X1 _62648_ (.D(_01290_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1421]),
    .QN(_29216_));
 DFF_X1 _62649_ (.D(_01291_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1422]),
    .QN(_29217_));
 DFF_X1 _62650_ (.D(_01292_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1423]),
    .QN(_29218_));
 DFF_X1 _62651_ (.D(_01293_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1424]),
    .QN(_29219_));
 DFF_X1 _62652_ (.D(_01294_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1425]),
    .QN(_29220_));
 DFF_X1 _62653_ (.D(_01295_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1426]),
    .QN(_29221_));
 DFF_X1 _62654_ (.D(_01296_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1427]),
    .QN(_29222_));
 DFF_X1 _62655_ (.D(_01297_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1428]),
    .QN(_29223_));
 DFF_X1 _62656_ (.D(_01298_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1429]),
    .QN(_29224_));
 DFF_X1 _62657_ (.D(_01300_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1430]),
    .QN(_29225_));
 DFF_X1 _62658_ (.D(_01301_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1431]),
    .QN(_29226_));
 DFF_X1 _62659_ (.D(_01302_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1432]),
    .QN(_29227_));
 DFF_X1 _62660_ (.D(_01303_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1433]),
    .QN(_29228_));
 DFF_X1 _62661_ (.D(_01304_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1434]),
    .QN(_29229_));
 DFF_X1 _62662_ (.D(_01305_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1435]),
    .QN(_29230_));
 DFF_X1 _62663_ (.D(_01306_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1436]),
    .QN(_29231_));
 DFF_X1 _62664_ (.D(_01307_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1437]),
    .QN(_29232_));
 DFF_X1 _62665_ (.D(_01308_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1438]),
    .QN(_29233_));
 DFF_X1 _62666_ (.D(_01309_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1439]),
    .QN(_29234_));
 DFF_X1 _62667_ (.D(_01311_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1440]),
    .QN(_29235_));
 DFF_X1 _62668_ (.D(_01312_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1441]),
    .QN(_29236_));
 DFF_X1 _62669_ (.D(_01313_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1442]),
    .QN(_29237_));
 DFF_X1 _62670_ (.D(_01314_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1443]),
    .QN(_29238_));
 DFF_X1 _62671_ (.D(_01315_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1444]),
    .QN(_29239_));
 DFF_X1 _62672_ (.D(_01316_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1445]),
    .QN(_29240_));
 DFF_X1 _62673_ (.D(_01317_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1446]),
    .QN(_29241_));
 DFF_X1 _62674_ (.D(_01318_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1447]),
    .QN(_29242_));
 DFF_X1 _62675_ (.D(_01319_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1448]),
    .QN(_29243_));
 DFF_X1 _62676_ (.D(_01320_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1449]),
    .QN(_29244_));
 DFF_X1 _62677_ (.D(_01322_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1450]),
    .QN(_29245_));
 DFF_X1 _62678_ (.D(_01323_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1451]),
    .QN(_29246_));
 DFF_X1 _62679_ (.D(_01324_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1452]),
    .QN(_29247_));
 DFF_X1 _62680_ (.D(_01325_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1453]),
    .QN(_29248_));
 DFF_X1 _62681_ (.D(_01326_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1454]),
    .QN(_29249_));
 DFF_X1 _62682_ (.D(_01327_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1455]),
    .QN(_29250_));
 DFF_X1 _62683_ (.D(_01328_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1456]),
    .QN(_29251_));
 DFF_X1 _62684_ (.D(_01329_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1457]),
    .QN(_29252_));
 DFF_X1 _62685_ (.D(_01330_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1458]),
    .QN(_29253_));
 DFF_X1 _62686_ (.D(_01331_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1459]),
    .QN(_29254_));
 DFF_X1 _62687_ (.D(_01333_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1460]),
    .QN(_29255_));
 DFF_X1 _62688_ (.D(_01334_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1461]),
    .QN(_29256_));
 DFF_X1 _62689_ (.D(_01335_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1462]),
    .QN(_29257_));
 DFF_X1 _62690_ (.D(_01336_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1463]),
    .QN(_29258_));
 DFF_X1 _62691_ (.D(_01337_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1464]),
    .QN(_29259_));
 DFF_X1 _62692_ (.D(_01338_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1465]),
    .QN(_29260_));
 DFF_X1 _62693_ (.D(_01339_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1466]),
    .QN(_29261_));
 DFF_X1 _62694_ (.D(_01340_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1467]),
    .QN(_29262_));
 DFF_X1 _62695_ (.D(_01341_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1468]),
    .QN(_29263_));
 DFF_X1 _62696_ (.D(_01342_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1469]),
    .QN(_29264_));
 DFF_X1 _62697_ (.D(_01344_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1470]),
    .QN(_29265_));
 DFF_X1 _62698_ (.D(_01345_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1471]),
    .QN(_29266_));
 DFF_X1 _62699_ (.D(_01346_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1472]),
    .QN(_29267_));
 DFF_X1 _62700_ (.D(_01347_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1473]),
    .QN(_29268_));
 DFF_X1 _62701_ (.D(_01348_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1474]),
    .QN(_29269_));
 DFF_X1 _62702_ (.D(_01349_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1475]),
    .QN(_29270_));
 DFF_X1 _62703_ (.D(_01350_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1476]),
    .QN(_29271_));
 DFF_X1 _62704_ (.D(_01351_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1477]),
    .QN(_29272_));
 DFF_X1 _62705_ (.D(_01352_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1478]),
    .QN(_29273_));
 DFF_X1 _62706_ (.D(_01353_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1479]),
    .QN(_29274_));
 DFF_X1 _62707_ (.D(_01355_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1480]),
    .QN(_29275_));
 DFF_X1 _62708_ (.D(_01356_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1481]),
    .QN(_29276_));
 DFF_X1 _62709_ (.D(_01357_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1482]),
    .QN(_29277_));
 DFF_X1 _62710_ (.D(_01358_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1483]),
    .QN(_29278_));
 DFF_X1 _62711_ (.D(_01359_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1484]),
    .QN(_29279_));
 DFF_X1 _62712_ (.D(_01360_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1485]),
    .QN(_29280_));
 DFF_X1 _62713_ (.D(_01361_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1486]),
    .QN(_29281_));
 DFF_X1 _62714_ (.D(_01362_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1487]),
    .QN(_29282_));
 DFF_X1 _62715_ (.D(_01363_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1488]),
    .QN(_29283_));
 DFF_X1 _62716_ (.D(_01364_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1489]),
    .QN(_29284_));
 DFF_X1 _62717_ (.D(_01366_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1490]),
    .QN(_29285_));
 DFF_X1 _62718_ (.D(_01367_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1491]),
    .QN(_29286_));
 DFF_X1 _62719_ (.D(_01368_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1492]),
    .QN(_29287_));
 DFF_X1 _62720_ (.D(_01369_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1493]),
    .QN(_29288_));
 DFF_X1 _62721_ (.D(_01370_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1494]),
    .QN(_29289_));
 DFF_X1 _62722_ (.D(_01371_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1495]),
    .QN(_29290_));
 DFF_X1 _62723_ (.D(_01372_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1496]),
    .QN(_29291_));
 DFF_X1 _62724_ (.D(_01373_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1497]),
    .QN(_29292_));
 DFF_X1 _62725_ (.D(_01374_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1498]),
    .QN(_29293_));
 DFF_X1 _62726_ (.D(_01375_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1499]),
    .QN(_29294_));
 DFF_X1 _62727_ (.D(_01378_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1500]),
    .QN(_29295_));
 DFF_X1 _62728_ (.D(_01379_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1501]),
    .QN(_29296_));
 DFF_X1 _62729_ (.D(_01380_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1502]),
    .QN(_29297_));
 DFF_X1 _62730_ (.D(_01381_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1503]),
    .QN(_29298_));
 DFF_X1 _62731_ (.D(_01382_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1504]),
    .QN(_29299_));
 DFF_X1 _62732_ (.D(_01383_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1505]),
    .QN(_29300_));
 DFF_X1 _62733_ (.D(_01384_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1506]),
    .QN(_29301_));
 DFF_X1 _62734_ (.D(_01385_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1507]),
    .QN(_29302_));
 DFF_X1 _62735_ (.D(_01386_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1508]),
    .QN(_29303_));
 DFF_X1 _62736_ (.D(_01387_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1509]),
    .QN(_29304_));
 DFF_X1 _62737_ (.D(_01389_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1510]),
    .QN(_29305_));
 DFF_X1 _62738_ (.D(_01390_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1511]),
    .QN(_29306_));
 DFF_X1 _62739_ (.D(_01391_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1512]),
    .QN(_29307_));
 DFF_X1 _62740_ (.D(_01392_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1513]),
    .QN(_29308_));
 DFF_X1 _62741_ (.D(_01393_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1514]),
    .QN(_29309_));
 DFF_X1 _62742_ (.D(_01394_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1515]),
    .QN(_29310_));
 DFF_X1 _62743_ (.D(_01395_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1516]),
    .QN(_29311_));
 DFF_X1 _62744_ (.D(_01396_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1517]),
    .QN(_29312_));
 DFF_X1 _62745_ (.D(_01397_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1518]),
    .QN(_29313_));
 DFF_X1 _62746_ (.D(_01398_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1519]),
    .QN(_29314_));
 DFF_X1 _62747_ (.D(_01400_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1520]),
    .QN(_29315_));
 DFF_X1 _62748_ (.D(_01401_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1521]),
    .QN(_29316_));
 DFF_X1 _62749_ (.D(_01402_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1522]),
    .QN(_29317_));
 DFF_X1 _62750_ (.D(_01403_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1523]),
    .QN(_29318_));
 DFF_X1 _62751_ (.D(_01404_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1524]),
    .QN(_29319_));
 DFF_X1 _62752_ (.D(_01405_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1525]),
    .QN(_29320_));
 DFF_X1 _62753_ (.D(_01406_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1526]),
    .QN(_29321_));
 DFF_X1 _62754_ (.D(_01407_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1527]),
    .QN(_29322_));
 DFF_X1 _62755_ (.D(_01408_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1528]),
    .QN(_29323_));
 DFF_X1 _62756_ (.D(_01409_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1529]),
    .QN(_29324_));
 DFF_X1 _62757_ (.D(_01411_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1530]),
    .QN(_29325_));
 DFF_X1 _62758_ (.D(_01412_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1531]),
    .QN(_29326_));
 DFF_X1 _62759_ (.D(_01413_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1532]),
    .QN(_29327_));
 DFF_X1 _62760_ (.D(_01414_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1533]),
    .QN(_29328_));
 DFF_X1 _62761_ (.D(_01415_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1534]),
    .QN(_29329_));
 DFF_X1 _62762_ (.D(_01416_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1535]),
    .QN(_29330_));
 DFF_X1 _62763_ (.D(_01417_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1536]),
    .QN(_29331_));
 DFF_X1 _62764_ (.D(_01418_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1537]),
    .QN(_29332_));
 DFF_X1 _62765_ (.D(_01419_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1538]),
    .QN(_29333_));
 DFF_X1 _62766_ (.D(_01420_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1539]),
    .QN(_29334_));
 DFF_X1 _62767_ (.D(_01422_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1540]),
    .QN(_29335_));
 DFF_X1 _62768_ (.D(_01423_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1541]),
    .QN(_29336_));
 DFF_X1 _62769_ (.D(_01424_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1542]),
    .QN(_29337_));
 DFF_X1 _62770_ (.D(_01425_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1543]),
    .QN(_29338_));
 DFF_X1 _62771_ (.D(_01426_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1544]),
    .QN(_29339_));
 DFF_X1 _62772_ (.D(_01427_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1545]),
    .QN(_29340_));
 DFF_X1 _62773_ (.D(_01428_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1546]),
    .QN(_29341_));
 DFF_X1 _62774_ (.D(_01429_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1547]),
    .QN(_29342_));
 DFF_X1 _62775_ (.D(_01430_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1548]),
    .QN(_29343_));
 DFF_X1 _62776_ (.D(_01431_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1549]),
    .QN(_29344_));
 DFF_X1 _62777_ (.D(_01433_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1550]),
    .QN(_29345_));
 DFF_X1 _62778_ (.D(_01434_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1551]),
    .QN(_29346_));
 DFF_X1 _62779_ (.D(_01435_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1552]),
    .QN(_29347_));
 DFF_X1 _62780_ (.D(_01436_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1553]),
    .QN(_29348_));
 DFF_X1 _62781_ (.D(_01437_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1554]),
    .QN(_29349_));
 DFF_X1 _62782_ (.D(_01438_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1555]),
    .QN(_29350_));
 DFF_X1 _62783_ (.D(_01439_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1556]),
    .QN(_29351_));
 DFF_X1 _62784_ (.D(_01440_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1557]),
    .QN(_29352_));
 DFF_X1 _62785_ (.D(_01441_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1558]),
    .QN(_29353_));
 DFF_X1 _62786_ (.D(_01442_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1559]),
    .QN(_29354_));
 DFF_X1 _62787_ (.D(_01444_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1560]),
    .QN(_29355_));
 DFF_X1 _62788_ (.D(_01445_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1561]),
    .QN(_29356_));
 DFF_X1 _62789_ (.D(_01446_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1562]),
    .QN(_29357_));
 DFF_X1 _62790_ (.D(_01447_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1563]),
    .QN(_29358_));
 DFF_X1 _62791_ (.D(_01448_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1564]),
    .QN(_29359_));
 DFF_X1 _62792_ (.D(_01449_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1565]),
    .QN(_29360_));
 DFF_X1 _62793_ (.D(_01450_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1566]),
    .QN(_29361_));
 DFF_X1 _62794_ (.D(_01451_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1567]),
    .QN(_29362_));
 DFF_X1 _62795_ (.D(_01452_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1568]),
    .QN(_29363_));
 DFF_X1 _62796_ (.D(_01453_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1569]),
    .QN(_29364_));
 DFF_X1 _62797_ (.D(_01455_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1570]),
    .QN(_29365_));
 DFF_X1 _62798_ (.D(_01456_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1571]),
    .QN(_29366_));
 DFF_X1 _62799_ (.D(_01457_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1572]),
    .QN(_29367_));
 DFF_X1 _62800_ (.D(_01458_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1573]),
    .QN(_29368_));
 DFF_X1 _62801_ (.D(_01459_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1574]),
    .QN(_29369_));
 DFF_X1 _62802_ (.D(_01460_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1575]),
    .QN(_29370_));
 DFF_X1 _62803_ (.D(_01461_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1576]),
    .QN(_29371_));
 DFF_X1 _62804_ (.D(_01462_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1577]),
    .QN(_29372_));
 DFF_X1 _62805_ (.D(_01463_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1578]),
    .QN(_29373_));
 DFF_X1 _62806_ (.D(_01464_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1579]),
    .QN(_29374_));
 DFF_X1 _62807_ (.D(_01466_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1580]),
    .QN(_29375_));
 DFF_X1 _62808_ (.D(_01467_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1581]),
    .QN(_29376_));
 DFF_X1 _62809_ (.D(_01468_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1582]),
    .QN(_29377_));
 DFF_X1 _62810_ (.D(_01469_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1583]),
    .QN(_29378_));
 DFF_X1 _62811_ (.D(_01470_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1584]),
    .QN(_29379_));
 DFF_X1 _62812_ (.D(_01471_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1585]),
    .QN(_29380_));
 DFF_X1 _62813_ (.D(_01472_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1586]),
    .QN(_29381_));
 DFF_X1 _62814_ (.D(_01473_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1587]),
    .QN(_29382_));
 DFF_X1 _62815_ (.D(_01474_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1588]),
    .QN(_29383_));
 DFF_X1 _62816_ (.D(_01475_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1589]),
    .QN(_29384_));
 DFF_X1 _62817_ (.D(_01477_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1590]),
    .QN(_29385_));
 DFF_X1 _62818_ (.D(_01478_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1591]),
    .QN(_29386_));
 DFF_X1 _62819_ (.D(_01479_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1592]),
    .QN(_29387_));
 DFF_X1 _62820_ (.D(_01480_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1593]),
    .QN(_29388_));
 DFF_X1 _62821_ (.D(_01481_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1594]),
    .QN(_29389_));
 DFF_X1 _62822_ (.D(_01482_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1595]),
    .QN(_29390_));
 DFF_X1 _62823_ (.D(_01483_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1596]),
    .QN(_29391_));
 DFF_X1 _62824_ (.D(_01484_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1597]),
    .QN(_29392_));
 DFF_X1 _62825_ (.D(_01485_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1598]),
    .QN(_29393_));
 DFF_X1 _62826_ (.D(_01486_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1599]),
    .QN(_29394_));
 DFF_X1 _62827_ (.D(_01489_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1600]),
    .QN(_29395_));
 DFF_X1 _62828_ (.D(_01490_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1601]),
    .QN(_29396_));
 DFF_X1 _62829_ (.D(_01491_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1602]),
    .QN(_29397_));
 DFF_X1 _62830_ (.D(_01492_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1603]),
    .QN(_29398_));
 DFF_X1 _62831_ (.D(_01493_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1604]),
    .QN(_29399_));
 DFF_X1 _62832_ (.D(_01494_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1605]),
    .QN(_29400_));
 DFF_X1 _62833_ (.D(_01495_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1606]),
    .QN(_29401_));
 DFF_X1 _62834_ (.D(_01496_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1607]),
    .QN(_29402_));
 DFF_X1 _62835_ (.D(_01497_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1608]),
    .QN(_29403_));
 DFF_X1 _62836_ (.D(_01498_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1609]),
    .QN(_29404_));
 DFF_X1 _62837_ (.D(_01500_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1610]),
    .QN(_29405_));
 DFF_X1 _62838_ (.D(_01501_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1611]),
    .QN(_29406_));
 DFF_X1 _62839_ (.D(_01502_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1612]),
    .QN(_29407_));
 DFF_X1 _62840_ (.D(_01503_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1613]),
    .QN(_29408_));
 DFF_X1 _62841_ (.D(_01504_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1614]),
    .QN(_29409_));
 DFF_X1 _62842_ (.D(_01505_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1615]),
    .QN(_29410_));
 DFF_X1 _62843_ (.D(_01506_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1616]),
    .QN(_29411_));
 DFF_X1 _62844_ (.D(_01507_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1617]),
    .QN(_29412_));
 DFF_X1 _62845_ (.D(_01508_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1618]),
    .QN(_29413_));
 DFF_X1 _62846_ (.D(_01509_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1619]),
    .QN(_29414_));
 DFF_X1 _62847_ (.D(_01511_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1620]),
    .QN(_29415_));
 DFF_X1 _62848_ (.D(_01512_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1621]),
    .QN(_29416_));
 DFF_X1 _62849_ (.D(_01513_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1622]),
    .QN(_29417_));
 DFF_X1 _62850_ (.D(_01514_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1623]),
    .QN(_29418_));
 DFF_X1 _62851_ (.D(_01515_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1624]),
    .QN(_29419_));
 DFF_X1 _62852_ (.D(_01516_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1625]),
    .QN(_29420_));
 DFF_X1 _62853_ (.D(_01517_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1626]),
    .QN(_29421_));
 DFF_X1 _62854_ (.D(_01518_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1627]),
    .QN(_29422_));
 DFF_X1 _62855_ (.D(_01519_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1628]),
    .QN(_29423_));
 DFF_X1 _62856_ (.D(_01520_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1629]),
    .QN(_29424_));
 DFF_X1 _62857_ (.D(_01522_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1630]),
    .QN(_29425_));
 DFF_X1 _62858_ (.D(_01523_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1631]),
    .QN(_29426_));
 DFF_X1 _62859_ (.D(_01524_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1632]),
    .QN(_29427_));
 DFF_X1 _62860_ (.D(_01525_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1633]),
    .QN(_29428_));
 DFF_X1 _62861_ (.D(_01526_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1634]),
    .QN(_29429_));
 DFF_X1 _62862_ (.D(_01527_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1635]),
    .QN(_29430_));
 DFF_X1 _62863_ (.D(_01528_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1636]),
    .QN(_29431_));
 DFF_X1 _62864_ (.D(_01529_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1637]),
    .QN(_29432_));
 DFF_X1 _62865_ (.D(_01530_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1638]),
    .QN(_29433_));
 DFF_X1 _62866_ (.D(_01531_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1639]),
    .QN(_29434_));
 DFF_X1 _62867_ (.D(_01533_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1640]),
    .QN(_29435_));
 DFF_X1 _62868_ (.D(_01534_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1641]),
    .QN(_29436_));
 DFF_X1 _62869_ (.D(_01535_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1642]),
    .QN(_29437_));
 DFF_X1 _62870_ (.D(_01536_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1643]),
    .QN(_29438_));
 DFF_X1 _62871_ (.D(_01537_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1644]),
    .QN(_29439_));
 DFF_X1 _62872_ (.D(_01538_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1645]),
    .QN(_29440_));
 DFF_X1 _62873_ (.D(_01539_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1646]),
    .QN(_29441_));
 DFF_X1 _62874_ (.D(_01540_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1647]),
    .QN(_29442_));
 DFF_X1 _62875_ (.D(_01541_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1648]),
    .QN(_29443_));
 DFF_X1 _62876_ (.D(_01542_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1649]),
    .QN(_29444_));
 DFF_X1 _62877_ (.D(_01544_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1650]),
    .QN(_29445_));
 DFF_X1 _62878_ (.D(_01545_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1651]),
    .QN(_29446_));
 DFF_X1 _62879_ (.D(_01546_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1652]),
    .QN(_29447_));
 DFF_X1 _62880_ (.D(_01547_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1653]),
    .QN(_29448_));
 DFF_X1 _62881_ (.D(_01548_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1654]),
    .QN(_29449_));
 DFF_X1 _62882_ (.D(_01549_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1655]),
    .QN(_29450_));
 DFF_X1 _62883_ (.D(_01550_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1656]),
    .QN(_29451_));
 DFF_X1 _62884_ (.D(_01551_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1657]),
    .QN(_29452_));
 DFF_X1 _62885_ (.D(_01552_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1658]),
    .QN(_29453_));
 DFF_X1 _62886_ (.D(_01553_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1659]),
    .QN(_29454_));
 DFF_X1 _62887_ (.D(_01555_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1660]),
    .QN(_29455_));
 DFF_X1 _62888_ (.D(_01556_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1661]),
    .QN(_29456_));
 DFF_X1 _62889_ (.D(_01557_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1662]),
    .QN(_29457_));
 DFF_X1 _62890_ (.D(_01558_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1663]),
    .QN(_29458_));
 DFF_X1 _62891_ (.D(_01559_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1664]),
    .QN(_29459_));
 DFF_X1 _62892_ (.D(_01560_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1665]),
    .QN(_29460_));
 DFF_X1 _62893_ (.D(_01561_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1666]),
    .QN(_29461_));
 DFF_X1 _62894_ (.D(_01562_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1667]),
    .QN(_29462_));
 DFF_X1 _62895_ (.D(_01563_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1668]),
    .QN(_29463_));
 DFF_X1 _62896_ (.D(_01564_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1669]),
    .QN(_29464_));
 DFF_X1 _62897_ (.D(_01566_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1670]),
    .QN(_29465_));
 DFF_X1 _62898_ (.D(_01567_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1671]),
    .QN(_29466_));
 DFF_X1 _62899_ (.D(_01568_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1672]),
    .QN(_29467_));
 DFF_X1 _62900_ (.D(_01569_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1673]),
    .QN(_29468_));
 DFF_X1 _62901_ (.D(_01570_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1674]),
    .QN(_29469_));
 DFF_X1 _62902_ (.D(_01571_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1675]),
    .QN(_29470_));
 DFF_X1 _62903_ (.D(_01572_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1676]),
    .QN(_29471_));
 DFF_X1 _62904_ (.D(_01573_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1677]),
    .QN(_29472_));
 DFF_X1 _62905_ (.D(_01574_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1678]),
    .QN(_29473_));
 DFF_X1 _62906_ (.D(_01575_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1679]),
    .QN(_29474_));
 DFF_X1 _62907_ (.D(_01577_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1680]),
    .QN(_29475_));
 DFF_X1 _62908_ (.D(_01578_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1681]),
    .QN(_29476_));
 DFF_X1 _62909_ (.D(_01579_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1682]),
    .QN(_29477_));
 DFF_X1 _62910_ (.D(_01580_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1683]),
    .QN(_29478_));
 DFF_X1 _62911_ (.D(_01581_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1684]),
    .QN(_29479_));
 DFF_X1 _62912_ (.D(_01582_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1685]),
    .QN(_29480_));
 DFF_X1 _62913_ (.D(_01583_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1686]),
    .QN(_29481_));
 DFF_X1 _62914_ (.D(_01584_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1687]),
    .QN(_29482_));
 DFF_X1 _62915_ (.D(_01585_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1688]),
    .QN(_29483_));
 DFF_X1 _62916_ (.D(_01586_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1689]),
    .QN(_29484_));
 DFF_X1 _62917_ (.D(_01588_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1690]),
    .QN(_29485_));
 DFF_X1 _62918_ (.D(_01589_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1691]),
    .QN(_29486_));
 DFF_X1 _62919_ (.D(_01590_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1692]),
    .QN(_29487_));
 DFF_X1 _62920_ (.D(_01591_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1693]),
    .QN(_29488_));
 DFF_X1 _62921_ (.D(_01592_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1694]),
    .QN(_29489_));
 DFF_X1 _62922_ (.D(_01593_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1695]),
    .QN(_29490_));
 DFF_X1 _62923_ (.D(_01594_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1696]),
    .QN(_29491_));
 DFF_X1 _62924_ (.D(_01595_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1697]),
    .QN(_29492_));
 DFF_X1 _62925_ (.D(_01596_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1698]),
    .QN(_29493_));
 DFF_X1 _62926_ (.D(_01597_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1699]),
    .QN(_29494_));
 DFF_X1 _62927_ (.D(_01600_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1700]),
    .QN(_29495_));
 DFF_X1 _62928_ (.D(_01601_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1701]),
    .QN(_29496_));
 DFF_X1 _62929_ (.D(_01602_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1702]),
    .QN(_29497_));
 DFF_X1 _62930_ (.D(_01603_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1703]),
    .QN(_29498_));
 DFF_X1 _62931_ (.D(_01604_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1704]),
    .QN(_29499_));
 DFF_X1 _62932_ (.D(_01605_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1705]),
    .QN(_29500_));
 DFF_X1 _62933_ (.D(_01606_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1706]),
    .QN(_29501_));
 DFF_X1 _62934_ (.D(_01607_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1707]),
    .QN(_29502_));
 DFF_X1 _62935_ (.D(_01608_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1708]),
    .QN(_29503_));
 DFF_X1 _62936_ (.D(_01609_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1709]),
    .QN(_29504_));
 DFF_X1 _62937_ (.D(_01611_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1710]),
    .QN(_29505_));
 DFF_X1 _62938_ (.D(_01612_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1711]),
    .QN(_29506_));
 DFF_X1 _62939_ (.D(_01613_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1712]),
    .QN(_29507_));
 DFF_X1 _62940_ (.D(_01614_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1713]),
    .QN(_29508_));
 DFF_X1 _62941_ (.D(_01615_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1714]),
    .QN(_29509_));
 DFF_X1 _62942_ (.D(_01616_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1715]),
    .QN(_29510_));
 DFF_X1 _62943_ (.D(_01617_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1716]),
    .QN(_29511_));
 DFF_X1 _62944_ (.D(_01618_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1717]),
    .QN(_29512_));
 DFF_X1 _62945_ (.D(_01619_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1718]),
    .QN(_29513_));
 DFF_X1 _62946_ (.D(_01620_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1719]),
    .QN(_29514_));
 DFF_X1 _62947_ (.D(_01622_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1720]),
    .QN(_29515_));
 DFF_X1 _62948_ (.D(_01623_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1721]),
    .QN(_29516_));
 DFF_X1 _62949_ (.D(_01624_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1722]),
    .QN(_29517_));
 DFF_X1 _62950_ (.D(_01625_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1723]),
    .QN(_29518_));
 DFF_X1 _62951_ (.D(_01626_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1724]),
    .QN(_29519_));
 DFF_X1 _62952_ (.D(_01627_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1725]),
    .QN(_29520_));
 DFF_X1 _62953_ (.D(_01628_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1726]),
    .QN(_29521_));
 DFF_X1 _62954_ (.D(_01629_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1727]),
    .QN(_29522_));
 DFF_X1 _62955_ (.D(_01630_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1728]),
    .QN(_29523_));
 DFF_X1 _62956_ (.D(_01631_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1729]),
    .QN(_29524_));
 DFF_X1 _62957_ (.D(_01633_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1730]),
    .QN(_29525_));
 DFF_X1 _62958_ (.D(_01634_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1731]),
    .QN(_29526_));
 DFF_X1 _62959_ (.D(_01635_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1732]),
    .QN(_29527_));
 DFF_X1 _62960_ (.D(_01636_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1733]),
    .QN(_29528_));
 DFF_X1 _62961_ (.D(_01637_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1734]),
    .QN(_29529_));
 DFF_X1 _62962_ (.D(_01638_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1735]),
    .QN(_29530_));
 DFF_X1 _62963_ (.D(_01639_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1736]),
    .QN(_29531_));
 DFF_X1 _62964_ (.D(_01640_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1737]),
    .QN(_29532_));
 DFF_X1 _62965_ (.D(_01641_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1738]),
    .QN(_29533_));
 DFF_X1 _62966_ (.D(_01642_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1739]),
    .QN(_29534_));
 DFF_X1 _62967_ (.D(_01644_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1740]),
    .QN(_29535_));
 DFF_X1 _62968_ (.D(_01645_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1741]),
    .QN(_29536_));
 DFF_X1 _62969_ (.D(_01646_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1742]),
    .QN(_29537_));
 DFF_X1 _62970_ (.D(_01647_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1743]),
    .QN(_29538_));
 DFF_X1 _62971_ (.D(_01648_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1744]),
    .QN(_29539_));
 DFF_X1 _62972_ (.D(_01649_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1745]),
    .QN(_29540_));
 DFF_X1 _62973_ (.D(_01650_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1746]),
    .QN(_29541_));
 DFF_X1 _62974_ (.D(_01651_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1747]),
    .QN(_29542_));
 DFF_X1 _62975_ (.D(_01652_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1748]),
    .QN(_29543_));
 DFF_X1 _62976_ (.D(_01653_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1749]),
    .QN(_29544_));
 DFF_X1 _62977_ (.D(_01655_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1750]),
    .QN(_29545_));
 DFF_X1 _62978_ (.D(_01656_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1751]),
    .QN(_29546_));
 DFF_X1 _62979_ (.D(_01657_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1752]),
    .QN(_29547_));
 DFF_X1 _62980_ (.D(_01658_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1753]),
    .QN(_29548_));
 DFF_X1 _62981_ (.D(_01659_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1754]),
    .QN(_29549_));
 DFF_X1 _62982_ (.D(_01660_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1755]),
    .QN(_29550_));
 DFF_X1 _62983_ (.D(_01661_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1756]),
    .QN(_29551_));
 DFF_X1 _62984_ (.D(_01662_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1757]),
    .QN(_29552_));
 DFF_X1 _62985_ (.D(_01663_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1758]),
    .QN(_29553_));
 DFF_X1 _62986_ (.D(_01664_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1759]),
    .QN(_29554_));
 DFF_X1 _62987_ (.D(_01666_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1760]),
    .QN(_29555_));
 DFF_X1 _62988_ (.D(_01667_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1761]),
    .QN(_29556_));
 DFF_X1 _62989_ (.D(_01668_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1762]),
    .QN(_29557_));
 DFF_X1 _62990_ (.D(_01669_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1763]),
    .QN(_29558_));
 DFF_X1 _62991_ (.D(_01670_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1764]),
    .QN(_29559_));
 DFF_X1 _62992_ (.D(_01671_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1765]),
    .QN(_29560_));
 DFF_X1 _62993_ (.D(_01672_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1766]),
    .QN(_29561_));
 DFF_X1 _62994_ (.D(_01673_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1767]),
    .QN(_29562_));
 DFF_X1 _62995_ (.D(_01674_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1768]),
    .QN(_29563_));
 DFF_X1 _62996_ (.D(_01675_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1769]),
    .QN(_29564_));
 DFF_X1 _62997_ (.D(_01677_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1770]),
    .QN(_29565_));
 DFF_X1 _62998_ (.D(_01678_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1771]),
    .QN(_29566_));
 DFF_X1 _62999_ (.D(_01679_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1772]),
    .QN(_29567_));
 DFF_X1 _63000_ (.D(_01680_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1773]),
    .QN(_29568_));
 DFF_X1 _63001_ (.D(_01681_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1774]),
    .QN(_29569_));
 DFF_X1 _63002_ (.D(_01682_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1775]),
    .QN(_29570_));
 DFF_X1 _63003_ (.D(_01683_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1776]),
    .QN(_29571_));
 DFF_X1 _63004_ (.D(_01684_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1777]),
    .QN(_29572_));
 DFF_X1 _63005_ (.D(_01685_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1778]),
    .QN(_29573_));
 DFF_X1 _63006_ (.D(_01686_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1779]),
    .QN(_29574_));
 DFF_X1 _63007_ (.D(_01688_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1780]),
    .QN(_29575_));
 DFF_X1 _63008_ (.D(_01689_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1781]),
    .QN(_29576_));
 DFF_X1 _63009_ (.D(_01690_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1782]),
    .QN(_29577_));
 DFF_X1 _63010_ (.D(_01691_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1783]),
    .QN(_29578_));
 DFF_X1 _63011_ (.D(_01692_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1784]),
    .QN(_29579_));
 DFF_X1 _63012_ (.D(_01693_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1785]),
    .QN(_29580_));
 DFF_X1 _63013_ (.D(_01694_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1786]),
    .QN(_29581_));
 DFF_X1 _63014_ (.D(_01695_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1787]),
    .QN(_29582_));
 DFF_X1 _63015_ (.D(_01696_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1788]),
    .QN(_29583_));
 DFF_X1 _63016_ (.D(_01697_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1789]),
    .QN(_29584_));
 DFF_X1 _63017_ (.D(_01699_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1790]),
    .QN(_29585_));
 DFF_X1 _63018_ (.D(_01700_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1791]),
    .QN(_29586_));
 DFF_X1 _63019_ (.D(_01701_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1792]),
    .QN(_29587_));
 DFF_X1 _63020_ (.D(_01702_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1793]),
    .QN(_29588_));
 DFF_X1 _63021_ (.D(_01703_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1794]),
    .QN(_29589_));
 DFF_X1 _63022_ (.D(_01704_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1795]),
    .QN(_29590_));
 DFF_X1 _63023_ (.D(_01705_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1796]),
    .QN(_29591_));
 DFF_X1 _63024_ (.D(_01706_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1797]),
    .QN(_29592_));
 DFF_X1 _63025_ (.D(_01707_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1798]),
    .QN(_29593_));
 DFF_X1 _63026_ (.D(_01708_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1799]),
    .QN(_29594_));
 DFF_X1 _63027_ (.D(_01711_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1800]),
    .QN(_29595_));
 DFF_X1 _63028_ (.D(_01712_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1801]),
    .QN(_29596_));
 DFF_X1 _63029_ (.D(_01713_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1802]),
    .QN(_29597_));
 DFF_X1 _63030_ (.D(_01714_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1803]),
    .QN(_29598_));
 DFF_X1 _63031_ (.D(_01715_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1804]),
    .QN(_29599_));
 DFF_X1 _63032_ (.D(_01716_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1805]),
    .QN(_29600_));
 DFF_X1 _63033_ (.D(_01717_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1806]),
    .QN(_29601_));
 DFF_X1 _63034_ (.D(_01718_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1807]),
    .QN(_29602_));
 DFF_X1 _63035_ (.D(_01719_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1808]),
    .QN(_29603_));
 DFF_X1 _63036_ (.D(_01720_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1809]),
    .QN(_29604_));
 DFF_X1 _63037_ (.D(_01722_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1810]),
    .QN(_29605_));
 DFF_X1 _63038_ (.D(_01723_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1811]),
    .QN(_29606_));
 DFF_X1 _63039_ (.D(_01724_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1812]),
    .QN(_29607_));
 DFF_X1 _63040_ (.D(_01725_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1813]),
    .QN(_29608_));
 DFF_X1 _63041_ (.D(_01726_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1814]),
    .QN(_29609_));
 DFF_X1 _63042_ (.D(_01727_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1815]),
    .QN(_29610_));
 DFF_X1 _63043_ (.D(_01728_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1816]),
    .QN(_29611_));
 DFF_X1 _63044_ (.D(_01729_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1817]),
    .QN(_29612_));
 DFF_X1 _63045_ (.D(_01730_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1818]),
    .QN(_29613_));
 DFF_X1 _63046_ (.D(_01731_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1819]),
    .QN(_29614_));
 DFF_X1 _63047_ (.D(_01733_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1820]),
    .QN(_29615_));
 DFF_X1 _63048_ (.D(_01734_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1821]),
    .QN(_29616_));
 DFF_X1 _63049_ (.D(_01735_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1822]),
    .QN(_29617_));
 DFF_X1 _63050_ (.D(_01736_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1823]),
    .QN(_29618_));
 DFF_X1 _63051_ (.D(_01737_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1824]),
    .QN(_29619_));
 DFF_X1 _63052_ (.D(_01738_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1825]),
    .QN(_29620_));
 DFF_X1 _63053_ (.D(_01739_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1826]),
    .QN(_29621_));
 DFF_X1 _63054_ (.D(_01740_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1827]),
    .QN(_29622_));
 DFF_X1 _63055_ (.D(_01741_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1828]),
    .QN(_29623_));
 DFF_X1 _63056_ (.D(_01742_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1829]),
    .QN(_29624_));
 DFF_X1 _63057_ (.D(_01744_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1830]),
    .QN(_29625_));
 DFF_X1 _63058_ (.D(_01745_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1831]),
    .QN(_29626_));
 DFF_X1 _63059_ (.D(_01746_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1832]),
    .QN(_29627_));
 DFF_X1 _63060_ (.D(_01747_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1833]),
    .QN(_29628_));
 DFF_X1 _63061_ (.D(_01748_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1834]),
    .QN(_29629_));
 DFF_X1 _63062_ (.D(_01749_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1835]),
    .QN(_29630_));
 DFF_X1 _63063_ (.D(_01750_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1836]),
    .QN(_29631_));
 DFF_X1 _63064_ (.D(_01751_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1837]),
    .QN(_29632_));
 DFF_X1 _63065_ (.D(_01752_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1838]),
    .QN(_29633_));
 DFF_X1 _63066_ (.D(_01753_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1839]),
    .QN(_29634_));
 DFF_X1 _63067_ (.D(_01755_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1840]),
    .QN(_29635_));
 DFF_X1 _63068_ (.D(_01756_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1841]),
    .QN(_29636_));
 DFF_X1 _63069_ (.D(_01757_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1842]),
    .QN(_29637_));
 DFF_X1 _63070_ (.D(_01758_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1843]),
    .QN(_29638_));
 DFF_X1 _63071_ (.D(_01759_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1844]),
    .QN(_29639_));
 DFF_X1 _63072_ (.D(_01760_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1845]),
    .QN(_29640_));
 DFF_X1 _63073_ (.D(_01761_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1846]),
    .QN(_29641_));
 DFF_X1 _63074_ (.D(_01762_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1847]),
    .QN(_29642_));
 DFF_X1 _63075_ (.D(_01763_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1848]),
    .QN(_29643_));
 DFF_X1 _63076_ (.D(_01764_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1849]),
    .QN(_29644_));
 DFF_X1 _63077_ (.D(_01766_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1850]),
    .QN(_29645_));
 DFF_X1 _63078_ (.D(_01767_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1851]),
    .QN(_29646_));
 DFF_X1 _63079_ (.D(_01768_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1852]),
    .QN(_29647_));
 DFF_X1 _63080_ (.D(_01769_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1853]),
    .QN(_29648_));
 DFF_X1 _63081_ (.D(_01770_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1854]),
    .QN(_29649_));
 DFF_X1 _63082_ (.D(_01771_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1855]),
    .QN(_29650_));
 DFF_X1 _63083_ (.D(_01772_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1856]),
    .QN(_29651_));
 DFF_X1 _63084_ (.D(_01773_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1857]),
    .QN(_29652_));
 DFF_X1 _63085_ (.D(_01774_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1858]),
    .QN(_29653_));
 DFF_X1 _63086_ (.D(_01775_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1859]),
    .QN(_29654_));
 DFF_X1 _63087_ (.D(_01777_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1860]),
    .QN(_29655_));
 DFF_X1 _63088_ (.D(_01778_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1861]),
    .QN(_29656_));
 DFF_X1 _63089_ (.D(_01779_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1862]),
    .QN(_29657_));
 DFF_X1 _63090_ (.D(_01780_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1863]),
    .QN(_29658_));
 DFF_X1 _63091_ (.D(_01781_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1864]),
    .QN(_29659_));
 DFF_X1 _63092_ (.D(_01782_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1865]),
    .QN(_29660_));
 DFF_X1 _63093_ (.D(_01783_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1866]),
    .QN(_29661_));
 DFF_X1 _63094_ (.D(_01784_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1867]),
    .QN(_29662_));
 DFF_X1 _63095_ (.D(_01785_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1868]),
    .QN(_29663_));
 DFF_X1 _63096_ (.D(_01786_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1869]),
    .QN(_29664_));
 DFF_X1 _63097_ (.D(_01788_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1870]),
    .QN(_29665_));
 DFF_X1 _63098_ (.D(_01789_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1871]),
    .QN(_29666_));
 DFF_X1 _63099_ (.D(_01790_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1872]),
    .QN(_29667_));
 DFF_X1 _63100_ (.D(_01791_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1873]),
    .QN(_29668_));
 DFF_X1 _63101_ (.D(_01792_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1874]),
    .QN(_29669_));
 DFF_X1 _63102_ (.D(_01793_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1875]),
    .QN(_29670_));
 DFF_X1 _63103_ (.D(_01794_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1876]),
    .QN(_29671_));
 DFF_X1 _63104_ (.D(_01795_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1877]),
    .QN(_29672_));
 DFF_X1 _63105_ (.D(_01796_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1878]),
    .QN(_29673_));
 DFF_X1 _63106_ (.D(_01797_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1879]),
    .QN(_29674_));
 DFF_X1 _63107_ (.D(_01799_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1880]),
    .QN(_29675_));
 DFF_X1 _63108_ (.D(_01800_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1881]),
    .QN(_29676_));
 DFF_X1 _63109_ (.D(_01801_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1882]),
    .QN(_29677_));
 DFF_X1 _63110_ (.D(_01802_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1883]),
    .QN(_29678_));
 DFF_X1 _63111_ (.D(_01803_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1884]),
    .QN(_29679_));
 DFF_X1 _63112_ (.D(_01804_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1885]),
    .QN(_29680_));
 DFF_X1 _63113_ (.D(_01805_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1886]),
    .QN(_29681_));
 DFF_X1 _63114_ (.D(_01806_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1887]),
    .QN(_29682_));
 DFF_X1 _63115_ (.D(_01807_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1888]),
    .QN(_29683_));
 DFF_X1 _63116_ (.D(_01808_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1889]),
    .QN(_29684_));
 DFF_X1 _63117_ (.D(_01810_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1890]),
    .QN(_29685_));
 DFF_X1 _63118_ (.D(_01811_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1891]),
    .QN(_29686_));
 DFF_X1 _63119_ (.D(_01812_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1892]),
    .QN(_29687_));
 DFF_X1 _63120_ (.D(_01813_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1893]),
    .QN(_29688_));
 DFF_X1 _63121_ (.D(_01814_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1894]),
    .QN(_29689_));
 DFF_X1 _63122_ (.D(_01815_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1895]),
    .QN(_29690_));
 DFF_X1 _63123_ (.D(_01816_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1896]),
    .QN(_29691_));
 DFF_X1 _63124_ (.D(_01817_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1897]),
    .QN(_29692_));
 DFF_X1 _63125_ (.D(_01818_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1898]),
    .QN(_29693_));
 DFF_X1 _63126_ (.D(_01819_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1899]),
    .QN(_29694_));
 DFF_X1 _63127_ (.D(_01822_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1900]),
    .QN(_29695_));
 DFF_X1 _63128_ (.D(_01823_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1901]),
    .QN(_29696_));
 DFF_X1 _63129_ (.D(_01824_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1902]),
    .QN(_29697_));
 DFF_X1 _63130_ (.D(_01825_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1903]),
    .QN(_29698_));
 DFF_X1 _63131_ (.D(_01826_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1904]),
    .QN(_29699_));
 DFF_X1 _63132_ (.D(_01827_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1905]),
    .QN(_29700_));
 DFF_X1 _63133_ (.D(_01828_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1906]),
    .QN(_29701_));
 DFF_X1 _63134_ (.D(_01829_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1907]),
    .QN(_29702_));
 DFF_X1 _63135_ (.D(_01830_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1908]),
    .QN(_29703_));
 DFF_X1 _63136_ (.D(_01831_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1909]),
    .QN(_29704_));
 DFF_X1 _63137_ (.D(_01833_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1910]),
    .QN(_29705_));
 DFF_X1 _63138_ (.D(_01834_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1911]),
    .QN(_29706_));
 DFF_X1 _63139_ (.D(_01835_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1912]),
    .QN(_29707_));
 DFF_X1 _63140_ (.D(_01836_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1913]),
    .QN(_29708_));
 DFF_X1 _63141_ (.D(_01837_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1914]),
    .QN(_29709_));
 DFF_X1 _63142_ (.D(_01838_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1915]),
    .QN(_29710_));
 DFF_X1 _63143_ (.D(_01839_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1916]),
    .QN(_29711_));
 DFF_X1 _63144_ (.D(_01840_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1917]),
    .QN(_29712_));
 DFF_X1 _63145_ (.D(_01841_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1918]),
    .QN(_29713_));
 DFF_X1 _63146_ (.D(_01842_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1919]),
    .QN(_29714_));
 DFF_X1 _63147_ (.D(_01844_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1920]),
    .QN(_29715_));
 DFF_X1 _63148_ (.D(_01845_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1921]),
    .QN(_29716_));
 DFF_X1 _63149_ (.D(_01846_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1922]),
    .QN(_29717_));
 DFF_X1 _63150_ (.D(_01847_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1923]),
    .QN(_29718_));
 DFF_X1 _63151_ (.D(_01848_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1924]),
    .QN(_29719_));
 DFF_X1 _63152_ (.D(_01849_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1925]),
    .QN(_29720_));
 DFF_X1 _63153_ (.D(_01850_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1926]),
    .QN(_29721_));
 DFF_X1 _63154_ (.D(_01851_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1927]),
    .QN(_29722_));
 DFF_X1 _63155_ (.D(_01852_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1928]),
    .QN(_29723_));
 DFF_X1 _63156_ (.D(_01853_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1929]),
    .QN(_29724_));
 DFF_X1 _63157_ (.D(_01855_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1930]),
    .QN(_29725_));
 DFF_X1 _63158_ (.D(_01856_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1931]),
    .QN(_29726_));
 DFF_X1 _63159_ (.D(_01857_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1932]),
    .QN(_29727_));
 DFF_X1 _63160_ (.D(_01858_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1933]),
    .QN(_29728_));
 DFF_X1 _63161_ (.D(_01859_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1934]),
    .QN(_29729_));
 DFF_X1 _63162_ (.D(_01860_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1935]),
    .QN(_29730_));
 DFF_X1 _63163_ (.D(_01861_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1936]),
    .QN(_29731_));
 DFF_X1 _63164_ (.D(_01862_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1937]),
    .QN(_29732_));
 DFF_X1 _63165_ (.D(_01863_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1938]),
    .QN(_29733_));
 DFF_X1 _63166_ (.D(_01864_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1939]),
    .QN(_29734_));
 DFF_X1 _63167_ (.D(_01866_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1940]),
    .QN(_29735_));
 DFF_X1 _63168_ (.D(_01867_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1941]),
    .QN(_29736_));
 DFF_X1 _63169_ (.D(_01868_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1942]),
    .QN(_29737_));
 DFF_X1 _63170_ (.D(_01869_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1943]),
    .QN(_29738_));
 DFF_X1 _63171_ (.D(_01870_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1944]),
    .QN(_29739_));
 DFF_X1 _63172_ (.D(_01871_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1945]),
    .QN(_29740_));
 DFF_X1 _63173_ (.D(_01872_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1946]),
    .QN(_29741_));
 DFF_X1 _63174_ (.D(_01873_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1947]),
    .QN(_29742_));
 DFF_X1 _63175_ (.D(_01874_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1948]),
    .QN(_29743_));
 DFF_X1 _63176_ (.D(_01875_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1949]),
    .QN(_29744_));
 DFF_X1 _63177_ (.D(_01877_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1950]),
    .QN(_29745_));
 DFF_X1 _63178_ (.D(_01878_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1951]),
    .QN(_29746_));
 DFF_X1 _63179_ (.D(_01879_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1952]),
    .QN(_29747_));
 DFF_X1 _63180_ (.D(_01880_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1953]),
    .QN(_29748_));
 DFF_X1 _63181_ (.D(_01881_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1954]),
    .QN(_29749_));
 DFF_X1 _63182_ (.D(_01882_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1955]),
    .QN(_29750_));
 DFF_X1 _63183_ (.D(_01883_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1956]),
    .QN(_29751_));
 DFF_X1 _63184_ (.D(_01884_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1957]),
    .QN(_29752_));
 DFF_X1 _63185_ (.D(_01885_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1958]),
    .QN(_29753_));
 DFF_X1 _63186_ (.D(_01886_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1959]),
    .QN(_29754_));
 DFF_X1 _63187_ (.D(_01888_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1960]),
    .QN(_29755_));
 DFF_X1 _63188_ (.D(_01889_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1961]),
    .QN(_29756_));
 DFF_X1 _63189_ (.D(_01890_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1962]),
    .QN(_29757_));
 DFF_X1 _63190_ (.D(_01891_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1963]),
    .QN(_29758_));
 DFF_X1 _63191_ (.D(_01892_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1964]),
    .QN(_29759_));
 DFF_X1 _63192_ (.D(_01893_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1965]),
    .QN(_29760_));
 DFF_X1 _63193_ (.D(_01894_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1966]),
    .QN(_29761_));
 DFF_X1 _63194_ (.D(_01895_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1967]),
    .QN(_29762_));
 DFF_X1 _63195_ (.D(_01896_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1968]),
    .QN(_29763_));
 DFF_X1 _63196_ (.D(_01897_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1969]),
    .QN(_29764_));
 DFF_X1 _63197_ (.D(_01899_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1970]),
    .QN(_29765_));
 DFF_X1 _63198_ (.D(_01900_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1971]),
    .QN(_29766_));
 DFF_X1 _63199_ (.D(_01901_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1972]),
    .QN(_29767_));
 DFF_X1 _63200_ (.D(_01902_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1973]),
    .QN(_29768_));
 DFF_X1 _63201_ (.D(_01903_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1974]),
    .QN(_29769_));
 DFF_X1 _63202_ (.D(_01904_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1975]),
    .QN(_29770_));
 DFF_X1 _63203_ (.D(_01905_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1976]),
    .QN(_29771_));
 DFF_X1 _63204_ (.D(_01906_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1977]),
    .QN(_29772_));
 DFF_X1 _63205_ (.D(_01907_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1978]),
    .QN(_29773_));
 DFF_X1 _63206_ (.D(_01908_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1979]),
    .QN(_29774_));
 DFF_X1 _63207_ (.D(_01910_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1980]),
    .QN(_29775_));
 DFF_X1 _63208_ (.D(_01911_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1981]),
    .QN(_29776_));
 DFF_X1 _63209_ (.D(_01912_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1982]),
    .QN(_29777_));
 DFF_X1 _63210_ (.D(_01913_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1983]),
    .QN(_29778_));
 DFF_X1 _63211_ (.D(_01914_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1984]),
    .QN(_29779_));
 DFF_X1 _63212_ (.D(_01915_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1985]),
    .QN(_29780_));
 DFF_X1 _63213_ (.D(_01916_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1986]),
    .QN(_29781_));
 DFF_X1 _63214_ (.D(_01917_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1987]),
    .QN(_29782_));
 DFF_X1 _63215_ (.D(_01918_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1988]),
    .QN(_29783_));
 DFF_X1 _63216_ (.D(_01919_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1989]),
    .QN(_29784_));
 DFF_X1 _63217_ (.D(_01921_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1990]),
    .QN(_29785_));
 DFF_X1 _63218_ (.D(_01922_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1991]),
    .QN(_29786_));
 DFF_X1 _63219_ (.D(_01923_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1992]),
    .QN(_29787_));
 DFF_X1 _63220_ (.D(_01924_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1993]),
    .QN(_29788_));
 DFF_X1 _63221_ (.D(_01925_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1994]),
    .QN(_29789_));
 DFF_X1 _63222_ (.D(_01926_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1995]),
    .QN(_29790_));
 DFF_X1 _63223_ (.D(_01927_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1996]),
    .QN(_29791_));
 DFF_X1 _63224_ (.D(_01928_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1997]),
    .QN(_29792_));
 DFF_X1 _63225_ (.D(_01929_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1998]),
    .QN(_29793_));
 DFF_X1 _63226_ (.D(_01930_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [1999]),
    .QN(_29794_));
 DFF_X1 _63227_ (.D(_01934_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2000]),
    .QN(_29795_));
 DFF_X1 _63228_ (.D(_01935_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2001]),
    .QN(_29796_));
 DFF_X1 _63229_ (.D(_01936_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2002]),
    .QN(_29797_));
 DFF_X1 _63230_ (.D(_01937_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2003]),
    .QN(_29798_));
 DFF_X1 _63231_ (.D(_01938_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2004]),
    .QN(_29799_));
 DFF_X1 _63232_ (.D(_01939_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2005]),
    .QN(_29800_));
 DFF_X1 _63233_ (.D(_01940_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2006]),
    .QN(_29801_));
 DFF_X1 _63234_ (.D(_01941_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2007]),
    .QN(_29802_));
 DFF_X1 _63235_ (.D(_01942_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2008]),
    .QN(_29803_));
 DFF_X1 _63236_ (.D(_01943_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2009]),
    .QN(_29804_));
 DFF_X1 _63237_ (.D(_01945_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2010]),
    .QN(_29805_));
 DFF_X1 _63238_ (.D(_01946_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2011]),
    .QN(_29806_));
 DFF_X1 _63239_ (.D(_01947_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2012]),
    .QN(_29807_));
 DFF_X1 _63240_ (.D(_01948_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2013]),
    .QN(_29808_));
 DFF_X1 _63241_ (.D(_01949_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2014]),
    .QN(_29809_));
 DFF_X1 _63242_ (.D(_01950_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2015]),
    .QN(_29810_));
 DFF_X1 _63243_ (.D(_01951_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2016]),
    .QN(_29811_));
 DFF_X1 _63244_ (.D(_01952_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2017]),
    .QN(_29812_));
 DFF_X1 _63245_ (.D(_01953_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2018]),
    .QN(_29813_));
 DFF_X1 _63246_ (.D(_01954_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2019]),
    .QN(_29814_));
 DFF_X1 _63247_ (.D(_01956_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2020]),
    .QN(_29815_));
 DFF_X1 _63248_ (.D(_01957_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2021]),
    .QN(_29816_));
 DFF_X1 _63249_ (.D(_01958_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2022]),
    .QN(_29817_));
 DFF_X1 _63250_ (.D(_01959_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2023]),
    .QN(_29818_));
 DFF_X1 _63251_ (.D(_01960_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2024]),
    .QN(_29819_));
 DFF_X1 _63252_ (.D(_01961_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2025]),
    .QN(_29820_));
 DFF_X1 _63253_ (.D(_01962_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2026]),
    .QN(_29821_));
 DFF_X1 _63254_ (.D(_01963_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2027]),
    .QN(_29822_));
 DFF_X1 _63255_ (.D(_01964_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2028]),
    .QN(_29823_));
 DFF_X1 _63256_ (.D(_01965_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2029]),
    .QN(_29824_));
 DFF_X1 _63257_ (.D(_01967_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2030]),
    .QN(_29825_));
 DFF_X1 _63258_ (.D(_01968_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2031]),
    .QN(_29826_));
 DFF_X1 _63259_ (.D(_01969_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2032]),
    .QN(_29827_));
 DFF_X1 _63260_ (.D(_01970_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2033]),
    .QN(_29828_));
 DFF_X1 _63261_ (.D(_01971_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2034]),
    .QN(_29829_));
 DFF_X1 _63262_ (.D(_01972_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2035]),
    .QN(_29830_));
 DFF_X1 _63263_ (.D(_01973_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2036]),
    .QN(_29831_));
 DFF_X1 _63264_ (.D(_01974_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2037]),
    .QN(_29832_));
 DFF_X1 _63265_ (.D(_01975_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2038]),
    .QN(_29833_));
 DFF_X1 _63266_ (.D(_01976_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2039]),
    .QN(_29834_));
 DFF_X1 _63267_ (.D(_01978_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2040]),
    .QN(_29835_));
 DFF_X1 _63268_ (.D(_01979_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2041]),
    .QN(_29836_));
 DFF_X1 _63269_ (.D(_01980_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2042]),
    .QN(_29837_));
 DFF_X1 _63270_ (.D(_01981_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2043]),
    .QN(_29838_));
 DFF_X1 _63271_ (.D(_01982_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2044]),
    .QN(_29839_));
 DFF_X1 _63272_ (.D(_01983_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2045]),
    .QN(_29840_));
 DFF_X1 _63273_ (.D(_01984_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2046]),
    .QN(_29841_));
 DFF_X1 _63274_ (.D(_01985_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2047]),
    .QN(_29842_));
 DFF_X1 _63275_ (.D(_01986_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2048]),
    .QN(_29843_));
 DFF_X1 _63276_ (.D(_01987_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2049]),
    .QN(_29844_));
 DFF_X1 _63277_ (.D(_01989_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2050]),
    .QN(_29845_));
 DFF_X1 _63278_ (.D(_01990_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2051]),
    .QN(_29846_));
 DFF_X1 _63279_ (.D(_01991_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2052]),
    .QN(_29847_));
 DFF_X1 _63280_ (.D(_01992_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2053]),
    .QN(_29848_));
 DFF_X1 _63281_ (.D(_01993_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2054]),
    .QN(_29849_));
 DFF_X1 _63282_ (.D(_01994_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2055]),
    .QN(_29850_));
 DFF_X1 _63283_ (.D(_01995_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2056]),
    .QN(_29851_));
 DFF_X1 _63284_ (.D(_01996_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2057]),
    .QN(_29852_));
 DFF_X1 _63285_ (.D(_01997_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2058]),
    .QN(_29853_));
 DFF_X1 _63286_ (.D(_01998_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2059]),
    .QN(_29854_));
 DFF_X1 _63287_ (.D(_02000_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2060]),
    .QN(_29855_));
 DFF_X1 _63288_ (.D(_02001_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2061]),
    .QN(_29856_));
 DFF_X1 _63289_ (.D(_02002_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2062]),
    .QN(_29857_));
 DFF_X1 _63290_ (.D(_02003_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2063]),
    .QN(_29858_));
 DFF_X1 _63291_ (.D(_02004_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2064]),
    .QN(_29859_));
 DFF_X1 _63292_ (.D(_02005_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2065]),
    .QN(_29860_));
 DFF_X1 _63293_ (.D(_02006_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2066]),
    .QN(_29861_));
 DFF_X1 _63294_ (.D(_02007_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2067]),
    .QN(_29862_));
 DFF_X1 _63295_ (.D(_02008_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2068]),
    .QN(_29863_));
 DFF_X1 _63296_ (.D(_02009_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2069]),
    .QN(_29864_));
 DFF_X1 _63297_ (.D(_02011_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2070]),
    .QN(_29865_));
 DFF_X1 _63298_ (.D(_02012_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2071]),
    .QN(_29866_));
 DFF_X1 _63299_ (.D(_02013_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2072]),
    .QN(_29867_));
 DFF_X1 _63300_ (.D(_02014_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2073]),
    .QN(_29868_));
 DFF_X1 _63301_ (.D(_02015_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2074]),
    .QN(_29869_));
 DFF_X1 _63302_ (.D(_02016_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2075]),
    .QN(_29870_));
 DFF_X1 _63303_ (.D(_02017_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2076]),
    .QN(_29871_));
 DFF_X1 _63304_ (.D(_02018_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2077]),
    .QN(_29872_));
 DFF_X1 _63305_ (.D(_02019_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2078]),
    .QN(_29873_));
 DFF_X1 _63306_ (.D(_02020_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2079]),
    .QN(_29874_));
 DFF_X1 _63307_ (.D(_02022_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2080]),
    .QN(_29875_));
 DFF_X1 _63308_ (.D(_02023_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2081]),
    .QN(_29876_));
 DFF_X1 _63309_ (.D(_02024_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2082]),
    .QN(_29877_));
 DFF_X1 _63310_ (.D(_02025_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2083]),
    .QN(_29878_));
 DFF_X1 _63311_ (.D(_02026_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2084]),
    .QN(_29879_));
 DFF_X1 _63312_ (.D(_02027_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2085]),
    .QN(_29880_));
 DFF_X1 _63313_ (.D(_02028_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2086]),
    .QN(_29881_));
 DFF_X1 _63314_ (.D(_02029_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2087]),
    .QN(_29882_));
 DFF_X1 _63315_ (.D(_02030_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2088]),
    .QN(_29883_));
 DFF_X1 _63316_ (.D(_02031_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2089]),
    .QN(_29884_));
 DFF_X1 _63317_ (.D(_02033_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2090]),
    .QN(_29885_));
 DFF_X1 _63318_ (.D(_02034_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2091]),
    .QN(_29886_));
 DFF_X1 _63319_ (.D(_02035_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2092]),
    .QN(_29887_));
 DFF_X1 _63320_ (.D(_02036_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2093]),
    .QN(_29888_));
 DFF_X1 _63321_ (.D(_02037_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2094]),
    .QN(_29889_));
 DFF_X1 _63322_ (.D(_02038_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2095]),
    .QN(_29890_));
 DFF_X1 _63323_ (.D(_02039_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2096]),
    .QN(_29891_));
 DFF_X1 _63324_ (.D(_02040_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2097]),
    .QN(_29892_));
 DFF_X1 _63325_ (.D(_02041_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2098]),
    .QN(_29893_));
 DFF_X1 _63326_ (.D(_02042_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2099]),
    .QN(_29894_));
 DFF_X1 _63327_ (.D(_02045_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2100]),
    .QN(_29895_));
 DFF_X1 _63328_ (.D(_02046_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2101]),
    .QN(_29896_));
 DFF_X1 _63329_ (.D(_02047_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2102]),
    .QN(_29897_));
 DFF_X1 _63330_ (.D(_02048_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2103]),
    .QN(_29898_));
 DFF_X1 _63331_ (.D(_02049_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2104]),
    .QN(_29899_));
 DFF_X1 _63332_ (.D(_02050_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2105]),
    .QN(_29900_));
 DFF_X1 _63333_ (.D(_02051_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2106]),
    .QN(_29901_));
 DFF_X1 _63334_ (.D(_02052_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2107]),
    .QN(_29902_));
 DFF_X1 _63335_ (.D(_02053_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2108]),
    .QN(_29903_));
 DFF_X1 _63336_ (.D(_02054_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2109]),
    .QN(_29904_));
 DFF_X1 _63337_ (.D(_02056_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2110]),
    .QN(_29905_));
 DFF_X1 _63338_ (.D(_02057_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2111]),
    .QN(_29906_));
 DFF_X1 _63339_ (.D(_02058_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2112]),
    .QN(_29907_));
 DFF_X1 _63340_ (.D(_02059_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2113]),
    .QN(_29908_));
 DFF_X1 _63341_ (.D(_02060_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2114]),
    .QN(_29909_));
 DFF_X1 _63342_ (.D(_02061_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2115]),
    .QN(_29910_));
 DFF_X1 _63343_ (.D(_02062_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2116]),
    .QN(_29911_));
 DFF_X1 _63344_ (.D(_02063_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2117]),
    .QN(_29912_));
 DFF_X1 _63345_ (.D(_02064_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2118]),
    .QN(_29913_));
 DFF_X1 _63346_ (.D(_02065_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2119]),
    .QN(_29914_));
 DFF_X1 _63347_ (.D(_02067_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2120]),
    .QN(_29915_));
 DFF_X1 _63348_ (.D(_02068_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2121]),
    .QN(_29916_));
 DFF_X1 _63349_ (.D(_02069_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2122]),
    .QN(_29917_));
 DFF_X1 _63350_ (.D(_02070_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2123]),
    .QN(_29918_));
 DFF_X1 _63351_ (.D(_02071_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2124]),
    .QN(_29919_));
 DFF_X1 _63352_ (.D(_02072_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2125]),
    .QN(_29920_));
 DFF_X1 _63353_ (.D(_02073_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2126]),
    .QN(_29921_));
 DFF_X1 _63354_ (.D(_02074_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2127]),
    .QN(_29922_));
 DFF_X1 _63355_ (.D(_02075_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2128]),
    .QN(_29923_));
 DFF_X1 _63356_ (.D(_02076_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2129]),
    .QN(_29924_));
 DFF_X1 _63357_ (.D(_02078_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2130]),
    .QN(_29925_));
 DFF_X1 _63358_ (.D(_02079_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2131]),
    .QN(_29926_));
 DFF_X1 _63359_ (.D(_02080_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2132]),
    .QN(_29927_));
 DFF_X1 _63360_ (.D(_02081_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2133]),
    .QN(_29928_));
 DFF_X1 _63361_ (.D(_02082_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2134]),
    .QN(_29929_));
 DFF_X1 _63362_ (.D(_02083_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2135]),
    .QN(_29930_));
 DFF_X1 _63363_ (.D(_02084_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2136]),
    .QN(_29931_));
 DFF_X1 _63364_ (.D(_02085_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2137]),
    .QN(_29932_));
 DFF_X1 _63365_ (.D(_02086_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2138]),
    .QN(_29933_));
 DFF_X1 _63366_ (.D(_02087_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2139]),
    .QN(_29934_));
 DFF_X1 _63367_ (.D(_02089_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2140]),
    .QN(_29935_));
 DFF_X1 _63368_ (.D(_02090_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2141]),
    .QN(_29936_));
 DFF_X1 _63369_ (.D(_02091_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2142]),
    .QN(_29937_));
 DFF_X1 _63370_ (.D(_02092_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2143]),
    .QN(_29938_));
 DFF_X1 _63371_ (.D(_02093_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2144]),
    .QN(_29939_));
 DFF_X1 _63372_ (.D(_02094_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2145]),
    .QN(_29940_));
 DFF_X1 _63373_ (.D(_02095_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2146]),
    .QN(_29941_));
 DFF_X1 _63374_ (.D(_02096_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2147]),
    .QN(_29942_));
 DFF_X1 _63375_ (.D(_02097_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2148]),
    .QN(_29943_));
 DFF_X1 _63376_ (.D(_02098_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2149]),
    .QN(_29944_));
 DFF_X1 _63377_ (.D(_02100_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2150]),
    .QN(_29945_));
 DFF_X1 _63378_ (.D(_02101_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2151]),
    .QN(_29946_));
 DFF_X1 _63379_ (.D(_02102_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2152]),
    .QN(_29947_));
 DFF_X1 _63380_ (.D(_02103_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2153]),
    .QN(_29948_));
 DFF_X1 _63381_ (.D(_02104_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2154]),
    .QN(_29949_));
 DFF_X1 _63382_ (.D(_02105_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2155]),
    .QN(_29950_));
 DFF_X1 _63383_ (.D(_02106_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2156]),
    .QN(_29951_));
 DFF_X1 _63384_ (.D(_02107_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2157]),
    .QN(_29952_));
 DFF_X1 _63385_ (.D(_02108_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2158]),
    .QN(_29953_));
 DFF_X1 _63386_ (.D(_02109_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2159]),
    .QN(_29954_));
 DFF_X1 _63387_ (.D(_02111_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2160]),
    .QN(_29955_));
 DFF_X1 _63388_ (.D(_02112_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2161]),
    .QN(_29956_));
 DFF_X1 _63389_ (.D(_02113_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2162]),
    .QN(_29957_));
 DFF_X1 _63390_ (.D(_02114_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2163]),
    .QN(_29958_));
 DFF_X1 _63391_ (.D(_02115_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2164]),
    .QN(_29959_));
 DFF_X1 _63392_ (.D(_02116_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2165]),
    .QN(_29960_));
 DFF_X1 _63393_ (.D(_02117_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2166]),
    .QN(_29961_));
 DFF_X1 _63394_ (.D(_02118_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2167]),
    .QN(_29962_));
 DFF_X1 _63395_ (.D(_02119_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2168]),
    .QN(_29963_));
 DFF_X1 _63396_ (.D(_02120_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2169]),
    .QN(_29964_));
 DFF_X1 _63397_ (.D(_02122_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2170]),
    .QN(_29965_));
 DFF_X1 _63398_ (.D(_02123_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2171]),
    .QN(_29966_));
 DFF_X1 _63399_ (.D(_02124_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2172]),
    .QN(_29967_));
 DFF_X1 _63400_ (.D(_02125_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2173]),
    .QN(_29968_));
 DFF_X1 _63401_ (.D(_02126_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2174]),
    .QN(_29969_));
 DFF_X1 _63402_ (.D(_02127_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2175]),
    .QN(_29970_));
 DFF_X1 _63403_ (.D(_02128_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2176]),
    .QN(_29971_));
 DFF_X1 _63404_ (.D(_02129_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2177]),
    .QN(_29972_));
 DFF_X1 _63405_ (.D(_02130_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2178]),
    .QN(_29973_));
 DFF_X1 _63406_ (.D(_02131_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2179]),
    .QN(_29974_));
 DFF_X1 _63407_ (.D(_02133_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2180]),
    .QN(_29975_));
 DFF_X1 _63408_ (.D(_02134_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2181]),
    .QN(_29976_));
 DFF_X1 _63409_ (.D(_02135_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2182]),
    .QN(_29977_));
 DFF_X1 _63410_ (.D(_02136_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2183]),
    .QN(_29978_));
 DFF_X1 _63411_ (.D(_02137_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2184]),
    .QN(_29979_));
 DFF_X1 _63412_ (.D(_02138_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2185]),
    .QN(_29980_));
 DFF_X1 _63413_ (.D(_02139_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2186]),
    .QN(_29981_));
 DFF_X1 _63414_ (.D(_02140_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2187]),
    .QN(_29982_));
 DFF_X1 _63415_ (.D(_02141_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2188]),
    .QN(_29983_));
 DFF_X1 _63416_ (.D(_02142_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2189]),
    .QN(_29984_));
 DFF_X1 _63417_ (.D(_02144_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2190]),
    .QN(_29985_));
 DFF_X1 _63418_ (.D(_02145_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2191]),
    .QN(_29986_));
 DFF_X1 _63419_ (.D(_02146_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2192]),
    .QN(_29987_));
 DFF_X1 _63420_ (.D(_02147_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2193]),
    .QN(_29988_));
 DFF_X1 _63421_ (.D(_02148_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2194]),
    .QN(_29989_));
 DFF_X1 _63422_ (.D(_02149_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2195]),
    .QN(_29990_));
 DFF_X1 _63423_ (.D(_02150_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2196]),
    .QN(_29991_));
 DFF_X1 _63424_ (.D(_02151_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2197]),
    .QN(_29992_));
 DFF_X1 _63425_ (.D(_02152_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2198]),
    .QN(_29993_));
 DFF_X1 _63426_ (.D(_02153_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2199]),
    .QN(_29994_));
 DFF_X1 _63427_ (.D(_02156_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2200]),
    .QN(_29995_));
 DFF_X1 _63428_ (.D(_02157_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2201]),
    .QN(_29996_));
 DFF_X1 _63429_ (.D(_02158_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2202]),
    .QN(_29997_));
 DFF_X1 _63430_ (.D(_02159_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2203]),
    .QN(_29998_));
 DFF_X1 _63431_ (.D(_02160_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2204]),
    .QN(_29999_));
 DFF_X1 _63432_ (.D(_02161_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2205]),
    .QN(_30000_));
 DFF_X1 _63433_ (.D(_02162_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2206]),
    .QN(_30001_));
 DFF_X1 _63434_ (.D(_02163_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2207]),
    .QN(_30002_));
 DFF_X1 _63435_ (.D(_02164_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2208]),
    .QN(_30003_));
 DFF_X1 _63436_ (.D(_02165_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2209]),
    .QN(_30004_));
 DFF_X1 _63437_ (.D(_02167_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2210]),
    .QN(_30005_));
 DFF_X1 _63438_ (.D(_02168_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2211]),
    .QN(_30006_));
 DFF_X1 _63439_ (.D(_02169_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2212]),
    .QN(_30007_));
 DFF_X1 _63440_ (.D(_02170_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2213]),
    .QN(_30008_));
 DFF_X1 _63441_ (.D(_02171_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2214]),
    .QN(_30009_));
 DFF_X1 _63442_ (.D(_02172_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2215]),
    .QN(_30010_));
 DFF_X1 _63443_ (.D(_02173_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2216]),
    .QN(_30011_));
 DFF_X1 _63444_ (.D(_02174_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2217]),
    .QN(_30012_));
 DFF_X1 _63445_ (.D(_02175_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2218]),
    .QN(_30013_));
 DFF_X1 _63446_ (.D(_02176_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2219]),
    .QN(_30014_));
 DFF_X1 _63447_ (.D(_02178_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2220]),
    .QN(_30015_));
 DFF_X1 _63448_ (.D(_02179_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2221]),
    .QN(_30016_));
 DFF_X1 _63449_ (.D(_02180_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2222]),
    .QN(_30017_));
 DFF_X1 _63450_ (.D(_02181_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2223]),
    .QN(_30018_));
 DFF_X1 _63451_ (.D(_02182_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2224]),
    .QN(_30019_));
 DFF_X1 _63452_ (.D(_02183_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2225]),
    .QN(_30020_));
 DFF_X1 _63453_ (.D(_02184_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2226]),
    .QN(_30021_));
 DFF_X1 _63454_ (.D(_02185_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2227]),
    .QN(_30022_));
 DFF_X1 _63455_ (.D(_02186_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2228]),
    .QN(_30023_));
 DFF_X1 _63456_ (.D(_02187_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2229]),
    .QN(_30024_));
 DFF_X1 _63457_ (.D(_02189_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2230]),
    .QN(_30025_));
 DFF_X1 _63458_ (.D(_02190_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2231]),
    .QN(_30026_));
 DFF_X1 _63459_ (.D(_02191_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2232]),
    .QN(_30027_));
 DFF_X1 _63460_ (.D(_02192_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2233]),
    .QN(_30028_));
 DFF_X1 _63461_ (.D(_02193_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2234]),
    .QN(_30029_));
 DFF_X1 _63462_ (.D(_02194_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2235]),
    .QN(_30030_));
 DFF_X1 _63463_ (.D(_02195_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2236]),
    .QN(_30031_));
 DFF_X1 _63464_ (.D(_02196_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2237]),
    .QN(_30032_));
 DFF_X1 _63465_ (.D(_02197_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2238]),
    .QN(_30033_));
 DFF_X1 _63466_ (.D(_02198_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2239]),
    .QN(_30034_));
 DFF_X1 _63467_ (.D(_02200_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2240]),
    .QN(_30035_));
 DFF_X1 _63468_ (.D(_02201_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2241]),
    .QN(_30036_));
 DFF_X1 _63469_ (.D(_02202_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2242]),
    .QN(_30037_));
 DFF_X1 _63470_ (.D(_02203_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2243]),
    .QN(_30038_));
 DFF_X1 _63471_ (.D(_02204_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2244]),
    .QN(_30039_));
 DFF_X1 _63472_ (.D(_02205_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2245]),
    .QN(_30040_));
 DFF_X1 _63473_ (.D(_02206_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2246]),
    .QN(_30041_));
 DFF_X1 _63474_ (.D(_02207_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2247]),
    .QN(_30042_));
 DFF_X1 _63475_ (.D(_02208_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2248]),
    .QN(_30043_));
 DFF_X1 _63476_ (.D(_02209_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2249]),
    .QN(_30044_));
 DFF_X1 _63477_ (.D(_02211_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2250]),
    .QN(_30045_));
 DFF_X1 _63478_ (.D(_02212_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2251]),
    .QN(_30046_));
 DFF_X1 _63479_ (.D(_02213_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2252]),
    .QN(_30047_));
 DFF_X1 _63480_ (.D(_02214_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2253]),
    .QN(_30048_));
 DFF_X1 _63481_ (.D(_02215_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2254]),
    .QN(_30049_));
 DFF_X1 _63482_ (.D(_02216_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2255]),
    .QN(_30050_));
 DFF_X1 _63483_ (.D(_02217_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2256]),
    .QN(_30051_));
 DFF_X1 _63484_ (.D(_02218_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2257]),
    .QN(_30052_));
 DFF_X1 _63485_ (.D(_02219_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2258]),
    .QN(_30053_));
 DFF_X1 _63486_ (.D(_02220_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2259]),
    .QN(_30054_));
 DFF_X1 _63487_ (.D(_02222_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2260]),
    .QN(_30055_));
 DFF_X1 _63488_ (.D(_02223_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2261]),
    .QN(_30056_));
 DFF_X1 _63489_ (.D(_02224_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2262]),
    .QN(_30057_));
 DFF_X1 _63490_ (.D(_02225_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2263]),
    .QN(_30058_));
 DFF_X1 _63491_ (.D(_02226_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2264]),
    .QN(_30059_));
 DFF_X1 _63492_ (.D(_02227_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2265]),
    .QN(_30060_));
 DFF_X1 _63493_ (.D(_02228_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2266]),
    .QN(_30061_));
 DFF_X1 _63494_ (.D(_02229_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2267]),
    .QN(_30062_));
 DFF_X1 _63495_ (.D(_02230_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2268]),
    .QN(_30063_));
 DFF_X1 _63496_ (.D(_02231_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2269]),
    .QN(_30064_));
 DFF_X1 _63497_ (.D(_02233_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2270]),
    .QN(_30065_));
 DFF_X1 _63498_ (.D(_02234_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2271]),
    .QN(_30066_));
 DFF_X1 _63499_ (.D(_02235_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2272]),
    .QN(_30067_));
 DFF_X1 _63500_ (.D(_02236_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2273]),
    .QN(_30068_));
 DFF_X1 _63501_ (.D(_02237_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2274]),
    .QN(_30069_));
 DFF_X1 _63502_ (.D(_02238_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2275]),
    .QN(_30070_));
 DFF_X1 _63503_ (.D(_02239_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2276]),
    .QN(_30071_));
 DFF_X1 _63504_ (.D(_02240_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2277]),
    .QN(_30072_));
 DFF_X1 _63505_ (.D(_02241_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2278]),
    .QN(_30073_));
 DFF_X1 _63506_ (.D(_02242_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2279]),
    .QN(_30074_));
 DFF_X1 _63507_ (.D(_02244_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2280]),
    .QN(_30075_));
 DFF_X1 _63508_ (.D(_02245_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2281]),
    .QN(_30076_));
 DFF_X1 _63509_ (.D(_02246_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2282]),
    .QN(_30077_));
 DFF_X1 _63510_ (.D(_02247_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2283]),
    .QN(_30078_));
 DFF_X1 _63511_ (.D(_02248_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2284]),
    .QN(_30079_));
 DFF_X1 _63512_ (.D(_02249_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2285]),
    .QN(_30080_));
 DFF_X1 _63513_ (.D(_02250_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2286]),
    .QN(_30081_));
 DFF_X1 _63514_ (.D(_02251_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2287]),
    .QN(_30082_));
 DFF_X1 _63515_ (.D(_02252_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2288]),
    .QN(_30083_));
 DFF_X1 _63516_ (.D(_02253_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2289]),
    .QN(_30084_));
 DFF_X1 _63517_ (.D(_02255_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2290]),
    .QN(_30085_));
 DFF_X1 _63518_ (.D(_02256_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2291]),
    .QN(_30086_));
 DFF_X1 _63519_ (.D(_02257_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2292]),
    .QN(_30087_));
 DFF_X1 _63520_ (.D(_02258_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2293]),
    .QN(_30088_));
 DFF_X1 _63521_ (.D(_02259_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2294]),
    .QN(_30089_));
 DFF_X1 _63522_ (.D(_02260_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2295]),
    .QN(_30090_));
 DFF_X1 _63523_ (.D(_02261_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2296]),
    .QN(_30091_));
 DFF_X1 _63524_ (.D(_02262_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2297]),
    .QN(_30092_));
 DFF_X1 _63525_ (.D(_02263_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2298]),
    .QN(_30093_));
 DFF_X1 _63526_ (.D(_02264_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2299]),
    .QN(_30094_));
 DFF_X1 _63527_ (.D(_02267_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2300]),
    .QN(_30095_));
 DFF_X1 _63528_ (.D(_02268_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2301]),
    .QN(_30096_));
 DFF_X1 _63529_ (.D(_02269_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2302]),
    .QN(_30097_));
 DFF_X1 _63530_ (.D(_02270_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2303]),
    .QN(_30098_));
 DFF_X1 _63531_ (.D(_02271_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2304]),
    .QN(_30099_));
 DFF_X1 _63532_ (.D(_02272_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2305]),
    .QN(_30100_));
 DFF_X1 _63533_ (.D(_02273_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2306]),
    .QN(_30101_));
 DFF_X1 _63534_ (.D(_02274_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2307]),
    .QN(_30102_));
 DFF_X1 _63535_ (.D(_02275_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2308]),
    .QN(_30103_));
 DFF_X1 _63536_ (.D(_02276_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2309]),
    .QN(_30104_));
 DFF_X1 _63537_ (.D(_02278_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2310]),
    .QN(_30105_));
 DFF_X1 _63538_ (.D(_02279_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2311]),
    .QN(_30106_));
 DFF_X1 _63539_ (.D(_02280_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2312]),
    .QN(_30107_));
 DFF_X1 _63540_ (.D(_02281_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2313]),
    .QN(_30108_));
 DFF_X1 _63541_ (.D(_02282_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2314]),
    .QN(_30109_));
 DFF_X1 _63542_ (.D(_02283_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2315]),
    .QN(_30110_));
 DFF_X1 _63543_ (.D(_02284_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2316]),
    .QN(_30111_));
 DFF_X1 _63544_ (.D(_02285_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2317]),
    .QN(_30112_));
 DFF_X1 _63545_ (.D(_02286_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2318]),
    .QN(_30113_));
 DFF_X1 _63546_ (.D(_02287_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2319]),
    .QN(_30114_));
 DFF_X1 _63547_ (.D(_02289_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2320]),
    .QN(_30115_));
 DFF_X1 _63548_ (.D(_02290_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2321]),
    .QN(_30116_));
 DFF_X1 _63549_ (.D(_02291_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2322]),
    .QN(_30117_));
 DFF_X1 _63550_ (.D(_02292_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2323]),
    .QN(_30118_));
 DFF_X1 _63551_ (.D(_02293_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2324]),
    .QN(_30119_));
 DFF_X1 _63552_ (.D(_02294_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2325]),
    .QN(_30120_));
 DFF_X1 _63553_ (.D(_02295_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2326]),
    .QN(_30121_));
 DFF_X1 _63554_ (.D(_02296_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2327]),
    .QN(_30122_));
 DFF_X1 _63555_ (.D(_02297_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2328]),
    .QN(_30123_));
 DFF_X1 _63556_ (.D(_02298_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2329]),
    .QN(_30124_));
 DFF_X1 _63557_ (.D(_02300_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2330]),
    .QN(_30125_));
 DFF_X1 _63558_ (.D(_02301_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2331]),
    .QN(_30126_));
 DFF_X1 _63559_ (.D(_02302_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2332]),
    .QN(_30127_));
 DFF_X1 _63560_ (.D(_02303_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2333]),
    .QN(_30128_));
 DFF_X1 _63561_ (.D(_02304_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2334]),
    .QN(_30129_));
 DFF_X1 _63562_ (.D(_02305_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2335]),
    .QN(_30130_));
 DFF_X1 _63563_ (.D(_02306_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2336]),
    .QN(_30131_));
 DFF_X1 _63564_ (.D(_02307_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2337]),
    .QN(_30132_));
 DFF_X1 _63565_ (.D(_02308_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2338]),
    .QN(_30133_));
 DFF_X1 _63566_ (.D(_02309_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2339]),
    .QN(_30134_));
 DFF_X1 _63567_ (.D(_02311_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2340]),
    .QN(_30135_));
 DFF_X1 _63568_ (.D(_02312_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2341]),
    .QN(_30136_));
 DFF_X1 _63569_ (.D(_02313_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2342]),
    .QN(_30137_));
 DFF_X1 _63570_ (.D(_02314_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2343]),
    .QN(_30138_));
 DFF_X1 _63571_ (.D(_02315_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2344]),
    .QN(_30139_));
 DFF_X1 _63572_ (.D(_02316_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2345]),
    .QN(_30140_));
 DFF_X1 _63573_ (.D(_02317_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2346]),
    .QN(_30141_));
 DFF_X1 _63574_ (.D(_02318_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2347]),
    .QN(_30142_));
 DFF_X1 _63575_ (.D(_02319_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2348]),
    .QN(_30143_));
 DFF_X1 _63576_ (.D(_02320_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2349]),
    .QN(_30144_));
 DFF_X1 _63577_ (.D(_02322_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2350]),
    .QN(_30145_));
 DFF_X1 _63578_ (.D(_02323_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2351]),
    .QN(_30146_));
 DFF_X1 _63579_ (.D(_02324_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2352]),
    .QN(_30147_));
 DFF_X1 _63580_ (.D(_02325_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2353]),
    .QN(_30148_));
 DFF_X1 _63581_ (.D(_02326_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2354]),
    .QN(_30149_));
 DFF_X1 _63582_ (.D(_02327_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2355]),
    .QN(_30150_));
 DFF_X1 _63583_ (.D(_02328_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2356]),
    .QN(_30151_));
 DFF_X1 _63584_ (.D(_02329_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2357]),
    .QN(_30152_));
 DFF_X1 _63585_ (.D(_02330_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2358]),
    .QN(_30153_));
 DFF_X1 _63586_ (.D(_02331_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2359]),
    .QN(_30154_));
 DFF_X1 _63587_ (.D(_02333_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2360]),
    .QN(_30155_));
 DFF_X1 _63588_ (.D(_02334_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2361]),
    .QN(_30156_));
 DFF_X1 _63589_ (.D(_02335_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2362]),
    .QN(_30157_));
 DFF_X1 _63590_ (.D(_02336_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2363]),
    .QN(_30158_));
 DFF_X1 _63591_ (.D(_02337_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2364]),
    .QN(_30159_));
 DFF_X1 _63592_ (.D(_02338_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2365]),
    .QN(_30160_));
 DFF_X1 _63593_ (.D(_02339_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2366]),
    .QN(_30161_));
 DFF_X1 _63594_ (.D(_02340_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2367]),
    .QN(_30162_));
 DFF_X1 _63595_ (.D(_02341_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2368]),
    .QN(_30163_));
 DFF_X1 _63596_ (.D(_02342_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2369]),
    .QN(_30164_));
 DFF_X1 _63597_ (.D(_02344_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2370]),
    .QN(_30165_));
 DFF_X1 _63598_ (.D(_02345_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2371]),
    .QN(_30166_));
 DFF_X1 _63599_ (.D(_02346_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2372]),
    .QN(_30167_));
 DFF_X1 _63600_ (.D(_02347_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2373]),
    .QN(_30168_));
 DFF_X1 _63601_ (.D(_02348_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2374]),
    .QN(_30169_));
 DFF_X1 _63602_ (.D(_02349_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2375]),
    .QN(_30170_));
 DFF_X1 _63603_ (.D(_02350_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2376]),
    .QN(_30171_));
 DFF_X1 _63604_ (.D(_02351_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2377]),
    .QN(_30172_));
 DFF_X1 _63605_ (.D(_02352_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2378]),
    .QN(_30173_));
 DFF_X1 _63606_ (.D(_02353_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2379]),
    .QN(_30174_));
 DFF_X1 _63607_ (.D(_02355_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2380]),
    .QN(_30175_));
 DFF_X1 _63608_ (.D(_02356_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2381]),
    .QN(_30176_));
 DFF_X1 _63609_ (.D(_02357_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2382]),
    .QN(_30177_));
 DFF_X1 _63610_ (.D(_02358_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2383]),
    .QN(_30178_));
 DFF_X1 _63611_ (.D(_02359_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2384]),
    .QN(_30179_));
 DFF_X1 _63612_ (.D(_02360_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2385]),
    .QN(_30180_));
 DFF_X1 _63613_ (.D(_02361_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2386]),
    .QN(_30181_));
 DFF_X1 _63614_ (.D(_02362_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2387]),
    .QN(_30182_));
 DFF_X1 _63615_ (.D(_02363_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2388]),
    .QN(_30183_));
 DFF_X1 _63616_ (.D(_02364_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2389]),
    .QN(_30184_));
 DFF_X1 _63617_ (.D(_02366_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2390]),
    .QN(_30185_));
 DFF_X1 _63618_ (.D(_02367_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2391]),
    .QN(_30186_));
 DFF_X1 _63619_ (.D(_02368_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2392]),
    .QN(_30187_));
 DFF_X1 _63620_ (.D(_02369_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2393]),
    .QN(_30188_));
 DFF_X1 _63621_ (.D(_02370_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2394]),
    .QN(_30189_));
 DFF_X1 _63622_ (.D(_02371_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2395]),
    .QN(_30190_));
 DFF_X1 _63623_ (.D(_02372_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2396]),
    .QN(_30191_));
 DFF_X1 _63624_ (.D(_02373_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2397]),
    .QN(_30192_));
 DFF_X1 _63625_ (.D(_02374_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2398]),
    .QN(_30193_));
 DFF_X1 _63626_ (.D(_02375_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2399]),
    .QN(_30194_));
 DFF_X1 _63627_ (.D(_02378_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2400]),
    .QN(_30195_));
 DFF_X1 _63628_ (.D(_02379_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2401]),
    .QN(_30196_));
 DFF_X1 _63629_ (.D(_02380_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2402]),
    .QN(_30197_));
 DFF_X1 _63630_ (.D(_02381_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2403]),
    .QN(_30198_));
 DFF_X1 _63631_ (.D(_02382_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2404]),
    .QN(_30199_));
 DFF_X1 _63632_ (.D(_02383_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2405]),
    .QN(_30200_));
 DFF_X1 _63633_ (.D(_02384_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2406]),
    .QN(_30201_));
 DFF_X1 _63634_ (.D(_02385_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2407]),
    .QN(_30202_));
 DFF_X1 _63635_ (.D(_02386_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2408]),
    .QN(_30203_));
 DFF_X1 _63636_ (.D(_02387_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2409]),
    .QN(_30204_));
 DFF_X1 _63637_ (.D(_02389_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2410]),
    .QN(_30205_));
 DFF_X1 _63638_ (.D(_02390_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2411]),
    .QN(_30206_));
 DFF_X1 _63639_ (.D(_02391_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2412]),
    .QN(_30207_));
 DFF_X1 _63640_ (.D(_02392_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2413]),
    .QN(_30208_));
 DFF_X1 _63641_ (.D(_02393_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2414]),
    .QN(_30209_));
 DFF_X1 _63642_ (.D(_02394_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2415]),
    .QN(_30210_));
 DFF_X1 _63643_ (.D(_02395_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2416]),
    .QN(_30211_));
 DFF_X1 _63644_ (.D(_02396_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2417]),
    .QN(_30212_));
 DFF_X1 _63645_ (.D(_02397_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2418]),
    .QN(_30213_));
 DFF_X1 _63646_ (.D(_02398_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2419]),
    .QN(_30214_));
 DFF_X1 _63647_ (.D(_02400_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2420]),
    .QN(_30215_));
 DFF_X1 _63648_ (.D(_02401_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2421]),
    .QN(_30216_));
 DFF_X1 _63649_ (.D(_02402_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2422]),
    .QN(_30217_));
 DFF_X1 _63650_ (.D(_02403_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2423]),
    .QN(_30218_));
 DFF_X1 _63651_ (.D(_02404_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2424]),
    .QN(_30219_));
 DFF_X1 _63652_ (.D(_02405_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2425]),
    .QN(_30220_));
 DFF_X1 _63653_ (.D(_02406_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2426]),
    .QN(_30221_));
 DFF_X1 _63654_ (.D(_02407_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2427]),
    .QN(_30222_));
 DFF_X1 _63655_ (.D(_02408_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2428]),
    .QN(_30223_));
 DFF_X1 _63656_ (.D(_02409_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2429]),
    .QN(_30224_));
 DFF_X1 _63657_ (.D(_02411_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2430]),
    .QN(_30225_));
 DFF_X1 _63658_ (.D(_02412_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2431]),
    .QN(_30226_));
 DFF_X1 _63659_ (.D(_02413_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2432]),
    .QN(_30227_));
 DFF_X1 _63660_ (.D(_02414_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2433]),
    .QN(_30228_));
 DFF_X1 _63661_ (.D(_02415_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2434]),
    .QN(_30229_));
 DFF_X1 _63662_ (.D(_02416_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2435]),
    .QN(_30230_));
 DFF_X1 _63663_ (.D(_02417_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2436]),
    .QN(_30231_));
 DFF_X1 _63664_ (.D(_02418_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2437]),
    .QN(_30232_));
 DFF_X1 _63665_ (.D(_02419_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2438]),
    .QN(_30233_));
 DFF_X1 _63666_ (.D(_02420_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2439]),
    .QN(_30234_));
 DFF_X1 _63667_ (.D(_02422_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2440]),
    .QN(_30235_));
 DFF_X1 _63668_ (.D(_02423_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2441]),
    .QN(_30236_));
 DFF_X1 _63669_ (.D(_02424_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2442]),
    .QN(_30237_));
 DFF_X1 _63670_ (.D(_02425_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2443]),
    .QN(_30238_));
 DFF_X1 _63671_ (.D(_02426_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2444]),
    .QN(_30239_));
 DFF_X1 _63672_ (.D(_02427_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2445]),
    .QN(_30240_));
 DFF_X1 _63673_ (.D(_02428_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2446]),
    .QN(_30241_));
 DFF_X1 _63674_ (.D(_02429_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2447]),
    .QN(_30242_));
 DFF_X1 _63675_ (.D(_02430_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2448]),
    .QN(_30243_));
 DFF_X1 _63676_ (.D(_02431_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2449]),
    .QN(_30244_));
 DFF_X1 _63677_ (.D(_02433_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2450]),
    .QN(_30245_));
 DFF_X1 _63678_ (.D(_02434_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2451]),
    .QN(_30246_));
 DFF_X1 _63679_ (.D(_02435_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2452]),
    .QN(_30247_));
 DFF_X1 _63680_ (.D(_02436_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2453]),
    .QN(_30248_));
 DFF_X1 _63681_ (.D(_02437_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2454]),
    .QN(_30249_));
 DFF_X1 _63682_ (.D(_02438_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2455]),
    .QN(_30250_));
 DFF_X1 _63683_ (.D(_02439_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2456]),
    .QN(_30251_));
 DFF_X1 _63684_ (.D(_02440_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2457]),
    .QN(_30252_));
 DFF_X1 _63685_ (.D(_02441_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2458]),
    .QN(_30253_));
 DFF_X1 _63686_ (.D(_02442_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2459]),
    .QN(_30254_));
 DFF_X1 _63687_ (.D(_02444_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2460]),
    .QN(_30255_));
 DFF_X1 _63688_ (.D(_02445_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2461]),
    .QN(_30256_));
 DFF_X1 _63689_ (.D(_02446_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2462]),
    .QN(_30257_));
 DFF_X1 _63690_ (.D(_02447_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2463]),
    .QN(_30258_));
 DFF_X1 _63691_ (.D(_02448_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2464]),
    .QN(_30259_));
 DFF_X1 _63692_ (.D(_02449_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2465]),
    .QN(_30260_));
 DFF_X1 _63693_ (.D(_02450_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2466]),
    .QN(_30261_));
 DFF_X1 _63694_ (.D(_02451_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2467]),
    .QN(_30262_));
 DFF_X1 _63695_ (.D(_02452_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2468]),
    .QN(_30263_));
 DFF_X1 _63696_ (.D(_02453_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2469]),
    .QN(_30264_));
 DFF_X1 _63697_ (.D(_02455_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2470]),
    .QN(_30265_));
 DFF_X1 _63698_ (.D(_02456_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2471]),
    .QN(_30266_));
 DFF_X1 _63699_ (.D(_02457_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2472]),
    .QN(_30267_));
 DFF_X1 _63700_ (.D(_02458_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2473]),
    .QN(_30268_));
 DFF_X1 _63701_ (.D(_02459_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2474]),
    .QN(_30269_));
 DFF_X1 _63702_ (.D(_02460_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2475]),
    .QN(_30270_));
 DFF_X1 _63703_ (.D(_02461_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2476]),
    .QN(_30271_));
 DFF_X1 _63704_ (.D(_02462_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2477]),
    .QN(_30272_));
 DFF_X1 _63705_ (.D(_02463_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2478]),
    .QN(_30273_));
 DFF_X1 _63706_ (.D(_02464_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2479]),
    .QN(_30274_));
 DFF_X1 _63707_ (.D(_02466_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2480]),
    .QN(_30275_));
 DFF_X1 _63708_ (.D(_02467_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2481]),
    .QN(_30276_));
 DFF_X1 _63709_ (.D(_02468_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2482]),
    .QN(_30277_));
 DFF_X1 _63710_ (.D(_02469_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2483]),
    .QN(_30278_));
 DFF_X1 _63711_ (.D(_02470_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2484]),
    .QN(_30279_));
 DFF_X1 _63712_ (.D(_02471_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2485]),
    .QN(_30280_));
 DFF_X1 _63713_ (.D(_02472_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2486]),
    .QN(_30281_));
 DFF_X1 _63714_ (.D(_02473_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2487]),
    .QN(_30282_));
 DFF_X1 _63715_ (.D(_02474_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2488]),
    .QN(_30283_));
 DFF_X1 _63716_ (.D(_02475_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2489]),
    .QN(_30284_));
 DFF_X1 _63717_ (.D(_02477_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2490]),
    .QN(_30285_));
 DFF_X1 _63718_ (.D(_02478_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2491]),
    .QN(_30286_));
 DFF_X1 _63719_ (.D(_02479_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2492]),
    .QN(_30287_));
 DFF_X1 _63720_ (.D(_02480_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2493]),
    .QN(_30288_));
 DFF_X1 _63721_ (.D(_02481_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2494]),
    .QN(_30289_));
 DFF_X1 _63722_ (.D(_02482_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2495]),
    .QN(_30290_));
 DFF_X1 _63723_ (.D(_02483_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2496]),
    .QN(_30291_));
 DFF_X1 _63724_ (.D(_02484_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2497]),
    .QN(_30292_));
 DFF_X1 _63725_ (.D(_02485_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2498]),
    .QN(_30293_));
 DFF_X1 _63726_ (.D(_02486_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2499]),
    .QN(_30294_));
 DFF_X1 _63727_ (.D(_02489_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2500]),
    .QN(_30295_));
 DFF_X1 _63728_ (.D(_02490_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2501]),
    .QN(_30296_));
 DFF_X1 _63729_ (.D(_02491_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2502]),
    .QN(_30297_));
 DFF_X1 _63730_ (.D(_02492_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2503]),
    .QN(_30298_));
 DFF_X1 _63731_ (.D(_02493_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2504]),
    .QN(_30299_));
 DFF_X1 _63732_ (.D(_02494_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2505]),
    .QN(_30300_));
 DFF_X1 _63733_ (.D(_02495_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2506]),
    .QN(_30301_));
 DFF_X1 _63734_ (.D(_02496_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2507]),
    .QN(_30302_));
 DFF_X1 _63735_ (.D(_02497_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2508]),
    .QN(_30303_));
 DFF_X1 _63736_ (.D(_02498_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2509]),
    .QN(_30304_));
 DFF_X1 _63737_ (.D(_02500_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2510]),
    .QN(_30305_));
 DFF_X1 _63738_ (.D(_02501_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2511]),
    .QN(_30306_));
 DFF_X1 _63739_ (.D(_02502_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2512]),
    .QN(_30307_));
 DFF_X1 _63740_ (.D(_02503_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2513]),
    .QN(_30308_));
 DFF_X1 _63741_ (.D(_02504_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2514]),
    .QN(_30309_));
 DFF_X1 _63742_ (.D(_02505_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2515]),
    .QN(_30310_));
 DFF_X1 _63743_ (.D(_02506_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2516]),
    .QN(_30311_));
 DFF_X1 _63744_ (.D(_02507_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2517]),
    .QN(_30312_));
 DFF_X1 _63745_ (.D(_02508_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2518]),
    .QN(_30313_));
 DFF_X1 _63746_ (.D(_02509_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2519]),
    .QN(_30314_));
 DFF_X1 _63747_ (.D(_02511_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2520]),
    .QN(_30315_));
 DFF_X1 _63748_ (.D(_02512_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2521]),
    .QN(_30316_));
 DFF_X1 _63749_ (.D(_02513_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2522]),
    .QN(_30317_));
 DFF_X1 _63750_ (.D(_02514_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2523]),
    .QN(_30318_));
 DFF_X1 _63751_ (.D(_02515_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2524]),
    .QN(_30319_));
 DFF_X1 _63752_ (.D(_02516_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2525]),
    .QN(_30320_));
 DFF_X1 _63753_ (.D(_02517_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2526]),
    .QN(_30321_));
 DFF_X1 _63754_ (.D(_02518_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2527]),
    .QN(_30322_));
 DFF_X1 _63755_ (.D(_02519_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2528]),
    .QN(_30323_));
 DFF_X1 _63756_ (.D(_02520_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2529]),
    .QN(_30324_));
 DFF_X1 _63757_ (.D(_02522_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2530]),
    .QN(_30325_));
 DFF_X1 _63758_ (.D(_02523_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2531]),
    .QN(_30326_));
 DFF_X1 _63759_ (.D(_02524_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2532]),
    .QN(_30327_));
 DFF_X1 _63760_ (.D(_02525_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2533]),
    .QN(_30328_));
 DFF_X1 _63761_ (.D(_02526_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2534]),
    .QN(_30329_));
 DFF_X1 _63762_ (.D(_02527_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2535]),
    .QN(_30330_));
 DFF_X1 _63763_ (.D(_02528_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2536]),
    .QN(_30331_));
 DFF_X1 _63764_ (.D(_02529_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2537]),
    .QN(_30332_));
 DFF_X1 _63765_ (.D(_02530_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2538]),
    .QN(_30333_));
 DFF_X1 _63766_ (.D(_02531_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2539]),
    .QN(_30334_));
 DFF_X1 _63767_ (.D(_02533_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2540]),
    .QN(_30335_));
 DFF_X1 _63768_ (.D(_02534_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2541]),
    .QN(_30336_));
 DFF_X1 _63769_ (.D(_02535_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2542]),
    .QN(_30337_));
 DFF_X1 _63770_ (.D(_02536_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2543]),
    .QN(_30338_));
 DFF_X1 _63771_ (.D(_02537_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2544]),
    .QN(_30339_));
 DFF_X1 _63772_ (.D(_02538_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2545]),
    .QN(_30340_));
 DFF_X1 _63773_ (.D(_02539_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2546]),
    .QN(_30341_));
 DFF_X1 _63774_ (.D(_02540_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2547]),
    .QN(_30342_));
 DFF_X1 _63775_ (.D(_02541_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2548]),
    .QN(_30343_));
 DFF_X1 _63776_ (.D(_02542_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2549]),
    .QN(_30344_));
 DFF_X1 _63777_ (.D(_02544_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2550]),
    .QN(_30345_));
 DFF_X1 _63778_ (.D(_02545_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2551]),
    .QN(_30346_));
 DFF_X1 _63779_ (.D(_02546_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2552]),
    .QN(_30347_));
 DFF_X1 _63780_ (.D(_02547_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2553]),
    .QN(_30348_));
 DFF_X1 _63781_ (.D(_02548_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2554]),
    .QN(_30349_));
 DFF_X1 _63782_ (.D(_02549_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2555]),
    .QN(_30350_));
 DFF_X1 _63783_ (.D(_02550_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2556]),
    .QN(_30351_));
 DFF_X1 _63784_ (.D(_02551_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2557]),
    .QN(_30352_));
 DFF_X1 _63785_ (.D(_02552_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2558]),
    .QN(_30353_));
 DFF_X1 _63786_ (.D(_02553_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2559]),
    .QN(_30354_));
 DFF_X1 _63787_ (.D(_02555_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2560]),
    .QN(_30355_));
 DFF_X1 _63788_ (.D(_02556_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2561]),
    .QN(_30356_));
 DFF_X1 _63789_ (.D(_02557_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2562]),
    .QN(_30357_));
 DFF_X1 _63790_ (.D(_02558_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2563]),
    .QN(_30358_));
 DFF_X1 _63791_ (.D(_02559_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2564]),
    .QN(_30359_));
 DFF_X1 _63792_ (.D(_02560_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2565]),
    .QN(_30360_));
 DFF_X1 _63793_ (.D(_02561_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2566]),
    .QN(_30361_));
 DFF_X1 _63794_ (.D(_02562_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2567]),
    .QN(_30362_));
 DFF_X1 _63795_ (.D(_02563_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2568]),
    .QN(_30363_));
 DFF_X1 _63796_ (.D(_02564_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2569]),
    .QN(_30364_));
 DFF_X1 _63797_ (.D(_02566_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2570]),
    .QN(_30365_));
 DFF_X1 _63798_ (.D(_02567_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2571]),
    .QN(_30366_));
 DFF_X1 _63799_ (.D(_02568_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2572]),
    .QN(_30367_));
 DFF_X1 _63800_ (.D(_02569_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2573]),
    .QN(_30368_));
 DFF_X1 _63801_ (.D(_02570_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2574]),
    .QN(_30369_));
 DFF_X1 _63802_ (.D(_02571_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2575]),
    .QN(_30370_));
 DFF_X1 _63803_ (.D(_02572_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2576]),
    .QN(_30371_));
 DFF_X1 _63804_ (.D(_02573_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2577]),
    .QN(_30372_));
 DFF_X1 _63805_ (.D(_02574_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2578]),
    .QN(_30373_));
 DFF_X1 _63806_ (.D(_02575_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2579]),
    .QN(_30374_));
 DFF_X1 _63807_ (.D(_02577_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2580]),
    .QN(_30375_));
 DFF_X1 _63808_ (.D(_02578_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2581]),
    .QN(_30376_));
 DFF_X1 _63809_ (.D(_02579_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2582]),
    .QN(_30377_));
 DFF_X1 _63810_ (.D(_02580_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2583]),
    .QN(_30378_));
 DFF_X1 _63811_ (.D(_02581_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2584]),
    .QN(_30379_));
 DFF_X1 _63812_ (.D(_02582_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2585]),
    .QN(_30380_));
 DFF_X1 _63813_ (.D(_02583_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2586]),
    .QN(_30381_));
 DFF_X1 _63814_ (.D(_02584_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2587]),
    .QN(_30382_));
 DFF_X1 _63815_ (.D(_02585_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2588]),
    .QN(_30383_));
 DFF_X1 _63816_ (.D(_02586_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2589]),
    .QN(_30384_));
 DFF_X1 _63817_ (.D(_02588_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2590]),
    .QN(_30385_));
 DFF_X1 _63818_ (.D(_02589_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2591]),
    .QN(_30386_));
 DFF_X1 _63819_ (.D(_02590_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2592]),
    .QN(_30387_));
 DFF_X1 _63820_ (.D(_02591_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2593]),
    .QN(_30388_));
 DFF_X1 _63821_ (.D(_02592_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2594]),
    .QN(_30389_));
 DFF_X1 _63822_ (.D(_02593_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2595]),
    .QN(_30390_));
 DFF_X1 _63823_ (.D(_02594_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2596]),
    .QN(_30391_));
 DFF_X1 _63824_ (.D(_02595_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2597]),
    .QN(_30392_));
 DFF_X1 _63825_ (.D(_02596_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2598]),
    .QN(_30393_));
 DFF_X1 _63826_ (.D(_02597_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2599]),
    .QN(_30394_));
 DFF_X1 _63827_ (.D(_02600_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2600]),
    .QN(_30395_));
 DFF_X1 _63828_ (.D(_02601_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2601]),
    .QN(_30396_));
 DFF_X1 _63829_ (.D(_02602_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2602]),
    .QN(_30397_));
 DFF_X1 _63830_ (.D(_02603_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2603]),
    .QN(_30398_));
 DFF_X1 _63831_ (.D(_02604_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2604]),
    .QN(_30399_));
 DFF_X1 _63832_ (.D(_02605_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2605]),
    .QN(_30400_));
 DFF_X1 _63833_ (.D(_02606_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2606]),
    .QN(_30401_));
 DFF_X1 _63834_ (.D(_02607_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2607]),
    .QN(_30402_));
 DFF_X1 _63835_ (.D(_02608_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2608]),
    .QN(_30403_));
 DFF_X1 _63836_ (.D(_02609_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2609]),
    .QN(_30404_));
 DFF_X1 _63837_ (.D(_02611_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2610]),
    .QN(_30405_));
 DFF_X1 _63838_ (.D(_02612_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2611]),
    .QN(_30406_));
 DFF_X1 _63839_ (.D(_02613_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2612]),
    .QN(_30407_));
 DFF_X1 _63840_ (.D(_02614_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2613]),
    .QN(_30408_));
 DFF_X1 _63841_ (.D(_02615_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2614]),
    .QN(_30409_));
 DFF_X1 _63842_ (.D(_02616_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2615]),
    .QN(_30410_));
 DFF_X1 _63843_ (.D(_02617_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2616]),
    .QN(_30411_));
 DFF_X1 _63844_ (.D(_02618_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2617]),
    .QN(_30412_));
 DFF_X1 _63845_ (.D(_02619_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2618]),
    .QN(_30413_));
 DFF_X1 _63846_ (.D(_02620_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2619]),
    .QN(_30414_));
 DFF_X1 _63847_ (.D(_02622_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2620]),
    .QN(_30415_));
 DFF_X1 _63848_ (.D(_02623_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2621]),
    .QN(_30416_));
 DFF_X1 _63849_ (.D(_02624_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2622]),
    .QN(_30417_));
 DFF_X1 _63850_ (.D(_02625_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2623]),
    .QN(_30418_));
 DFF_X1 _63851_ (.D(_02626_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2624]),
    .QN(_30419_));
 DFF_X1 _63852_ (.D(_02627_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2625]),
    .QN(_30420_));
 DFF_X1 _63853_ (.D(_02628_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2626]),
    .QN(_30421_));
 DFF_X1 _63854_ (.D(_02629_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2627]),
    .QN(_30422_));
 DFF_X1 _63855_ (.D(_02630_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2628]),
    .QN(_30423_));
 DFF_X1 _63856_ (.D(_02631_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2629]),
    .QN(_30424_));
 DFF_X1 _63857_ (.D(_02633_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2630]),
    .QN(_30425_));
 DFF_X1 _63858_ (.D(_02634_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2631]),
    .QN(_30426_));
 DFF_X1 _63859_ (.D(_02635_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2632]),
    .QN(_30427_));
 DFF_X1 _63860_ (.D(_02636_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2633]),
    .QN(_30428_));
 DFF_X1 _63861_ (.D(_02637_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2634]),
    .QN(_30429_));
 DFF_X1 _63862_ (.D(_02638_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2635]),
    .QN(_30430_));
 DFF_X1 _63863_ (.D(_02639_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2636]),
    .QN(_30431_));
 DFF_X1 _63864_ (.D(_02640_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2637]),
    .QN(_30432_));
 DFF_X1 _63865_ (.D(_02641_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2638]),
    .QN(_30433_));
 DFF_X1 _63866_ (.D(_02642_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2639]),
    .QN(_30434_));
 DFF_X1 _63867_ (.D(_02644_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2640]),
    .QN(_30435_));
 DFF_X1 _63868_ (.D(_02645_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2641]),
    .QN(_30436_));
 DFF_X1 _63869_ (.D(_02646_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2642]),
    .QN(_30437_));
 DFF_X1 _63870_ (.D(_02647_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2643]),
    .QN(_30438_));
 DFF_X1 _63871_ (.D(_02648_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2644]),
    .QN(_30439_));
 DFF_X1 _63872_ (.D(_02649_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2645]),
    .QN(_30440_));
 DFF_X1 _63873_ (.D(_02650_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2646]),
    .QN(_30441_));
 DFF_X1 _63874_ (.D(_02651_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2647]),
    .QN(_30442_));
 DFF_X1 _63875_ (.D(_02652_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2648]),
    .QN(_30443_));
 DFF_X1 _63876_ (.D(_02653_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2649]),
    .QN(_30444_));
 DFF_X1 _63877_ (.D(_02655_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2650]),
    .QN(_30445_));
 DFF_X1 _63878_ (.D(_02656_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2651]),
    .QN(_30446_));
 DFF_X1 _63879_ (.D(_02657_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2652]),
    .QN(_30447_));
 DFF_X1 _63880_ (.D(_02658_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2653]),
    .QN(_30448_));
 DFF_X1 _63881_ (.D(_02659_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2654]),
    .QN(_30449_));
 DFF_X1 _63882_ (.D(_02660_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2655]),
    .QN(_30450_));
 DFF_X1 _63883_ (.D(_02661_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2656]),
    .QN(_30451_));
 DFF_X1 _63884_ (.D(_02662_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2657]),
    .QN(_30452_));
 DFF_X1 _63885_ (.D(_02663_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2658]),
    .QN(_30453_));
 DFF_X1 _63886_ (.D(_02664_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2659]),
    .QN(_30454_));
 DFF_X1 _63887_ (.D(_02666_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2660]),
    .QN(_30455_));
 DFF_X1 _63888_ (.D(_02667_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2661]),
    .QN(_30456_));
 DFF_X1 _63889_ (.D(_02668_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2662]),
    .QN(_30457_));
 DFF_X1 _63890_ (.D(_02669_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2663]),
    .QN(_30458_));
 DFF_X1 _63891_ (.D(_02670_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2664]),
    .QN(_30459_));
 DFF_X1 _63892_ (.D(_02671_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2665]),
    .QN(_30460_));
 DFF_X1 _63893_ (.D(_02672_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2666]),
    .QN(_30461_));
 DFF_X1 _63894_ (.D(_02673_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2667]),
    .QN(_30462_));
 DFF_X1 _63895_ (.D(_02674_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2668]),
    .QN(_30463_));
 DFF_X1 _63896_ (.D(_02675_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2669]),
    .QN(_30464_));
 DFF_X1 _63897_ (.D(_02677_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2670]),
    .QN(_30465_));
 DFF_X1 _63898_ (.D(_02678_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2671]),
    .QN(_30466_));
 DFF_X1 _63899_ (.D(_02679_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2672]),
    .QN(_30467_));
 DFF_X1 _63900_ (.D(_02680_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2673]),
    .QN(_30468_));
 DFF_X1 _63901_ (.D(_02681_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2674]),
    .QN(_30469_));
 DFF_X1 _63902_ (.D(_02682_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2675]),
    .QN(_30470_));
 DFF_X1 _63903_ (.D(_02683_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2676]),
    .QN(_30471_));
 DFF_X1 _63904_ (.D(_02684_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2677]),
    .QN(_30472_));
 DFF_X1 _63905_ (.D(_02685_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2678]),
    .QN(_30473_));
 DFF_X1 _63906_ (.D(_02686_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2679]),
    .QN(_30474_));
 DFF_X1 _63907_ (.D(_02688_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2680]),
    .QN(_30475_));
 DFF_X1 _63908_ (.D(_02689_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2681]),
    .QN(_30476_));
 DFF_X1 _63909_ (.D(_02690_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2682]),
    .QN(_30477_));
 DFF_X1 _63910_ (.D(_02691_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2683]),
    .QN(_30478_));
 DFF_X1 _63911_ (.D(_02692_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2684]),
    .QN(_30479_));
 DFF_X1 _63912_ (.D(_02693_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2685]),
    .QN(_30480_));
 DFF_X1 _63913_ (.D(_02694_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2686]),
    .QN(_30481_));
 DFF_X1 _63914_ (.D(_02695_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2687]),
    .QN(_30482_));
 DFF_X1 _63915_ (.D(_02696_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2688]),
    .QN(_30483_));
 DFF_X1 _63916_ (.D(_02697_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2689]),
    .QN(_30484_));
 DFF_X1 _63917_ (.D(_02699_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2690]),
    .QN(_30485_));
 DFF_X1 _63918_ (.D(_02700_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2691]),
    .QN(_30486_));
 DFF_X1 _63919_ (.D(_02701_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2692]),
    .QN(_30487_));
 DFF_X1 _63920_ (.D(_02702_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2693]),
    .QN(_30488_));
 DFF_X1 _63921_ (.D(_02703_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2694]),
    .QN(_30489_));
 DFF_X1 _63922_ (.D(_02704_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2695]),
    .QN(_30490_));
 DFF_X1 _63923_ (.D(_02705_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2696]),
    .QN(_30491_));
 DFF_X1 _63924_ (.D(_02706_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2697]),
    .QN(_30492_));
 DFF_X1 _63925_ (.D(_02707_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2698]),
    .QN(_30493_));
 DFF_X1 _63926_ (.D(_02708_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2699]),
    .QN(_30494_));
 DFF_X1 _63927_ (.D(_02711_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2700]),
    .QN(_30495_));
 DFF_X1 _63928_ (.D(_02712_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2701]),
    .QN(_30496_));
 DFF_X1 _63929_ (.D(_02713_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2702]),
    .QN(_30497_));
 DFF_X1 _63930_ (.D(_02714_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2703]),
    .QN(_30498_));
 DFF_X1 _63931_ (.D(_02715_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2704]),
    .QN(_30499_));
 DFF_X1 _63932_ (.D(_02716_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2705]),
    .QN(_30500_));
 DFF_X1 _63933_ (.D(_02717_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2706]),
    .QN(_30501_));
 DFF_X1 _63934_ (.D(_02718_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2707]),
    .QN(_30502_));
 DFF_X1 _63935_ (.D(_02719_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2708]),
    .QN(_30503_));
 DFF_X1 _63936_ (.D(_02720_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2709]),
    .QN(_30504_));
 DFF_X1 _63937_ (.D(_02722_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2710]),
    .QN(_30505_));
 DFF_X1 _63938_ (.D(_02723_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2711]),
    .QN(_30506_));
 DFF_X1 _63939_ (.D(_02724_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2712]),
    .QN(_30507_));
 DFF_X1 _63940_ (.D(_02725_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2713]),
    .QN(_30508_));
 DFF_X1 _63941_ (.D(_02726_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2714]),
    .QN(_30509_));
 DFF_X1 _63942_ (.D(_02727_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2715]),
    .QN(_30510_));
 DFF_X1 _63943_ (.D(_02728_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2716]),
    .QN(_30511_));
 DFF_X1 _63944_ (.D(_02729_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2717]),
    .QN(_30512_));
 DFF_X1 _63945_ (.D(_02730_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2718]),
    .QN(_30513_));
 DFF_X1 _63946_ (.D(_02731_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2719]),
    .QN(_30514_));
 DFF_X1 _63947_ (.D(_02733_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2720]),
    .QN(_30515_));
 DFF_X1 _63948_ (.D(_02734_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2721]),
    .QN(_30516_));
 DFF_X1 _63949_ (.D(_02735_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2722]),
    .QN(_30517_));
 DFF_X1 _63950_ (.D(_02736_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2723]),
    .QN(_30518_));
 DFF_X1 _63951_ (.D(_02737_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2724]),
    .QN(_30519_));
 DFF_X1 _63952_ (.D(_02738_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2725]),
    .QN(_30520_));
 DFF_X1 _63953_ (.D(_02739_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2726]),
    .QN(_30521_));
 DFF_X1 _63954_ (.D(_02740_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2727]),
    .QN(_30522_));
 DFF_X1 _63955_ (.D(_02741_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2728]),
    .QN(_30523_));
 DFF_X1 _63956_ (.D(_02742_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2729]),
    .QN(_30524_));
 DFF_X1 _63957_ (.D(_02744_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2730]),
    .QN(_30525_));
 DFF_X1 _63958_ (.D(_02745_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2731]),
    .QN(_30526_));
 DFF_X1 _63959_ (.D(_02746_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2732]),
    .QN(_30527_));
 DFF_X1 _63960_ (.D(_02747_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2733]),
    .QN(_30528_));
 DFF_X1 _63961_ (.D(_02748_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2734]),
    .QN(_30529_));
 DFF_X1 _63962_ (.D(_02749_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2735]),
    .QN(_30530_));
 DFF_X1 _63963_ (.D(_02750_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2736]),
    .QN(_30531_));
 DFF_X1 _63964_ (.D(_02751_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2737]),
    .QN(_30532_));
 DFF_X1 _63965_ (.D(_02752_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2738]),
    .QN(_30533_));
 DFF_X1 _63966_ (.D(_02753_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2739]),
    .QN(_30534_));
 DFF_X1 _63967_ (.D(_02755_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2740]),
    .QN(_30535_));
 DFF_X1 _63968_ (.D(_02756_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2741]),
    .QN(_30536_));
 DFF_X1 _63969_ (.D(_02757_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2742]),
    .QN(_30537_));
 DFF_X1 _63970_ (.D(_02758_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2743]),
    .QN(_30538_));
 DFF_X1 _63971_ (.D(_02759_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2744]),
    .QN(_30539_));
 DFF_X1 _63972_ (.D(_02760_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2745]),
    .QN(_30540_));
 DFF_X1 _63973_ (.D(_02761_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2746]),
    .QN(_30541_));
 DFF_X1 _63974_ (.D(_02762_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2747]),
    .QN(_30542_));
 DFF_X1 _63975_ (.D(_02763_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2748]),
    .QN(_30543_));
 DFF_X1 _63976_ (.D(_02764_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2749]),
    .QN(_30544_));
 DFF_X1 _63977_ (.D(_02766_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2750]),
    .QN(_30545_));
 DFF_X1 _63978_ (.D(_02767_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2751]),
    .QN(_30546_));
 DFF_X1 _63979_ (.D(_02768_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2752]),
    .QN(_30547_));
 DFF_X1 _63980_ (.D(_02769_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2753]),
    .QN(_30548_));
 DFF_X1 _63981_ (.D(_02770_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2754]),
    .QN(_30549_));
 DFF_X1 _63982_ (.D(_02771_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2755]),
    .QN(_30550_));
 DFF_X1 _63983_ (.D(_02772_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2756]),
    .QN(_30551_));
 DFF_X1 _63984_ (.D(_02773_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2757]),
    .QN(_30552_));
 DFF_X1 _63985_ (.D(_02774_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2758]),
    .QN(_30553_));
 DFF_X1 _63986_ (.D(_02775_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2759]),
    .QN(_30554_));
 DFF_X1 _63987_ (.D(_02777_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2760]),
    .QN(_30555_));
 DFF_X1 _63988_ (.D(_02778_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2761]),
    .QN(_30556_));
 DFF_X1 _63989_ (.D(_02779_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2762]),
    .QN(_30557_));
 DFF_X1 _63990_ (.D(_02780_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2763]),
    .QN(_30558_));
 DFF_X1 _63991_ (.D(_02781_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2764]),
    .QN(_30559_));
 DFF_X1 _63992_ (.D(_02782_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2765]),
    .QN(_30560_));
 DFF_X1 _63993_ (.D(_02783_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2766]),
    .QN(_30561_));
 DFF_X1 _63994_ (.D(_02784_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2767]),
    .QN(_30562_));
 DFF_X1 _63995_ (.D(_02785_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2768]),
    .QN(_30563_));
 DFF_X1 _63996_ (.D(_02786_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2769]),
    .QN(_30564_));
 DFF_X1 _63997_ (.D(_02788_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2770]),
    .QN(_30565_));
 DFF_X1 _63998_ (.D(_02789_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2771]),
    .QN(_30566_));
 DFF_X1 _63999_ (.D(_02790_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2772]),
    .QN(_30567_));
 DFF_X1 _64000_ (.D(_02791_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2773]),
    .QN(_30568_));
 DFF_X1 _64001_ (.D(_02792_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2774]),
    .QN(_30569_));
 DFF_X1 _64002_ (.D(_02793_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2775]),
    .QN(_30570_));
 DFF_X1 _64003_ (.D(_02794_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2776]),
    .QN(_30571_));
 DFF_X1 _64004_ (.D(_02795_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2777]),
    .QN(_30572_));
 DFF_X1 _64005_ (.D(_02796_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2778]),
    .QN(_30573_));
 DFF_X1 _64006_ (.D(_02797_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2779]),
    .QN(_30574_));
 DFF_X1 _64007_ (.D(_02799_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2780]),
    .QN(_30575_));
 DFF_X1 _64008_ (.D(_02800_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2781]),
    .QN(_30576_));
 DFF_X1 _64009_ (.D(_02801_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2782]),
    .QN(_30577_));
 DFF_X1 _64010_ (.D(_02802_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2783]),
    .QN(_30578_));
 DFF_X1 _64011_ (.D(_02803_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2784]),
    .QN(_30579_));
 DFF_X1 _64012_ (.D(_02804_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2785]),
    .QN(_30580_));
 DFF_X1 _64013_ (.D(_02805_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2786]),
    .QN(_30581_));
 DFF_X1 _64014_ (.D(_02806_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2787]),
    .QN(_30582_));
 DFF_X1 _64015_ (.D(_02807_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2788]),
    .QN(_30583_));
 DFF_X1 _64016_ (.D(_02808_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2789]),
    .QN(_30584_));
 DFF_X1 _64017_ (.D(_02810_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2790]),
    .QN(_30585_));
 DFF_X1 _64018_ (.D(_02811_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2791]),
    .QN(_30586_));
 DFF_X1 _64019_ (.D(_02812_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2792]),
    .QN(_30587_));
 DFF_X1 _64020_ (.D(_02813_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2793]),
    .QN(_30588_));
 DFF_X1 _64021_ (.D(_02814_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2794]),
    .QN(_30589_));
 DFF_X1 _64022_ (.D(_02815_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2795]),
    .QN(_30590_));
 DFF_X1 _64023_ (.D(_02816_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2796]),
    .QN(_30591_));
 DFF_X1 _64024_ (.D(_02817_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2797]),
    .QN(_30592_));
 DFF_X1 _64025_ (.D(_02818_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2798]),
    .QN(_30593_));
 DFF_X1 _64026_ (.D(_02819_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2799]),
    .QN(_30594_));
 DFF_X1 _64027_ (.D(_02822_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2800]),
    .QN(_30595_));
 DFF_X1 _64028_ (.D(_02823_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2801]),
    .QN(_30596_));
 DFF_X1 _64029_ (.D(_02824_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2802]),
    .QN(_30597_));
 DFF_X1 _64030_ (.D(_02825_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2803]),
    .QN(_30598_));
 DFF_X1 _64031_ (.D(_02826_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2804]),
    .QN(_30599_));
 DFF_X1 _64032_ (.D(_02827_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2805]),
    .QN(_30600_));
 DFF_X1 _64033_ (.D(_02828_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2806]),
    .QN(_30601_));
 DFF_X1 _64034_ (.D(_02829_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2807]),
    .QN(_30602_));
 DFF_X1 _64035_ (.D(_02830_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2808]),
    .QN(_30603_));
 DFF_X1 _64036_ (.D(_02831_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2809]),
    .QN(_30604_));
 DFF_X1 _64037_ (.D(_02833_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2810]),
    .QN(_30605_));
 DFF_X1 _64038_ (.D(_02834_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2811]),
    .QN(_30606_));
 DFF_X1 _64039_ (.D(_02835_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2812]),
    .QN(_30607_));
 DFF_X1 _64040_ (.D(_02836_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2813]),
    .QN(_30608_));
 DFF_X1 _64041_ (.D(_02837_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2814]),
    .QN(_30609_));
 DFF_X1 _64042_ (.D(_02838_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2815]),
    .QN(_30610_));
 DFF_X1 _64043_ (.D(_02839_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2816]),
    .QN(_30611_));
 DFF_X1 _64044_ (.D(_02840_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2817]),
    .QN(_30612_));
 DFF_X1 _64045_ (.D(_02841_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2818]),
    .QN(_30613_));
 DFF_X1 _64046_ (.D(_02842_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2819]),
    .QN(_30614_));
 DFF_X1 _64047_ (.D(_02844_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2820]),
    .QN(_30615_));
 DFF_X1 _64048_ (.D(_02845_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2821]),
    .QN(_30616_));
 DFF_X1 _64049_ (.D(_02846_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2822]),
    .QN(_30617_));
 DFF_X1 _64050_ (.D(_02847_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2823]),
    .QN(_30618_));
 DFF_X1 _64051_ (.D(_02848_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2824]),
    .QN(_30619_));
 DFF_X1 _64052_ (.D(_02849_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2825]),
    .QN(_30620_));
 DFF_X1 _64053_ (.D(_02850_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2826]),
    .QN(_30621_));
 DFF_X1 _64054_ (.D(_02851_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2827]),
    .QN(_30622_));
 DFF_X1 _64055_ (.D(_02852_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2828]),
    .QN(_30623_));
 DFF_X1 _64056_ (.D(_02853_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2829]),
    .QN(_30624_));
 DFF_X1 _64057_ (.D(_02855_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2830]),
    .QN(_30625_));
 DFF_X1 _64058_ (.D(_02856_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2831]),
    .QN(_30626_));
 DFF_X1 _64059_ (.D(_02857_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2832]),
    .QN(_30627_));
 DFF_X1 _64060_ (.D(_02858_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2833]),
    .QN(_30628_));
 DFF_X1 _64061_ (.D(_02859_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2834]),
    .QN(_30629_));
 DFF_X1 _64062_ (.D(_02860_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2835]),
    .QN(_30630_));
 DFF_X1 _64063_ (.D(_02861_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2836]),
    .QN(_30631_));
 DFF_X1 _64064_ (.D(_02862_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2837]),
    .QN(_30632_));
 DFF_X1 _64065_ (.D(_02863_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2838]),
    .QN(_30633_));
 DFF_X1 _64066_ (.D(_02864_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2839]),
    .QN(_30634_));
 DFF_X1 _64067_ (.D(_02866_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2840]),
    .QN(_30635_));
 DFF_X1 _64068_ (.D(_02867_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2841]),
    .QN(_30636_));
 DFF_X1 _64069_ (.D(_02868_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2842]),
    .QN(_30637_));
 DFF_X1 _64070_ (.D(_02869_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2843]),
    .QN(_30638_));
 DFF_X1 _64071_ (.D(_02870_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2844]),
    .QN(_30639_));
 DFF_X1 _64072_ (.D(_02871_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2845]),
    .QN(_30640_));
 DFF_X1 _64073_ (.D(_02872_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2846]),
    .QN(_30641_));
 DFF_X1 _64074_ (.D(_02873_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2847]),
    .QN(_30642_));
 DFF_X1 _64075_ (.D(_02874_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2848]),
    .QN(_30643_));
 DFF_X1 _64076_ (.D(_02875_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2849]),
    .QN(_30644_));
 DFF_X1 _64077_ (.D(_02877_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2850]),
    .QN(_30645_));
 DFF_X1 _64078_ (.D(_02878_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2851]),
    .QN(_30646_));
 DFF_X1 _64079_ (.D(_02879_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2852]),
    .QN(_30647_));
 DFF_X1 _64080_ (.D(_02880_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2853]),
    .QN(_30648_));
 DFF_X1 _64081_ (.D(_02881_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2854]),
    .QN(_30649_));
 DFF_X1 _64082_ (.D(_02882_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2855]),
    .QN(_30650_));
 DFF_X1 _64083_ (.D(_02883_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2856]),
    .QN(_30651_));
 DFF_X1 _64084_ (.D(_02884_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2857]),
    .QN(_30652_));
 DFF_X1 _64085_ (.D(_02885_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2858]),
    .QN(_30653_));
 DFF_X1 _64086_ (.D(_02886_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2859]),
    .QN(_30654_));
 DFF_X1 _64087_ (.D(_02888_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2860]),
    .QN(_30655_));
 DFF_X1 _64088_ (.D(_02889_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2861]),
    .QN(_30656_));
 DFF_X1 _64089_ (.D(_02890_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2862]),
    .QN(_30657_));
 DFF_X1 _64090_ (.D(_02891_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2863]),
    .QN(_30658_));
 DFF_X1 _64091_ (.D(_02892_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2864]),
    .QN(_30659_));
 DFF_X1 _64092_ (.D(_02893_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2865]),
    .QN(_30660_));
 DFF_X1 _64093_ (.D(_02894_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2866]),
    .QN(_30661_));
 DFF_X1 _64094_ (.D(_02895_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2867]),
    .QN(_30662_));
 DFF_X1 _64095_ (.D(_02896_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2868]),
    .QN(_30663_));
 DFF_X1 _64096_ (.D(_02897_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2869]),
    .QN(_30664_));
 DFF_X1 _64097_ (.D(_02899_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2870]),
    .QN(_30665_));
 DFF_X1 _64098_ (.D(_02900_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2871]),
    .QN(_30666_));
 DFF_X1 _64099_ (.D(_02901_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2872]),
    .QN(_30667_));
 DFF_X1 _64100_ (.D(_02902_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2873]),
    .QN(_30668_));
 DFF_X1 _64101_ (.D(_02903_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2874]),
    .QN(_30669_));
 DFF_X1 _64102_ (.D(_02904_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2875]),
    .QN(_30670_));
 DFF_X1 _64103_ (.D(_02905_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2876]),
    .QN(_30671_));
 DFF_X1 _64104_ (.D(_02906_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2877]),
    .QN(_30672_));
 DFF_X1 _64105_ (.D(_02907_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2878]),
    .QN(_30673_));
 DFF_X1 _64106_ (.D(_02908_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2879]),
    .QN(_30674_));
 DFF_X1 _64107_ (.D(_02910_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2880]),
    .QN(_30675_));
 DFF_X1 _64108_ (.D(_02911_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2881]),
    .QN(_30676_));
 DFF_X1 _64109_ (.D(_02912_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2882]),
    .QN(_30677_));
 DFF_X1 _64110_ (.D(_02913_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2883]),
    .QN(_30678_));
 DFF_X1 _64111_ (.D(_02914_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2884]),
    .QN(_30679_));
 DFF_X1 _64112_ (.D(_02915_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2885]),
    .QN(_30680_));
 DFF_X1 _64113_ (.D(_02916_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2886]),
    .QN(_30681_));
 DFF_X1 _64114_ (.D(_02917_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2887]),
    .QN(_30682_));
 DFF_X1 _64115_ (.D(_02918_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2888]),
    .QN(_30683_));
 DFF_X1 _64116_ (.D(_02919_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2889]),
    .QN(_30684_));
 DFF_X1 _64117_ (.D(_02921_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2890]),
    .QN(_30685_));
 DFF_X1 _64118_ (.D(_02922_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2891]),
    .QN(_30686_));
 DFF_X1 _64119_ (.D(_02923_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2892]),
    .QN(_30687_));
 DFF_X1 _64120_ (.D(_02924_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2893]),
    .QN(_30688_));
 DFF_X1 _64121_ (.D(_02925_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2894]),
    .QN(_30689_));
 DFF_X1 _64122_ (.D(_02926_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2895]),
    .QN(_30690_));
 DFF_X1 _64123_ (.D(_02927_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2896]),
    .QN(_30691_));
 DFF_X1 _64124_ (.D(_02928_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2897]),
    .QN(_30692_));
 DFF_X1 _64125_ (.D(_02929_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2898]),
    .QN(_30693_));
 DFF_X1 _64126_ (.D(_02930_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2899]),
    .QN(_30694_));
 DFF_X1 _64127_ (.D(_02933_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2900]),
    .QN(_30695_));
 DFF_X1 _64128_ (.D(_02934_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2901]),
    .QN(_30696_));
 DFF_X1 _64129_ (.D(_02935_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2902]),
    .QN(_30697_));
 DFF_X1 _64130_ (.D(_02936_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2903]),
    .QN(_30698_));
 DFF_X1 _64131_ (.D(_02937_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2904]),
    .QN(_30699_));
 DFF_X1 _64132_ (.D(_02938_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2905]),
    .QN(_30700_));
 DFF_X1 _64133_ (.D(_02939_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2906]),
    .QN(_30701_));
 DFF_X1 _64134_ (.D(_02940_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2907]),
    .QN(_30702_));
 DFF_X1 _64135_ (.D(_02941_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2908]),
    .QN(_30703_));
 DFF_X1 _64136_ (.D(_02942_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2909]),
    .QN(_30704_));
 DFF_X1 _64137_ (.D(_02944_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2910]),
    .QN(_30705_));
 DFF_X1 _64138_ (.D(_02945_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2911]),
    .QN(_30706_));
 DFF_X1 _64139_ (.D(_02946_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2912]),
    .QN(_30707_));
 DFF_X1 _64140_ (.D(_02947_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2913]),
    .QN(_30708_));
 DFF_X1 _64141_ (.D(_02948_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2914]),
    .QN(_30709_));
 DFF_X1 _64142_ (.D(_02949_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2915]),
    .QN(_30710_));
 DFF_X1 _64143_ (.D(_02950_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2916]),
    .QN(_30711_));
 DFF_X1 _64144_ (.D(_02951_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2917]),
    .QN(_30712_));
 DFF_X1 _64145_ (.D(_02952_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2918]),
    .QN(_30713_));
 DFF_X1 _64146_ (.D(_02953_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2919]),
    .QN(_30714_));
 DFF_X1 _64147_ (.D(_02955_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2920]),
    .QN(_30715_));
 DFF_X1 _64148_ (.D(_02956_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2921]),
    .QN(_30716_));
 DFF_X1 _64149_ (.D(_02957_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2922]),
    .QN(_30717_));
 DFF_X1 _64150_ (.D(_02958_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2923]),
    .QN(_30718_));
 DFF_X1 _64151_ (.D(_02959_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2924]),
    .QN(_30719_));
 DFF_X1 _64152_ (.D(_02960_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2925]),
    .QN(_30720_));
 DFF_X1 _64153_ (.D(_02961_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2926]),
    .QN(_30721_));
 DFF_X1 _64154_ (.D(_02962_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2927]),
    .QN(_30722_));
 DFF_X1 _64155_ (.D(_02963_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2928]),
    .QN(_30723_));
 DFF_X1 _64156_ (.D(_02964_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2929]),
    .QN(_30724_));
 DFF_X1 _64157_ (.D(_02966_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2930]),
    .QN(_30725_));
 DFF_X1 _64158_ (.D(_02967_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2931]),
    .QN(_30726_));
 DFF_X1 _64159_ (.D(_02968_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2932]),
    .QN(_30727_));
 DFF_X1 _64160_ (.D(_02969_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2933]),
    .QN(_30728_));
 DFF_X1 _64161_ (.D(_02970_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2934]),
    .QN(_30729_));
 DFF_X1 _64162_ (.D(_02971_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2935]),
    .QN(_30730_));
 DFF_X1 _64163_ (.D(_02972_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2936]),
    .QN(_30731_));
 DFF_X1 _64164_ (.D(_02973_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2937]),
    .QN(_30732_));
 DFF_X1 _64165_ (.D(_02974_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2938]),
    .QN(_30733_));
 DFF_X1 _64166_ (.D(_02975_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2939]),
    .QN(_30734_));
 DFF_X1 _64167_ (.D(_02977_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2940]),
    .QN(_30735_));
 DFF_X1 _64168_ (.D(_02978_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2941]),
    .QN(_30736_));
 DFF_X1 _64169_ (.D(_02979_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2942]),
    .QN(_30737_));
 DFF_X1 _64170_ (.D(_02980_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2943]),
    .QN(_30738_));
 DFF_X1 _64171_ (.D(_02981_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2944]),
    .QN(_30739_));
 DFF_X1 _64172_ (.D(_02982_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2945]),
    .QN(_30740_));
 DFF_X1 _64173_ (.D(_02983_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2946]),
    .QN(_30741_));
 DFF_X1 _64174_ (.D(_02984_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2947]),
    .QN(_30742_));
 DFF_X1 _64175_ (.D(_02985_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2948]),
    .QN(_30743_));
 DFF_X1 _64176_ (.D(_02986_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2949]),
    .QN(_30744_));
 DFF_X1 _64177_ (.D(_02988_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2950]),
    .QN(_30745_));
 DFF_X1 _64178_ (.D(_02989_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2951]),
    .QN(_30746_));
 DFF_X1 _64179_ (.D(_02990_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2952]),
    .QN(_30747_));
 DFF_X1 _64180_ (.D(_02991_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2953]),
    .QN(_30748_));
 DFF_X1 _64181_ (.D(_02992_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2954]),
    .QN(_30749_));
 DFF_X1 _64182_ (.D(_02993_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2955]),
    .QN(_30750_));
 DFF_X1 _64183_ (.D(_02994_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2956]),
    .QN(_30751_));
 DFF_X1 _64184_ (.D(_02995_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2957]),
    .QN(_30752_));
 DFF_X1 _64185_ (.D(_02996_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2958]),
    .QN(_30753_));
 DFF_X1 _64186_ (.D(_02997_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2959]),
    .QN(_30754_));
 DFF_X1 _64187_ (.D(_02999_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2960]),
    .QN(_30755_));
 DFF_X1 _64188_ (.D(_03000_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2961]),
    .QN(_30756_));
 DFF_X1 _64189_ (.D(_03001_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2962]),
    .QN(_30757_));
 DFF_X1 _64190_ (.D(_03002_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2963]),
    .QN(_30758_));
 DFF_X1 _64191_ (.D(_03003_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2964]),
    .QN(_30759_));
 DFF_X1 _64192_ (.D(_03004_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2965]),
    .QN(_30760_));
 DFF_X1 _64193_ (.D(_03005_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2966]),
    .QN(_30761_));
 DFF_X1 _64194_ (.D(_03006_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2967]),
    .QN(_30762_));
 DFF_X1 _64195_ (.D(_03007_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2968]),
    .QN(_30763_));
 DFF_X1 _64196_ (.D(_03008_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2969]),
    .QN(_30764_));
 DFF_X1 _64197_ (.D(_03010_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2970]),
    .QN(_30765_));
 DFF_X1 _64198_ (.D(_03011_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2971]),
    .QN(_30766_));
 DFF_X1 _64199_ (.D(_03012_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2972]),
    .QN(_30767_));
 DFF_X1 _64200_ (.D(_03013_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2973]),
    .QN(_30768_));
 DFF_X1 _64201_ (.D(_03014_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2974]),
    .QN(_30769_));
 DFF_X1 _64202_ (.D(_03015_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2975]),
    .QN(_30770_));
 DFF_X1 _64203_ (.D(_03016_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2976]),
    .QN(_30771_));
 DFF_X1 _64204_ (.D(_03017_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2977]),
    .QN(_30772_));
 DFF_X1 _64205_ (.D(_03018_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2978]),
    .QN(_30773_));
 DFF_X1 _64206_ (.D(_03019_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2979]),
    .QN(_30774_));
 DFF_X1 _64207_ (.D(_03021_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2980]),
    .QN(_30775_));
 DFF_X1 _64208_ (.D(_03022_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2981]),
    .QN(_30776_));
 DFF_X1 _64209_ (.D(_03023_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2982]),
    .QN(_30777_));
 DFF_X1 _64210_ (.D(_03024_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2983]),
    .QN(_30778_));
 DFF_X1 _64211_ (.D(_03025_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2984]),
    .QN(_30779_));
 DFF_X1 _64212_ (.D(_03026_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2985]),
    .QN(_30780_));
 DFF_X1 _64213_ (.D(_03027_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2986]),
    .QN(_30781_));
 DFF_X1 _64214_ (.D(_03028_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2987]),
    .QN(_30782_));
 DFF_X1 _64215_ (.D(_03029_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2988]),
    .QN(_30783_));
 DFF_X1 _64216_ (.D(_03030_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2989]),
    .QN(_30784_));
 DFF_X1 _64217_ (.D(_03032_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2990]),
    .QN(_30785_));
 DFF_X1 _64218_ (.D(_03033_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2991]),
    .QN(_30786_));
 DFF_X1 _64219_ (.D(_03034_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2992]),
    .QN(_30787_));
 DFF_X1 _64220_ (.D(_03035_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2993]),
    .QN(_30788_));
 DFF_X1 _64221_ (.D(_03036_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2994]),
    .QN(_30789_));
 DFF_X1 _64222_ (.D(_03037_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2995]),
    .QN(_30790_));
 DFF_X1 _64223_ (.D(_03038_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2996]),
    .QN(_30791_));
 DFF_X1 _64224_ (.D(_03039_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2997]),
    .QN(_30792_));
 DFF_X1 _64225_ (.D(_03040_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2998]),
    .QN(_30793_));
 DFF_X1 _64226_ (.D(_03041_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [2999]),
    .QN(_30794_));
 DFF_X1 _64227_ (.D(_03045_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3000]),
    .QN(_30795_));
 DFF_X1 _64228_ (.D(_03046_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3001]),
    .QN(_30796_));
 DFF_X1 _64229_ (.D(_03047_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3002]),
    .QN(_30797_));
 DFF_X1 _64230_ (.D(_03048_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3003]),
    .QN(_30798_));
 DFF_X1 _64231_ (.D(_03049_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3004]),
    .QN(_30799_));
 DFF_X1 _64232_ (.D(_03050_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3005]),
    .QN(_30800_));
 DFF_X1 _64233_ (.D(_03051_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3006]),
    .QN(_30801_));
 DFF_X1 _64234_ (.D(_03052_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3007]),
    .QN(_30802_));
 DFF_X1 _64235_ (.D(_03053_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3008]),
    .QN(_30803_));
 DFF_X1 _64236_ (.D(_03054_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3009]),
    .QN(_30804_));
 DFF_X1 _64237_ (.D(_03056_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3010]),
    .QN(_30805_));
 DFF_X1 _64238_ (.D(_03057_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3011]),
    .QN(_30806_));
 DFF_X1 _64239_ (.D(_03058_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3012]),
    .QN(_30807_));
 DFF_X1 _64240_ (.D(_03059_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3013]),
    .QN(_30808_));
 DFF_X1 _64241_ (.D(_03060_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3014]),
    .QN(_30809_));
 DFF_X1 _64242_ (.D(_03061_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3015]),
    .QN(_30810_));
 DFF_X1 _64243_ (.D(_03062_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3016]),
    .QN(_30811_));
 DFF_X1 _64244_ (.D(_03063_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3017]),
    .QN(_30812_));
 DFF_X1 _64245_ (.D(_03064_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3018]),
    .QN(_30813_));
 DFF_X1 _64246_ (.D(_03065_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3019]),
    .QN(_30814_));
 DFF_X1 _64247_ (.D(_03067_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3020]),
    .QN(_30815_));
 DFF_X1 _64248_ (.D(_03068_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3021]),
    .QN(_30816_));
 DFF_X1 _64249_ (.D(_03069_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3022]),
    .QN(_30817_));
 DFF_X1 _64250_ (.D(_03070_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3023]),
    .QN(_30818_));
 DFF_X1 _64251_ (.D(_03071_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3024]),
    .QN(_30819_));
 DFF_X1 _64252_ (.D(_03072_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3025]),
    .QN(_30820_));
 DFF_X1 _64253_ (.D(_03073_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3026]),
    .QN(_30821_));
 DFF_X1 _64254_ (.D(_03074_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3027]),
    .QN(_30822_));
 DFF_X1 _64255_ (.D(_03075_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3028]),
    .QN(_30823_));
 DFF_X1 _64256_ (.D(_03076_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3029]),
    .QN(_30824_));
 DFF_X1 _64257_ (.D(_03078_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3030]),
    .QN(_30825_));
 DFF_X1 _64258_ (.D(_03079_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3031]),
    .QN(_30826_));
 DFF_X1 _64259_ (.D(_03080_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3032]),
    .QN(_30827_));
 DFF_X1 _64260_ (.D(_03081_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3033]),
    .QN(_30828_));
 DFF_X1 _64261_ (.D(_03082_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3034]),
    .QN(_30829_));
 DFF_X1 _64262_ (.D(_03083_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3035]),
    .QN(_30830_));
 DFF_X1 _64263_ (.D(_03084_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3036]),
    .QN(_30831_));
 DFF_X1 _64264_ (.D(_03085_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3037]),
    .QN(_30832_));
 DFF_X1 _64265_ (.D(_03086_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3038]),
    .QN(_30833_));
 DFF_X1 _64266_ (.D(_03087_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3039]),
    .QN(_30834_));
 DFF_X1 _64267_ (.D(_03089_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3040]),
    .QN(_30835_));
 DFF_X1 _64268_ (.D(_03090_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3041]),
    .QN(_30836_));
 DFF_X1 _64269_ (.D(_03091_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3042]),
    .QN(_30837_));
 DFF_X1 _64270_ (.D(_03092_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3043]),
    .QN(_30838_));
 DFF_X1 _64271_ (.D(_03093_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3044]),
    .QN(_30839_));
 DFF_X1 _64272_ (.D(_03094_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3045]),
    .QN(_30840_));
 DFF_X1 _64273_ (.D(_03095_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3046]),
    .QN(_30841_));
 DFF_X1 _64274_ (.D(_03096_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3047]),
    .QN(_30842_));
 DFF_X1 _64275_ (.D(_03097_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3048]),
    .QN(_30843_));
 DFF_X1 _64276_ (.D(_03098_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3049]),
    .QN(_30844_));
 DFF_X1 _64277_ (.D(_03100_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3050]),
    .QN(_30845_));
 DFF_X1 _64278_ (.D(_03101_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3051]),
    .QN(_30846_));
 DFF_X1 _64279_ (.D(_03102_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3052]),
    .QN(_30847_));
 DFF_X1 _64280_ (.D(_03103_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3053]),
    .QN(_30848_));
 DFF_X1 _64281_ (.D(_03104_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3054]),
    .QN(_30849_));
 DFF_X1 _64282_ (.D(_03105_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3055]),
    .QN(_30850_));
 DFF_X1 _64283_ (.D(_03106_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3056]),
    .QN(_30851_));
 DFF_X1 _64284_ (.D(_03107_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3057]),
    .QN(_30852_));
 DFF_X1 _64285_ (.D(_03108_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3058]),
    .QN(_30853_));
 DFF_X1 _64286_ (.D(_03109_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3059]),
    .QN(_30854_));
 DFF_X1 _64287_ (.D(_03111_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3060]),
    .QN(_30855_));
 DFF_X1 _64288_ (.D(_03112_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3061]),
    .QN(_30856_));
 DFF_X1 _64289_ (.D(_03113_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3062]),
    .QN(_30857_));
 DFF_X1 _64290_ (.D(_03114_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3063]),
    .QN(_30858_));
 DFF_X1 _64291_ (.D(_03115_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3064]),
    .QN(_30859_));
 DFF_X1 _64292_ (.D(_03116_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3065]),
    .QN(_30860_));
 DFF_X1 _64293_ (.D(_03117_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3066]),
    .QN(_30861_));
 DFF_X1 _64294_ (.D(_03118_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3067]),
    .QN(_30862_));
 DFF_X1 _64295_ (.D(_03119_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3068]),
    .QN(_30863_));
 DFF_X1 _64296_ (.D(_03120_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3069]),
    .QN(_30864_));
 DFF_X1 _64297_ (.D(_03122_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3070]),
    .QN(_30865_));
 DFF_X1 _64298_ (.D(_03123_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3071]),
    .QN(_30866_));
 DFF_X1 _64299_ (.D(_03124_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3072]),
    .QN(_30867_));
 DFF_X1 _64300_ (.D(_03125_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3073]),
    .QN(_30868_));
 DFF_X1 _64301_ (.D(_03126_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3074]),
    .QN(_30869_));
 DFF_X1 _64302_ (.D(_03127_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3075]),
    .QN(_30870_));
 DFF_X1 _64303_ (.D(_03128_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3076]),
    .QN(_30871_));
 DFF_X1 _64304_ (.D(_03129_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3077]),
    .QN(_30872_));
 DFF_X1 _64305_ (.D(_03130_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3078]),
    .QN(_30873_));
 DFF_X1 _64306_ (.D(_03131_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3079]),
    .QN(_30874_));
 DFF_X1 _64307_ (.D(_03133_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3080]),
    .QN(_30875_));
 DFF_X1 _64308_ (.D(_03134_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3081]),
    .QN(_30876_));
 DFF_X1 _64309_ (.D(_03135_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3082]),
    .QN(_30877_));
 DFF_X1 _64310_ (.D(_03136_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3083]),
    .QN(_30878_));
 DFF_X1 _64311_ (.D(_03137_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3084]),
    .QN(_30879_));
 DFF_X1 _64312_ (.D(_03138_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3085]),
    .QN(_30880_));
 DFF_X1 _64313_ (.D(_03139_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3086]),
    .QN(_30881_));
 DFF_X1 _64314_ (.D(_03140_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3087]),
    .QN(_30882_));
 DFF_X1 _64315_ (.D(_03141_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3088]),
    .QN(_30883_));
 DFF_X1 _64316_ (.D(_03142_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3089]),
    .QN(_30884_));
 DFF_X1 _64317_ (.D(_03144_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3090]),
    .QN(_30885_));
 DFF_X1 _64318_ (.D(_03145_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3091]),
    .QN(_30886_));
 DFF_X1 _64319_ (.D(_03146_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3092]),
    .QN(_30887_));
 DFF_X1 _64320_ (.D(_03147_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3093]),
    .QN(_30888_));
 DFF_X1 _64321_ (.D(_03148_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3094]),
    .QN(_30889_));
 DFF_X1 _64322_ (.D(_03149_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3095]),
    .QN(_30890_));
 DFF_X1 _64323_ (.D(_03150_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3096]),
    .QN(_30891_));
 DFF_X1 _64324_ (.D(_03151_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3097]),
    .QN(_30892_));
 DFF_X1 _64325_ (.D(_03152_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3098]),
    .QN(_30893_));
 DFF_X1 _64326_ (.D(_03153_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3099]),
    .QN(_30894_));
 DFF_X1 _64327_ (.D(_03156_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3100]),
    .QN(_30895_));
 DFF_X1 _64328_ (.D(_03157_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3101]),
    .QN(_30896_));
 DFF_X1 _64329_ (.D(_03158_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3102]),
    .QN(_30897_));
 DFF_X1 _64330_ (.D(_03159_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3103]),
    .QN(_30898_));
 DFF_X1 _64331_ (.D(_03160_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3104]),
    .QN(_30899_));
 DFF_X1 _64332_ (.D(_03161_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3105]),
    .QN(_30900_));
 DFF_X1 _64333_ (.D(_03162_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3106]),
    .QN(_30901_));
 DFF_X1 _64334_ (.D(_03163_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3107]),
    .QN(_30902_));
 DFF_X1 _64335_ (.D(_03164_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3108]),
    .QN(_30903_));
 DFF_X1 _64336_ (.D(_03165_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3109]),
    .QN(_30904_));
 DFF_X1 _64337_ (.D(_03167_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3110]),
    .QN(_30905_));
 DFF_X1 _64338_ (.D(_03168_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3111]),
    .QN(_30906_));
 DFF_X1 _64339_ (.D(_03169_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3112]),
    .QN(_30907_));
 DFF_X1 _64340_ (.D(_03170_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3113]),
    .QN(_30908_));
 DFF_X1 _64341_ (.D(_03171_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3114]),
    .QN(_30909_));
 DFF_X1 _64342_ (.D(_03172_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3115]),
    .QN(_30910_));
 DFF_X1 _64343_ (.D(_03173_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3116]),
    .QN(_30911_));
 DFF_X1 _64344_ (.D(_03174_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3117]),
    .QN(_30912_));
 DFF_X1 _64345_ (.D(_03175_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3118]),
    .QN(_30913_));
 DFF_X1 _64346_ (.D(_03176_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3119]),
    .QN(_30914_));
 DFF_X1 _64347_ (.D(_03178_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3120]),
    .QN(_30915_));
 DFF_X1 _64348_ (.D(_03179_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3121]),
    .QN(_30916_));
 DFF_X1 _64349_ (.D(_03180_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3122]),
    .QN(_30917_));
 DFF_X1 _64350_ (.D(_03181_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3123]),
    .QN(_30918_));
 DFF_X1 _64351_ (.D(_03182_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3124]),
    .QN(_30919_));
 DFF_X1 _64352_ (.D(_03183_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3125]),
    .QN(_30920_));
 DFF_X1 _64353_ (.D(_03184_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3126]),
    .QN(_30921_));
 DFF_X1 _64354_ (.D(_03185_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3127]),
    .QN(_30922_));
 DFF_X1 _64355_ (.D(_03186_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3128]),
    .QN(_30923_));
 DFF_X1 _64356_ (.D(_03187_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3129]),
    .QN(_30924_));
 DFF_X1 _64357_ (.D(_03189_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3130]),
    .QN(_30925_));
 DFF_X1 _64358_ (.D(_03190_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3131]),
    .QN(_30926_));
 DFF_X1 _64359_ (.D(_03191_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3132]),
    .QN(_30927_));
 DFF_X1 _64360_ (.D(_03192_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3133]),
    .QN(_30928_));
 DFF_X1 _64361_ (.D(_03193_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3134]),
    .QN(_30929_));
 DFF_X1 _64362_ (.D(_03194_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [3135]),
    .QN(_30930_));
 DFF_X1 _64363_ (.D(_05408_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [0]),
    .QN(_30931_));
 DFF_X1 _64364_ (.D(_05424_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [1]),
    .QN(_30932_));
 DFF_X1 _64365_ (.D(_05435_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [2]),
    .QN(_30933_));
 DFF_X1 _64366_ (.D(_05446_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [3]),
    .QN(_30934_));
 DFF_X1 _64367_ (.D(_05457_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [4]),
    .QN(_30935_));
 DFF_X1 _64368_ (.D(_05467_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [5]),
    .QN(_30936_));
 DFF_X1 _64369_ (.D(_05478_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [6]),
    .QN(_30937_));
 DFF_X1 _64370_ (.D(_05489_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [7]),
    .QN(_30938_));
 DFF_X1 _64371_ (.D(_05500_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [8]),
    .QN(_30939_));
 DFF_X1 _64372_ (.D(_05511_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [9]),
    .QN(_00583_));
 DFF_X1 _64373_ (.D(_05414_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [10]),
    .QN(_00585_));
 DFF_X1 _64374_ (.D(_05415_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [11]),
    .QN(_00587_));
 DFF_X1 _64375_ (.D(_05416_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [12]),
    .QN(_00589_));
 DFF_X1 _64376_ (.D(_05417_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [13]),
    .QN(_00591_));
 DFF_X1 _64377_ (.D(_05418_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [14]),
    .QN(_00593_));
 DFF_X1 _64378_ (.D(_05419_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [15]),
    .QN(_30940_));
 DFF_X1 _64379_ (.D(_05420_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [16]),
    .QN(_30941_));
 DFF_X1 _64380_ (.D(_05421_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [17]),
    .QN(_30942_));
 DFF_X1 _64381_ (.D(_05422_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [18]),
    .QN(_30943_));
 DFF_X1 _64382_ (.D(_05423_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [19]),
    .QN(_30944_));
 DFF_X1 _64383_ (.D(_05425_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [20]),
    .QN(_30945_));
 DFF_X1 _64384_ (.D(_05426_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [21]),
    .QN(_30946_));
 DFF_X1 _64385_ (.D(_05427_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [22]),
    .QN(_30947_));
 DFF_X1 _64386_ (.D(_05428_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [23]),
    .QN(_30948_));
 DFF_X1 _64387_ (.D(_05429_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [24]),
    .QN(_30949_));
 DFF_X1 _64388_ (.D(_05430_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [25]),
    .QN(_30950_));
 DFF_X1 _64389_ (.D(_05431_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [26]),
    .QN(_30951_));
 DFF_X1 _64390_ (.D(_05432_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [27]),
    .QN(_30952_));
 DFF_X1 _64391_ (.D(_05433_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [28]),
    .QN(_30953_));
 DFF_X1 _64392_ (.D(_05434_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [29]),
    .QN(_30954_));
 DFF_X1 _64393_ (.D(_05436_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [30]),
    .QN(_30955_));
 DFF_X1 _64394_ (.D(_05437_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [31]),
    .QN(_30956_));
 DFF_X1 _64395_ (.D(_05438_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [32]),
    .QN(_30957_));
 DFF_X1 _64396_ (.D(_05439_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [33]),
    .QN(_30958_));
 DFF_X1 _64397_ (.D(_05440_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [34]),
    .QN(_30959_));
 DFF_X1 _64398_ (.D(_05441_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [35]),
    .QN(_30960_));
 DFF_X1 _64399_ (.D(_05442_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [36]),
    .QN(_30961_));
 DFF_X1 _64400_ (.D(_05443_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [37]),
    .QN(_30962_));
 DFF_X1 _64401_ (.D(_05444_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [38]),
    .QN(_30963_));
 DFF_X1 _64402_ (.D(_05445_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [39]),
    .QN(_30964_));
 DFF_X1 _64403_ (.D(_05447_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [40]),
    .QN(_30965_));
 DFF_X1 _64404_ (.D(_05448_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [41]),
    .QN(_30966_));
 DFF_X1 _64405_ (.D(_05449_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [42]),
    .QN(_30967_));
 DFF_X1 _64406_ (.D(_05450_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [43]),
    .QN(_30968_));
 DFF_X1 _64407_ (.D(_05451_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [44]),
    .QN(_30969_));
 DFF_X1 _64408_ (.D(_05452_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [45]),
    .QN(_30970_));
 DFF_X1 _64409_ (.D(_05453_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [46]),
    .QN(_30971_));
 DFF_X1 _64410_ (.D(_05454_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [47]),
    .QN(_30972_));
 DFF_X1 _64411_ (.D(_05455_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [48]),
    .QN(_30973_));
 DFF_X1 _64412_ (.D(_05456_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [49]),
    .QN(_30974_));
 DFF_X1 _64413_ (.D(_05458_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [50]),
    .QN(_30975_));
 DFF_X1 _64414_ (.D(_05459_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [51]),
    .QN(_00595_));
 DFF_X1 _64415_ (.D(_05460_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [53]),
    .QN(_30976_));
 DFF_X1 _64416_ (.D(_05461_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [54]),
    .QN(_30977_));
 DFF_X1 _64417_ (.D(_05462_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [55]),
    .QN(_30978_));
 DFF_X1 _64418_ (.D(_05463_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [56]),
    .QN(_30979_));
 DFF_X1 _64419_ (.D(_05464_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [57]),
    .QN(_30980_));
 DFF_X1 _64420_ (.D(_05465_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [58]),
    .QN(_30981_));
 DFF_X1 _64421_ (.D(_05466_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [59]),
    .QN(_30982_));
 DFF_X1 _64422_ (.D(_05468_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [60]),
    .QN(_30983_));
 DFF_X1 _64423_ (.D(_05469_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [61]),
    .QN(_30984_));
 DFF_X1 _64424_ (.D(_05470_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [62]),
    .QN(_00584_));
 DFF_X1 _64425_ (.D(_05471_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [63]),
    .QN(_00586_));
 DFF_X1 _64426_ (.D(_05472_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [64]),
    .QN(_00588_));
 DFF_X1 _64427_ (.D(_05473_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [65]),
    .QN(_00590_));
 DFF_X1 _64428_ (.D(_05474_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [66]),
    .QN(_00592_));
 DFF_X1 _64429_ (.D(_05475_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [67]),
    .QN(_00594_));
 DFF_X1 _64430_ (.D(_05476_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [68]),
    .QN(_30985_));
 DFF_X1 _64431_ (.D(_05477_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [69]),
    .QN(_30986_));
 DFF_X1 _64432_ (.D(_05479_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [70]),
    .QN(_30987_));
 DFF_X1 _64433_ (.D(_05480_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [71]),
    .QN(_30988_));
 DFF_X1 _64434_ (.D(_05481_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [72]),
    .QN(_30989_));
 DFF_X1 _64435_ (.D(_05482_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [73]),
    .QN(_30990_));
 DFF_X1 _64436_ (.D(_05483_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [74]),
    .QN(_30991_));
 DFF_X1 _64437_ (.D(_05484_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [75]),
    .QN(_30992_));
 DFF_X1 _64438_ (.D(_05485_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [76]),
    .QN(_30993_));
 DFF_X1 _64439_ (.D(_05486_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [77]),
    .QN(_30994_));
 DFF_X1 _64440_ (.D(_05487_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [78]),
    .QN(_30995_));
 DFF_X1 _64441_ (.D(_05488_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [79]),
    .QN(_30996_));
 DFF_X1 _64442_ (.D(_05490_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [80]),
    .QN(_30997_));
 DFF_X1 _64443_ (.D(_05491_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [81]),
    .QN(_30998_));
 DFF_X1 _64444_ (.D(_05492_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [82]),
    .QN(_30999_));
 DFF_X1 _64445_ (.D(_05493_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [83]),
    .QN(_31000_));
 DFF_X1 _64446_ (.D(_05494_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [84]),
    .QN(_31001_));
 DFF_X1 _64447_ (.D(_05495_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [85]),
    .QN(_31002_));
 DFF_X1 _64448_ (.D(_05496_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [86]),
    .QN(_31003_));
 DFF_X1 _64449_ (.D(_05497_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [87]),
    .QN(_31004_));
 DFF_X1 _64450_ (.D(_05498_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [88]),
    .QN(_31005_));
 DFF_X1 _64451_ (.D(_05499_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [89]),
    .QN(_31006_));
 DFF_X1 _64452_ (.D(_05501_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [90]),
    .QN(_31007_));
 DFF_X1 _64453_ (.D(_05502_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [91]),
    .QN(_31008_));
 DFF_X1 _64454_ (.D(_05503_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [92]),
    .QN(_31009_));
 DFF_X1 _64455_ (.D(_05504_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [93]),
    .QN(_31010_));
 DFF_X1 _64456_ (.D(_05505_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [94]),
    .QN(_31011_));
 DFF_X1 _64457_ (.D(_05506_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [95]),
    .QN(_31012_));
 DFF_X1 _64458_ (.D(_05507_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [96]),
    .QN(_31013_));
 DFF_X1 _64459_ (.D(_05508_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [97]),
    .QN(_31014_));
 DFF_X1 _64460_ (.D(_05509_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [98]),
    .QN(_31015_));
 DFF_X1 _64461_ (.D(_05510_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [99]),
    .QN(_31016_));
 DFF_X1 _64462_ (.D(_05409_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [100]),
    .QN(_31017_));
 DFF_X1 _64463_ (.D(_05410_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [101]),
    .QN(_31018_));
 DFF_X1 _64464_ (.D(_05411_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [102]),
    .QN(_31019_));
 DFF_X1 _64465_ (.D(_05412_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [103]),
    .QN(_31020_));
 DFF_X1 _64466_ (.D(_05413_),
    .CK(clk_i),
    .Q(\icache.lce.lce_cmd_inst.rv_adapter.mem_1r1w.synth.mem [104]),
    .QN(_00596_));
 DFF_X1 _64467_ (.D(_05514_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [0]),
    .QN(_31021_));
 DFF_X1 _64468_ (.D(_05661_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1]),
    .QN(_31022_));
 DFF_X1 _64469_ (.D(_05772_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [2]),
    .QN(_31023_));
 DFF_X1 _64470_ (.D(_05883_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [3]),
    .QN(_31024_));
 DFF_X1 _64471_ (.D(_05994_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [4]),
    .QN(_31025_));
 DFF_X1 _64472_ (.D(_06214_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [6]),
    .QN(_31026_));
 DFF_X1 _64473_ (.D(_06325_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [7]),
    .QN(_31027_));
 DFF_X1 _64474_ (.D(_06436_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [8]),
    .QN(_31028_));
 DFF_X1 _64475_ (.D(_06547_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [9]),
    .QN(_31029_));
 DFF_X1 _64476_ (.D(_05561_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [10]),
    .QN(_31030_));
 DFF_X1 _64477_ (.D(_05572_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [11]),
    .QN(_31031_));
 DFF_X1 _64478_ (.D(_05583_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [12]),
    .QN(_31032_));
 DFF_X1 _64479_ (.D(_05594_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [13]),
    .QN(_31033_));
 DFF_X1 _64480_ (.D(_05605_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [14]),
    .QN(_31034_));
 DFF_X1 _64481_ (.D(_05616_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [15]),
    .QN(_31035_));
 DFF_X1 _64482_ (.D(_05627_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [16]),
    .QN(_31036_));
 DFF_X1 _64483_ (.D(_05638_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [17]),
    .QN(_31037_));
 DFF_X1 _64484_ (.D(_05649_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [18]),
    .QN(_31038_));
 DFF_X1 _64485_ (.D(_05660_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [19]),
    .QN(_31039_));
 DFF_X1 _64486_ (.D(_05672_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [20]),
    .QN(_31040_));
 DFF_X1 _64487_ (.D(_05683_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [21]),
    .QN(_31041_));
 DFF_X1 _64488_ (.D(_05694_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [22]),
    .QN(_31042_));
 DFF_X1 _64489_ (.D(_05705_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [23]),
    .QN(_31043_));
 DFF_X1 _64490_ (.D(_05716_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [24]),
    .QN(_31044_));
 DFF_X1 _64491_ (.D(_05727_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [25]),
    .QN(_31045_));
 DFF_X1 _64492_ (.D(_05738_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [26]),
    .QN(_31046_));
 DFF_X1 _64493_ (.D(_05749_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [27]),
    .QN(_31047_));
 DFF_X1 _64494_ (.D(_05760_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [28]),
    .QN(_31048_));
 DFF_X1 _64495_ (.D(_05771_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [29]),
    .QN(_31049_));
 DFF_X1 _64496_ (.D(_05783_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [30]),
    .QN(_31050_));
 DFF_X1 _64497_ (.D(_05794_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [31]),
    .QN(_31051_));
 DFF_X1 _64498_ (.D(_05805_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [32]),
    .QN(_31052_));
 DFF_X1 _64499_ (.D(_05816_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [33]),
    .QN(_31053_));
 DFF_X1 _64500_ (.D(_05827_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [34]),
    .QN(_31054_));
 DFF_X1 _64501_ (.D(_05838_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [35]),
    .QN(_31055_));
 DFF_X1 _64502_ (.D(_05849_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [36]),
    .QN(_31056_));
 DFF_X1 _64503_ (.D(_05860_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [37]),
    .QN(_31057_));
 DFF_X1 _64504_ (.D(_05871_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [38]),
    .QN(_31058_));
 DFF_X1 _64505_ (.D(_05882_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [39]),
    .QN(_31059_));
 DFF_X1 _64506_ (.D(_05894_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [40]),
    .QN(_31060_));
 DFF_X1 _64507_ (.D(_05905_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [41]),
    .QN(_31061_));
 DFF_X1 _64508_ (.D(_05916_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [42]),
    .QN(_31062_));
 DFF_X1 _64509_ (.D(_05927_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [43]),
    .QN(_31063_));
 DFF_X1 _64510_ (.D(_05938_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [44]),
    .QN(_31064_));
 DFF_X1 _64511_ (.D(_05949_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [45]),
    .QN(_31065_));
 DFF_X1 _64512_ (.D(_05960_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [46]),
    .QN(_31066_));
 DFF_X1 _64513_ (.D(_05971_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [47]),
    .QN(_31067_));
 DFF_X1 _64514_ (.D(_05982_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [48]),
    .QN(_31068_));
 DFF_X1 _64515_ (.D(_05993_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [49]),
    .QN(_31069_));
 DFF_X1 _64516_ (.D(_06005_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [50]),
    .QN(_31070_));
 DFF_X1 _64517_ (.D(_06016_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [51]),
    .QN(_31071_));
 DFF_X1 _64518_ (.D(_06026_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [52]),
    .QN(_31072_));
 DFF_X1 _64519_ (.D(_06037_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [53]),
    .QN(_31073_));
 DFF_X1 _64520_ (.D(_06048_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [54]),
    .QN(_31074_));
 DFF_X1 _64521_ (.D(_06059_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [55]),
    .QN(_31075_));
 DFF_X1 _64522_ (.D(_06070_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [56]),
    .QN(_31076_));
 DFF_X1 _64523_ (.D(_06081_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [57]),
    .QN(_31077_));
 DFF_X1 _64524_ (.D(_06092_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [58]),
    .QN(_31078_));
 DFF_X1 _64525_ (.D(_06103_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [59]),
    .QN(_31079_));
 DFF_X1 _64526_ (.D(_06114_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [60]),
    .QN(_31080_));
 DFF_X1 _64527_ (.D(_06125_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [61]),
    .QN(_31081_));
 DFF_X1 _64528_ (.D(_06136_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [62]),
    .QN(_31082_));
 DFF_X1 _64529_ (.D(_06147_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [63]),
    .QN(_31083_));
 DFF_X1 _64530_ (.D(_06158_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [64]),
    .QN(_31084_));
 DFF_X1 _64531_ (.D(_06169_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [65]),
    .QN(_31085_));
 DFF_X1 _64532_ (.D(_06180_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [66]),
    .QN(_31086_));
 DFF_X1 _64533_ (.D(_06191_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [67]),
    .QN(_31087_));
 DFF_X1 _64534_ (.D(_06202_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [68]),
    .QN(_31088_));
 DFF_X1 _64535_ (.D(_06213_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [69]),
    .QN(_31089_));
 DFF_X1 _64536_ (.D(_06225_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [70]),
    .QN(_31090_));
 DFF_X1 _64537_ (.D(_06236_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [71]),
    .QN(_31091_));
 DFF_X1 _64538_ (.D(_06247_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [72]),
    .QN(_31092_));
 DFF_X1 _64539_ (.D(_06258_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [73]),
    .QN(_31093_));
 DFF_X1 _64540_ (.D(_06269_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [74]),
    .QN(_31094_));
 DFF_X1 _64541_ (.D(_06280_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [75]),
    .QN(_31095_));
 DFF_X1 _64542_ (.D(_06291_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [76]),
    .QN(_31096_));
 DFF_X1 _64543_ (.D(_06302_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [77]),
    .QN(_31097_));
 DFF_X1 _64544_ (.D(_06313_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [78]),
    .QN(_31098_));
 DFF_X1 _64545_ (.D(_06324_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [79]),
    .QN(_31099_));
 DFF_X1 _64546_ (.D(_06336_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [80]),
    .QN(_31100_));
 DFF_X1 _64547_ (.D(_06347_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [81]),
    .QN(_31101_));
 DFF_X1 _64548_ (.D(_06358_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [82]),
    .QN(_31102_));
 DFF_X1 _64549_ (.D(_06369_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [83]),
    .QN(_31103_));
 DFF_X1 _64550_ (.D(_06380_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [84]),
    .QN(_31104_));
 DFF_X1 _64551_ (.D(_06391_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [85]),
    .QN(_31105_));
 DFF_X1 _64552_ (.D(_06402_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [86]),
    .QN(_31106_));
 DFF_X1 _64553_ (.D(_06413_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [87]),
    .QN(_31107_));
 DFF_X1 _64554_ (.D(_06424_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [88]),
    .QN(_31108_));
 DFF_X1 _64555_ (.D(_06435_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [89]),
    .QN(_31109_));
 DFF_X1 _64556_ (.D(_06447_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [90]),
    .QN(_31110_));
 DFF_X1 _64557_ (.D(_06458_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [91]),
    .QN(_31111_));
 DFF_X1 _64558_ (.D(_06469_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [92]),
    .QN(_31112_));
 DFF_X1 _64559_ (.D(_06480_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [93]),
    .QN(_31113_));
 DFF_X1 _64560_ (.D(_06491_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [94]),
    .QN(_31114_));
 DFF_X1 _64561_ (.D(_06502_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [95]),
    .QN(_31115_));
 DFF_X1 _64562_ (.D(_06513_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [96]),
    .QN(_31116_));
 DFF_X1 _64563_ (.D(_06524_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [97]),
    .QN(_31117_));
 DFF_X1 _64564_ (.D(_06535_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [98]),
    .QN(_31118_));
 DFF_X1 _64565_ (.D(_06546_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [99]),
    .QN(_31119_));
 DFF_X1 _64566_ (.D(_05525_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [100]),
    .QN(_31120_));
 DFF_X1 _64567_ (.D(_05536_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [101]),
    .QN(_31121_));
 DFF_X1 _64568_ (.D(_05547_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [102]),
    .QN(_31122_));
 DFF_X1 _64569_ (.D(_05554_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [103]),
    .QN(_31123_));
 DFF_X1 _64570_ (.D(_05555_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [104]),
    .QN(_31124_));
 DFF_X1 _64571_ (.D(_05556_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [105]),
    .QN(_31125_));
 DFF_X1 _64572_ (.D(_05557_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [106]),
    .QN(_31126_));
 DFF_X1 _64573_ (.D(_05558_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [107]),
    .QN(_31127_));
 DFF_X1 _64574_ (.D(_05559_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [108]),
    .QN(_31128_));
 DFF_X1 _64575_ (.D(_05560_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [109]),
    .QN(_31129_));
 DFF_X1 _64576_ (.D(_05562_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [110]),
    .QN(_31130_));
 DFF_X1 _64577_ (.D(_05563_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [111]),
    .QN(_31131_));
 DFF_X1 _64578_ (.D(_05564_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [112]),
    .QN(_31132_));
 DFF_X1 _64579_ (.D(_05565_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [113]),
    .QN(_31133_));
 DFF_X1 _64580_ (.D(_05566_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [114]),
    .QN(_31134_));
 DFF_X1 _64581_ (.D(_05567_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [115]),
    .QN(_31135_));
 DFF_X1 _64582_ (.D(_05568_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [116]),
    .QN(_31136_));
 DFF_X1 _64583_ (.D(_05569_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [117]),
    .QN(_31137_));
 DFF_X1 _64584_ (.D(_05570_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [118]),
    .QN(_31138_));
 DFF_X1 _64585_ (.D(_05571_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [119]),
    .QN(_31139_));
 DFF_X1 _64586_ (.D(_05573_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [120]),
    .QN(_31140_));
 DFF_X1 _64587_ (.D(_05574_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [121]),
    .QN(_31141_));
 DFF_X1 _64588_ (.D(_05575_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [122]),
    .QN(_31142_));
 DFF_X1 _64589_ (.D(_05576_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [123]),
    .QN(_31143_));
 DFF_X1 _64590_ (.D(_05577_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [124]),
    .QN(_31144_));
 DFF_X1 _64591_ (.D(_05578_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [125]),
    .QN(_31145_));
 DFF_X1 _64592_ (.D(_05579_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [126]),
    .QN(_31146_));
 DFF_X1 _64593_ (.D(_05580_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [127]),
    .QN(_31147_));
 DFF_X1 _64594_ (.D(_05581_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [128]),
    .QN(_31148_));
 DFF_X1 _64595_ (.D(_05582_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [129]),
    .QN(_31149_));
 DFF_X1 _64596_ (.D(_05584_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [130]),
    .QN(_31150_));
 DFF_X1 _64597_ (.D(_05585_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [131]),
    .QN(_31151_));
 DFF_X1 _64598_ (.D(_05586_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [132]),
    .QN(_31152_));
 DFF_X1 _64599_ (.D(_05587_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [133]),
    .QN(_31153_));
 DFF_X1 _64600_ (.D(_05588_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [134]),
    .QN(_31154_));
 DFF_X1 _64601_ (.D(_05589_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [135]),
    .QN(_31155_));
 DFF_X1 _64602_ (.D(_05590_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [136]),
    .QN(_31156_));
 DFF_X1 _64603_ (.D(_05591_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [137]),
    .QN(_31157_));
 DFF_X1 _64604_ (.D(_05592_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [138]),
    .QN(_31158_));
 DFF_X1 _64605_ (.D(_05593_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [139]),
    .QN(_31159_));
 DFF_X1 _64606_ (.D(_05595_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [140]),
    .QN(_31160_));
 DFF_X1 _64607_ (.D(_05596_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [141]),
    .QN(_31161_));
 DFF_X1 _64608_ (.D(_05597_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [142]),
    .QN(_31162_));
 DFF_X1 _64609_ (.D(_05598_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [143]),
    .QN(_31163_));
 DFF_X1 _64610_ (.D(_05599_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [144]),
    .QN(_31164_));
 DFF_X1 _64611_ (.D(_05600_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [145]),
    .QN(_31165_));
 DFF_X1 _64612_ (.D(_05601_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [146]),
    .QN(_31166_));
 DFF_X1 _64613_ (.D(_05602_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [147]),
    .QN(_31167_));
 DFF_X1 _64614_ (.D(_05603_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [148]),
    .QN(_31168_));
 DFF_X1 _64615_ (.D(_05604_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [149]),
    .QN(_31169_));
 DFF_X1 _64616_ (.D(_05606_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [150]),
    .QN(_31170_));
 DFF_X1 _64617_ (.D(_05607_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [151]),
    .QN(_31171_));
 DFF_X1 _64618_ (.D(_05608_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [152]),
    .QN(_31172_));
 DFF_X1 _64619_ (.D(_05609_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [153]),
    .QN(_31173_));
 DFF_X1 _64620_ (.D(_05610_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [154]),
    .QN(_31174_));
 DFF_X1 _64621_ (.D(_05611_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [155]),
    .QN(_31175_));
 DFF_X1 _64622_ (.D(_05612_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [156]),
    .QN(_31176_));
 DFF_X1 _64623_ (.D(_05613_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [157]),
    .QN(_31177_));
 DFF_X1 _64624_ (.D(_05614_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [158]),
    .QN(_31178_));
 DFF_X1 _64625_ (.D(_05615_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [159]),
    .QN(_31179_));
 DFF_X1 _64626_ (.D(_05617_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [160]),
    .QN(_31180_));
 DFF_X1 _64627_ (.D(_05618_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [161]),
    .QN(_31181_));
 DFF_X1 _64628_ (.D(_05619_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [162]),
    .QN(_31182_));
 DFF_X1 _64629_ (.D(_05620_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [163]),
    .QN(_31183_));
 DFF_X1 _64630_ (.D(_05621_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [164]),
    .QN(_31184_));
 DFF_X1 _64631_ (.D(_05622_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [165]),
    .QN(_31185_));
 DFF_X1 _64632_ (.D(_05623_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [166]),
    .QN(_31186_));
 DFF_X1 _64633_ (.D(_05624_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [167]),
    .QN(_31187_));
 DFF_X1 _64634_ (.D(_05625_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [168]),
    .QN(_31188_));
 DFF_X1 _64635_ (.D(_05626_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [169]),
    .QN(_31189_));
 DFF_X1 _64636_ (.D(_05628_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [170]),
    .QN(_31190_));
 DFF_X1 _64637_ (.D(_05629_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [171]),
    .QN(_31191_));
 DFF_X1 _64638_ (.D(_05630_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [172]),
    .QN(_31192_));
 DFF_X1 _64639_ (.D(_05631_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [173]),
    .QN(_31193_));
 DFF_X1 _64640_ (.D(_05632_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [174]),
    .QN(_31194_));
 DFF_X1 _64641_ (.D(_05633_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [175]),
    .QN(_31195_));
 DFF_X1 _64642_ (.D(_05634_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [176]),
    .QN(_31196_));
 DFF_X1 _64643_ (.D(_05635_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [177]),
    .QN(_31197_));
 DFF_X1 _64644_ (.D(_05636_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [178]),
    .QN(_31198_));
 DFF_X1 _64645_ (.D(_05637_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [179]),
    .QN(_31199_));
 DFF_X1 _64646_ (.D(_05639_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [180]),
    .QN(_31200_));
 DFF_X1 _64647_ (.D(_05640_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [181]),
    .QN(_31201_));
 DFF_X1 _64648_ (.D(_05641_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [182]),
    .QN(_31202_));
 DFF_X1 _64649_ (.D(_05642_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [183]),
    .QN(_31203_));
 DFF_X1 _64650_ (.D(_05643_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [184]),
    .QN(_31204_));
 DFF_X1 _64651_ (.D(_05644_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [185]),
    .QN(_31205_));
 DFF_X1 _64652_ (.D(_05645_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [186]),
    .QN(_31206_));
 DFF_X1 _64653_ (.D(_05646_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [187]),
    .QN(_31207_));
 DFF_X1 _64654_ (.D(_05647_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [188]),
    .QN(_31208_));
 DFF_X1 _64655_ (.D(_05648_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [189]),
    .QN(_31209_));
 DFF_X1 _64656_ (.D(_05650_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [190]),
    .QN(_31210_));
 DFF_X1 _64657_ (.D(_05651_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [191]),
    .QN(_31211_));
 DFF_X1 _64658_ (.D(_05652_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [192]),
    .QN(_31212_));
 DFF_X1 _64659_ (.D(_05653_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [193]),
    .QN(_31213_));
 DFF_X1 _64660_ (.D(_05654_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [194]),
    .QN(_31214_));
 DFF_X1 _64661_ (.D(_05655_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [195]),
    .QN(_31215_));
 DFF_X1 _64662_ (.D(_05656_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [196]),
    .QN(_31216_));
 DFF_X1 _64663_ (.D(_05657_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [197]),
    .QN(_31217_));
 DFF_X1 _64664_ (.D(_05658_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [198]),
    .QN(_31218_));
 DFF_X1 _64665_ (.D(_05659_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [199]),
    .QN(_31219_));
 DFF_X1 _64666_ (.D(_05662_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [200]),
    .QN(_31220_));
 DFF_X1 _64667_ (.D(_05663_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [201]),
    .QN(_31221_));
 DFF_X1 _64668_ (.D(_05664_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [202]),
    .QN(_31222_));
 DFF_X1 _64669_ (.D(_05665_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [203]),
    .QN(_31223_));
 DFF_X1 _64670_ (.D(_05666_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [204]),
    .QN(_31224_));
 DFF_X1 _64671_ (.D(_05667_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [205]),
    .QN(_31225_));
 DFF_X1 _64672_ (.D(_05668_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [206]),
    .QN(_31226_));
 DFF_X1 _64673_ (.D(_05669_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [207]),
    .QN(_31227_));
 DFF_X1 _64674_ (.D(_05670_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [208]),
    .QN(_31228_));
 DFF_X1 _64675_ (.D(_05671_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [209]),
    .QN(_31229_));
 DFF_X1 _64676_ (.D(_05673_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [210]),
    .QN(_31230_));
 DFF_X1 _64677_ (.D(_05674_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [211]),
    .QN(_31231_));
 DFF_X1 _64678_ (.D(_05675_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [212]),
    .QN(_31232_));
 DFF_X1 _64679_ (.D(_05676_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [213]),
    .QN(_31233_));
 DFF_X1 _64680_ (.D(_05677_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [214]),
    .QN(_31234_));
 DFF_X1 _64681_ (.D(_05678_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [215]),
    .QN(_31235_));
 DFF_X1 _64682_ (.D(_05679_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [216]),
    .QN(_31236_));
 DFF_X1 _64683_ (.D(_05680_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [217]),
    .QN(_31237_));
 DFF_X1 _64684_ (.D(_05681_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [218]),
    .QN(_31238_));
 DFF_X1 _64685_ (.D(_05682_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [219]),
    .QN(_31239_));
 DFF_X1 _64686_ (.D(_05684_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [220]),
    .QN(_31240_));
 DFF_X1 _64687_ (.D(_05685_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [221]),
    .QN(_31241_));
 DFF_X1 _64688_ (.D(_05686_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [222]),
    .QN(_31242_));
 DFF_X1 _64689_ (.D(_05687_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [223]),
    .QN(_31243_));
 DFF_X1 _64690_ (.D(_05688_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [224]),
    .QN(_31244_));
 DFF_X1 _64691_ (.D(_05689_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [225]),
    .QN(_31245_));
 DFF_X1 _64692_ (.D(_05690_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [226]),
    .QN(_31246_));
 DFF_X1 _64693_ (.D(_05691_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [227]),
    .QN(_31247_));
 DFF_X1 _64694_ (.D(_05692_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [228]),
    .QN(_31248_));
 DFF_X1 _64695_ (.D(_05693_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [229]),
    .QN(_31249_));
 DFF_X1 _64696_ (.D(_05695_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [230]),
    .QN(_31250_));
 DFF_X1 _64697_ (.D(_05696_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [231]),
    .QN(_31251_));
 DFF_X1 _64698_ (.D(_05697_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [232]),
    .QN(_31252_));
 DFF_X1 _64699_ (.D(_05698_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [233]),
    .QN(_31253_));
 DFF_X1 _64700_ (.D(_05699_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [234]),
    .QN(_31254_));
 DFF_X1 _64701_ (.D(_05700_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [235]),
    .QN(_31255_));
 DFF_X1 _64702_ (.D(_05701_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [236]),
    .QN(_31256_));
 DFF_X1 _64703_ (.D(_05702_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [237]),
    .QN(_31257_));
 DFF_X1 _64704_ (.D(_05703_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [238]),
    .QN(_31258_));
 DFF_X1 _64705_ (.D(_05704_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [239]),
    .QN(_31259_));
 DFF_X1 _64706_ (.D(_05706_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [240]),
    .QN(_31260_));
 DFF_X1 _64707_ (.D(_05707_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [241]),
    .QN(_31261_));
 DFF_X1 _64708_ (.D(_05708_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [242]),
    .QN(_31262_));
 DFF_X1 _64709_ (.D(_05709_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [243]),
    .QN(_31263_));
 DFF_X1 _64710_ (.D(_05710_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [244]),
    .QN(_31264_));
 DFF_X1 _64711_ (.D(_05711_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [245]),
    .QN(_31265_));
 DFF_X1 _64712_ (.D(_05712_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [246]),
    .QN(_31266_));
 DFF_X1 _64713_ (.D(_05713_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [247]),
    .QN(_31267_));
 DFF_X1 _64714_ (.D(_05714_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [248]),
    .QN(_31268_));
 DFF_X1 _64715_ (.D(_05715_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [249]),
    .QN(_31269_));
 DFF_X1 _64716_ (.D(_05717_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [250]),
    .QN(_31270_));
 DFF_X1 _64717_ (.D(_05718_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [251]),
    .QN(_31271_));
 DFF_X1 _64718_ (.D(_05719_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [252]),
    .QN(_31272_));
 DFF_X1 _64719_ (.D(_05720_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [253]),
    .QN(_31273_));
 DFF_X1 _64720_ (.D(_05721_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [254]),
    .QN(_31274_));
 DFF_X1 _64721_ (.D(_05722_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [255]),
    .QN(_31275_));
 DFF_X1 _64722_ (.D(_05723_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [256]),
    .QN(_31276_));
 DFF_X1 _64723_ (.D(_05724_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [257]),
    .QN(_31277_));
 DFF_X1 _64724_ (.D(_05725_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [258]),
    .QN(_31278_));
 DFF_X1 _64725_ (.D(_05726_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [259]),
    .QN(_31279_));
 DFF_X1 _64726_ (.D(_05728_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [260]),
    .QN(_31280_));
 DFF_X1 _64727_ (.D(_05729_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [261]),
    .QN(_31281_));
 DFF_X1 _64728_ (.D(_05730_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [262]),
    .QN(_31282_));
 DFF_X1 _64729_ (.D(_05731_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [263]),
    .QN(_31283_));
 DFF_X1 _64730_ (.D(_05732_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [264]),
    .QN(_31284_));
 DFF_X1 _64731_ (.D(_05733_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [265]),
    .QN(_31285_));
 DFF_X1 _64732_ (.D(_05734_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [266]),
    .QN(_31286_));
 DFF_X1 _64733_ (.D(_05735_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [267]),
    .QN(_31287_));
 DFF_X1 _64734_ (.D(_05736_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [268]),
    .QN(_31288_));
 DFF_X1 _64735_ (.D(_05737_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [269]),
    .QN(_31289_));
 DFF_X1 _64736_ (.D(_05739_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [270]),
    .QN(_31290_));
 DFF_X1 _64737_ (.D(_05740_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [271]),
    .QN(_31291_));
 DFF_X1 _64738_ (.D(_05741_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [272]),
    .QN(_31292_));
 DFF_X1 _64739_ (.D(_05742_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [273]),
    .QN(_31293_));
 DFF_X1 _64740_ (.D(_05743_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [274]),
    .QN(_31294_));
 DFF_X1 _64741_ (.D(_05744_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [275]),
    .QN(_31295_));
 DFF_X1 _64742_ (.D(_05745_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [276]),
    .QN(_31296_));
 DFF_X1 _64743_ (.D(_05746_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [277]),
    .QN(_31297_));
 DFF_X1 _64744_ (.D(_05747_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [278]),
    .QN(_31298_));
 DFF_X1 _64745_ (.D(_05748_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [279]),
    .QN(_31299_));
 DFF_X1 _64746_ (.D(_05750_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [280]),
    .QN(_31300_));
 DFF_X1 _64747_ (.D(_05751_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [281]),
    .QN(_31301_));
 DFF_X1 _64748_ (.D(_05752_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [282]),
    .QN(_31302_));
 DFF_X1 _64749_ (.D(_05753_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [283]),
    .QN(_31303_));
 DFF_X1 _64750_ (.D(_05754_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [284]),
    .QN(_31304_));
 DFF_X1 _64751_ (.D(_05755_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [285]),
    .QN(_31305_));
 DFF_X1 _64752_ (.D(_05756_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [286]),
    .QN(_31306_));
 DFF_X1 _64753_ (.D(_05757_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [287]),
    .QN(_31307_));
 DFF_X1 _64754_ (.D(_05758_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [288]),
    .QN(_31308_));
 DFF_X1 _64755_ (.D(_05759_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [289]),
    .QN(_31309_));
 DFF_X1 _64756_ (.D(_05761_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [290]),
    .QN(_31310_));
 DFF_X1 _64757_ (.D(_05762_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [291]),
    .QN(_31311_));
 DFF_X1 _64758_ (.D(_05763_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [292]),
    .QN(_31312_));
 DFF_X1 _64759_ (.D(_05764_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [293]),
    .QN(_31313_));
 DFF_X1 _64760_ (.D(_05765_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [294]),
    .QN(_31314_));
 DFF_X1 _64761_ (.D(_05766_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [295]),
    .QN(_31315_));
 DFF_X1 _64762_ (.D(_05767_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [296]),
    .QN(_31316_));
 DFF_X1 _64763_ (.D(_05768_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [297]),
    .QN(_31317_));
 DFF_X1 _64764_ (.D(_05769_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [298]),
    .QN(_31318_));
 DFF_X1 _64765_ (.D(_05770_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [299]),
    .QN(_31319_));
 DFF_X1 _64766_ (.D(_05773_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [300]),
    .QN(_31320_));
 DFF_X1 _64767_ (.D(_05774_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [301]),
    .QN(_31321_));
 DFF_X1 _64768_ (.D(_05775_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [302]),
    .QN(_31322_));
 DFF_X1 _64769_ (.D(_05776_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [303]),
    .QN(_31323_));
 DFF_X1 _64770_ (.D(_05777_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [304]),
    .QN(_31324_));
 DFF_X1 _64771_ (.D(_05778_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [305]),
    .QN(_31325_));
 DFF_X1 _64772_ (.D(_05779_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [306]),
    .QN(_31326_));
 DFF_X1 _64773_ (.D(_05780_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [307]),
    .QN(_31327_));
 DFF_X1 _64774_ (.D(_05781_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [308]),
    .QN(_31328_));
 DFF_X1 _64775_ (.D(_05782_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [309]),
    .QN(_31329_));
 DFF_X1 _64776_ (.D(_05784_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [310]),
    .QN(_31330_));
 DFF_X1 _64777_ (.D(_05785_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [311]),
    .QN(_31331_));
 DFF_X1 _64778_ (.D(_05786_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [312]),
    .QN(_31332_));
 DFF_X1 _64779_ (.D(_05787_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [313]),
    .QN(_31333_));
 DFF_X1 _64780_ (.D(_05788_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [314]),
    .QN(_31334_));
 DFF_X1 _64781_ (.D(_05789_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [315]),
    .QN(_31335_));
 DFF_X1 _64782_ (.D(_05790_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [316]),
    .QN(_31336_));
 DFF_X1 _64783_ (.D(_05791_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [317]),
    .QN(_31337_));
 DFF_X1 _64784_ (.D(_05792_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [318]),
    .QN(_31338_));
 DFF_X1 _64785_ (.D(_05793_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [319]),
    .QN(_31339_));
 DFF_X1 _64786_ (.D(_05795_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [320]),
    .QN(_31340_));
 DFF_X1 _64787_ (.D(_05796_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [321]),
    .QN(_31341_));
 DFF_X1 _64788_ (.D(_05797_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [322]),
    .QN(_31342_));
 DFF_X1 _64789_ (.D(_05798_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [323]),
    .QN(_31343_));
 DFF_X1 _64790_ (.D(_05799_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [324]),
    .QN(_31344_));
 DFF_X1 _64791_ (.D(_05800_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [325]),
    .QN(_31345_));
 DFF_X1 _64792_ (.D(_05801_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [326]),
    .QN(_31346_));
 DFF_X1 _64793_ (.D(_05802_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [327]),
    .QN(_31347_));
 DFF_X1 _64794_ (.D(_05803_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [328]),
    .QN(_31348_));
 DFF_X1 _64795_ (.D(_05804_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [329]),
    .QN(_31349_));
 DFF_X1 _64796_ (.D(_05806_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [330]),
    .QN(_31350_));
 DFF_X1 _64797_ (.D(_05807_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [331]),
    .QN(_31351_));
 DFF_X1 _64798_ (.D(_05808_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [332]),
    .QN(_31352_));
 DFF_X1 _64799_ (.D(_05809_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [333]),
    .QN(_31353_));
 DFF_X1 _64800_ (.D(_05810_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [334]),
    .QN(_31354_));
 DFF_X1 _64801_ (.D(_05811_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [335]),
    .QN(_31355_));
 DFF_X1 _64802_ (.D(_05812_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [336]),
    .QN(_31356_));
 DFF_X1 _64803_ (.D(_05813_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [337]),
    .QN(_31357_));
 DFF_X1 _64804_ (.D(_05814_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [338]),
    .QN(_31358_));
 DFF_X1 _64805_ (.D(_05815_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [339]),
    .QN(_31359_));
 DFF_X1 _64806_ (.D(_05817_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [340]),
    .QN(_31360_));
 DFF_X1 _64807_ (.D(_05818_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [341]),
    .QN(_31361_));
 DFF_X1 _64808_ (.D(_05819_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [342]),
    .QN(_31362_));
 DFF_X1 _64809_ (.D(_05820_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [343]),
    .QN(_31363_));
 DFF_X1 _64810_ (.D(_05821_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [344]),
    .QN(_31364_));
 DFF_X1 _64811_ (.D(_05822_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [345]),
    .QN(_31365_));
 DFF_X1 _64812_ (.D(_05823_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [346]),
    .QN(_31366_));
 DFF_X1 _64813_ (.D(_05824_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [347]),
    .QN(_31367_));
 DFF_X1 _64814_ (.D(_05825_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [348]),
    .QN(_31368_));
 DFF_X1 _64815_ (.D(_05826_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [349]),
    .QN(_31369_));
 DFF_X1 _64816_ (.D(_05828_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [350]),
    .QN(_31370_));
 DFF_X1 _64817_ (.D(_05829_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [351]),
    .QN(_31371_));
 DFF_X1 _64818_ (.D(_05830_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [352]),
    .QN(_31372_));
 DFF_X1 _64819_ (.D(_05831_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [353]),
    .QN(_31373_));
 DFF_X1 _64820_ (.D(_05832_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [354]),
    .QN(_31374_));
 DFF_X1 _64821_ (.D(_05833_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [355]),
    .QN(_31375_));
 DFF_X1 _64822_ (.D(_05834_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [356]),
    .QN(_31376_));
 DFF_X1 _64823_ (.D(_05835_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [357]),
    .QN(_31377_));
 DFF_X1 _64824_ (.D(_05836_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [358]),
    .QN(_31378_));
 DFF_X1 _64825_ (.D(_05837_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [359]),
    .QN(_31379_));
 DFF_X1 _64826_ (.D(_05839_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [360]),
    .QN(_31380_));
 DFF_X1 _64827_ (.D(_05840_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [361]),
    .QN(_31381_));
 DFF_X1 _64828_ (.D(_05841_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [362]),
    .QN(_31382_));
 DFF_X1 _64829_ (.D(_05842_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [363]),
    .QN(_31383_));
 DFF_X1 _64830_ (.D(_05843_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [364]),
    .QN(_31384_));
 DFF_X1 _64831_ (.D(_05844_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [365]),
    .QN(_31385_));
 DFF_X1 _64832_ (.D(_05845_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [366]),
    .QN(_31386_));
 DFF_X1 _64833_ (.D(_05846_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [367]),
    .QN(_31387_));
 DFF_X1 _64834_ (.D(_05847_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [368]),
    .QN(_31388_));
 DFF_X1 _64835_ (.D(_05848_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [369]),
    .QN(_31389_));
 DFF_X1 _64836_ (.D(_05850_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [370]),
    .QN(_31390_));
 DFF_X1 _64837_ (.D(_05851_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [371]),
    .QN(_31391_));
 DFF_X1 _64838_ (.D(_05852_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [372]),
    .QN(_31392_));
 DFF_X1 _64839_ (.D(_05853_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [373]),
    .QN(_31393_));
 DFF_X1 _64840_ (.D(_05854_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [374]),
    .QN(_31394_));
 DFF_X1 _64841_ (.D(_05855_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [375]),
    .QN(_31395_));
 DFF_X1 _64842_ (.D(_05856_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [376]),
    .QN(_31396_));
 DFF_X1 _64843_ (.D(_05857_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [377]),
    .QN(_31397_));
 DFF_X1 _64844_ (.D(_05858_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [378]),
    .QN(_31398_));
 DFF_X1 _64845_ (.D(_05859_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [379]),
    .QN(_31399_));
 DFF_X1 _64846_ (.D(_05861_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [380]),
    .QN(_31400_));
 DFF_X1 _64847_ (.D(_05862_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [381]),
    .QN(_31401_));
 DFF_X1 _64848_ (.D(_05863_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [382]),
    .QN(_31402_));
 DFF_X1 _64849_ (.D(_05864_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [383]),
    .QN(_31403_));
 DFF_X1 _64850_ (.D(_05865_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [384]),
    .QN(_31404_));
 DFF_X1 _64851_ (.D(_05866_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [385]),
    .QN(_31405_));
 DFF_X1 _64852_ (.D(_05867_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [386]),
    .QN(_31406_));
 DFF_X1 _64853_ (.D(_05868_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [387]),
    .QN(_31407_));
 DFF_X1 _64854_ (.D(_05869_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [388]),
    .QN(_31408_));
 DFF_X1 _64855_ (.D(_05870_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [389]),
    .QN(_31409_));
 DFF_X1 _64856_ (.D(_05872_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [390]),
    .QN(_31410_));
 DFF_X1 _64857_ (.D(_05873_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [391]),
    .QN(_31411_));
 DFF_X1 _64858_ (.D(_05874_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [392]),
    .QN(_31412_));
 DFF_X1 _64859_ (.D(_05875_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [393]),
    .QN(_31413_));
 DFF_X1 _64860_ (.D(_05876_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [394]),
    .QN(_31414_));
 DFF_X1 _64861_ (.D(_05877_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [395]),
    .QN(_31415_));
 DFF_X1 _64862_ (.D(_05878_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [396]),
    .QN(_31416_));
 DFF_X1 _64863_ (.D(_05879_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [397]),
    .QN(_31417_));
 DFF_X1 _64864_ (.D(_05880_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [398]),
    .QN(_31418_));
 DFF_X1 _64865_ (.D(_05881_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [399]),
    .QN(_31419_));
 DFF_X1 _64866_ (.D(_05884_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [400]),
    .QN(_31420_));
 DFF_X1 _64867_ (.D(_05885_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [401]),
    .QN(_31421_));
 DFF_X1 _64868_ (.D(_05886_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [402]),
    .QN(_31422_));
 DFF_X1 _64869_ (.D(_05887_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [403]),
    .QN(_31423_));
 DFF_X1 _64870_ (.D(_05888_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [404]),
    .QN(_31424_));
 DFF_X1 _64871_ (.D(_05889_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [405]),
    .QN(_31425_));
 DFF_X1 _64872_ (.D(_05890_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [406]),
    .QN(_31426_));
 DFF_X1 _64873_ (.D(_05891_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [407]),
    .QN(_31427_));
 DFF_X1 _64874_ (.D(_05892_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [408]),
    .QN(_31428_));
 DFF_X1 _64875_ (.D(_05893_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [409]),
    .QN(_31429_));
 DFF_X1 _64876_ (.D(_05895_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [410]),
    .QN(_31430_));
 DFF_X1 _64877_ (.D(_05896_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [411]),
    .QN(_31431_));
 DFF_X1 _64878_ (.D(_05897_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [412]),
    .QN(_31432_));
 DFF_X1 _64879_ (.D(_05898_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [413]),
    .QN(_31433_));
 DFF_X1 _64880_ (.D(_05899_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [414]),
    .QN(_31434_));
 DFF_X1 _64881_ (.D(_05900_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [415]),
    .QN(_31435_));
 DFF_X1 _64882_ (.D(_05901_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [416]),
    .QN(_31436_));
 DFF_X1 _64883_ (.D(_05902_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [417]),
    .QN(_31437_));
 DFF_X1 _64884_ (.D(_05903_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [418]),
    .QN(_31438_));
 DFF_X1 _64885_ (.D(_05904_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [419]),
    .QN(_31439_));
 DFF_X1 _64886_ (.D(_05906_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [420]),
    .QN(_31440_));
 DFF_X1 _64887_ (.D(_05907_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [421]),
    .QN(_31441_));
 DFF_X1 _64888_ (.D(_05908_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [422]),
    .QN(_31442_));
 DFF_X1 _64889_ (.D(_05909_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [423]),
    .QN(_31443_));
 DFF_X1 _64890_ (.D(_05910_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [424]),
    .QN(_31444_));
 DFF_X1 _64891_ (.D(_05911_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [425]),
    .QN(_31445_));
 DFF_X1 _64892_ (.D(_05912_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [426]),
    .QN(_31446_));
 DFF_X1 _64893_ (.D(_05913_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [427]),
    .QN(_31447_));
 DFF_X1 _64894_ (.D(_05914_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [428]),
    .QN(_31448_));
 DFF_X1 _64895_ (.D(_05915_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [429]),
    .QN(_31449_));
 DFF_X1 _64896_ (.D(_05917_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [430]),
    .QN(_31450_));
 DFF_X1 _64897_ (.D(_05918_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [431]),
    .QN(_31451_));
 DFF_X1 _64898_ (.D(_05919_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [432]),
    .QN(_31452_));
 DFF_X1 _64899_ (.D(_05920_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [433]),
    .QN(_31453_));
 DFF_X1 _64900_ (.D(_05921_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [434]),
    .QN(_31454_));
 DFF_X1 _64901_ (.D(_05922_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [435]),
    .QN(_31455_));
 DFF_X1 _64902_ (.D(_05923_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [436]),
    .QN(_31456_));
 DFF_X1 _64903_ (.D(_05924_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [437]),
    .QN(_31457_));
 DFF_X1 _64904_ (.D(_05925_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [438]),
    .QN(_31458_));
 DFF_X1 _64905_ (.D(_05926_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [439]),
    .QN(_31459_));
 DFF_X1 _64906_ (.D(_05928_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [440]),
    .QN(_31460_));
 DFF_X1 _64907_ (.D(_05929_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [441]),
    .QN(_31461_));
 DFF_X1 _64908_ (.D(_05930_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [442]),
    .QN(_31462_));
 DFF_X1 _64909_ (.D(_05931_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [443]),
    .QN(_31463_));
 DFF_X1 _64910_ (.D(_05932_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [444]),
    .QN(_31464_));
 DFF_X1 _64911_ (.D(_05933_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [445]),
    .QN(_31465_));
 DFF_X1 _64912_ (.D(_05934_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [446]),
    .QN(_31466_));
 DFF_X1 _64913_ (.D(_05935_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [447]),
    .QN(_31467_));
 DFF_X1 _64914_ (.D(_05936_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [448]),
    .QN(_31468_));
 DFF_X1 _64915_ (.D(_05937_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [449]),
    .QN(_31469_));
 DFF_X1 _64916_ (.D(_05939_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [450]),
    .QN(_31470_));
 DFF_X1 _64917_ (.D(_05940_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [451]),
    .QN(_31471_));
 DFF_X1 _64918_ (.D(_05941_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [452]),
    .QN(_31472_));
 DFF_X1 _64919_ (.D(_05942_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [453]),
    .QN(_31473_));
 DFF_X1 _64920_ (.D(_05943_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [454]),
    .QN(_31474_));
 DFF_X1 _64921_ (.D(_05944_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [455]),
    .QN(_31475_));
 DFF_X1 _64922_ (.D(_05945_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [456]),
    .QN(_31476_));
 DFF_X1 _64923_ (.D(_05946_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [457]),
    .QN(_31477_));
 DFF_X1 _64924_ (.D(_05947_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [458]),
    .QN(_31478_));
 DFF_X1 _64925_ (.D(_05948_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [459]),
    .QN(_31479_));
 DFF_X1 _64926_ (.D(_05950_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [460]),
    .QN(_31480_));
 DFF_X1 _64927_ (.D(_05951_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [461]),
    .QN(_31481_));
 DFF_X1 _64928_ (.D(_05952_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [462]),
    .QN(_31482_));
 DFF_X1 _64929_ (.D(_05953_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [463]),
    .QN(_31483_));
 DFF_X1 _64930_ (.D(_05954_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [464]),
    .QN(_31484_));
 DFF_X1 _64931_ (.D(_05955_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [465]),
    .QN(_31485_));
 DFF_X1 _64932_ (.D(_05956_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [466]),
    .QN(_31486_));
 DFF_X1 _64933_ (.D(_05957_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [467]),
    .QN(_31487_));
 DFF_X1 _64934_ (.D(_05958_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [468]),
    .QN(_31488_));
 DFF_X1 _64935_ (.D(_05959_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [469]),
    .QN(_31489_));
 DFF_X1 _64936_ (.D(_05961_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [470]),
    .QN(_31490_));
 DFF_X1 _64937_ (.D(_05962_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [471]),
    .QN(_31491_));
 DFF_X1 _64938_ (.D(_05963_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [472]),
    .QN(_31492_));
 DFF_X1 _64939_ (.D(_05964_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [473]),
    .QN(_31493_));
 DFF_X1 _64940_ (.D(_05965_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [474]),
    .QN(_31494_));
 DFF_X1 _64941_ (.D(_05966_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [475]),
    .QN(_31495_));
 DFF_X1 _64942_ (.D(_05967_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [476]),
    .QN(_31496_));
 DFF_X1 _64943_ (.D(_05968_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [477]),
    .QN(_31497_));
 DFF_X1 _64944_ (.D(_05969_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [478]),
    .QN(_31498_));
 DFF_X1 _64945_ (.D(_05970_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [479]),
    .QN(_31499_));
 DFF_X1 _64946_ (.D(_05972_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [480]),
    .QN(_31500_));
 DFF_X1 _64947_ (.D(_05973_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [481]),
    .QN(_31501_));
 DFF_X1 _64948_ (.D(_05974_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [482]),
    .QN(_31502_));
 DFF_X1 _64949_ (.D(_05975_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [483]),
    .QN(_31503_));
 DFF_X1 _64950_ (.D(_05976_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [484]),
    .QN(_31504_));
 DFF_X1 _64951_ (.D(_05977_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [485]),
    .QN(_31505_));
 DFF_X1 _64952_ (.D(_05978_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [486]),
    .QN(_31506_));
 DFF_X1 _64953_ (.D(_05979_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [487]),
    .QN(_31507_));
 DFF_X1 _64954_ (.D(_05980_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [488]),
    .QN(_31508_));
 DFF_X1 _64955_ (.D(_05981_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [489]),
    .QN(_31509_));
 DFF_X1 _64956_ (.D(_05983_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [490]),
    .QN(_31510_));
 DFF_X1 _64957_ (.D(_05984_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [491]),
    .QN(_31511_));
 DFF_X1 _64958_ (.D(_05985_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [492]),
    .QN(_31512_));
 DFF_X1 _64959_ (.D(_05986_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [493]),
    .QN(_31513_));
 DFF_X1 _64960_ (.D(_05987_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [494]),
    .QN(_31514_));
 DFF_X1 _64961_ (.D(_05988_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [495]),
    .QN(_31515_));
 DFF_X1 _64962_ (.D(_05989_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [496]),
    .QN(_31516_));
 DFF_X1 _64963_ (.D(_05990_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [497]),
    .QN(_31517_));
 DFF_X1 _64964_ (.D(_05991_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [498]),
    .QN(_31518_));
 DFF_X1 _64965_ (.D(_05992_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [499]),
    .QN(_31519_));
 DFF_X1 _64966_ (.D(_05995_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [500]),
    .QN(_31520_));
 DFF_X1 _64967_ (.D(_05996_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [501]),
    .QN(_31521_));
 DFF_X1 _64968_ (.D(_05997_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [502]),
    .QN(_31522_));
 DFF_X1 _64969_ (.D(_05998_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [503]),
    .QN(_31523_));
 DFF_X1 _64970_ (.D(_05999_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [504]),
    .QN(_31524_));
 DFF_X1 _64971_ (.D(_06000_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [505]),
    .QN(_31525_));
 DFF_X1 _64972_ (.D(_06001_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [506]),
    .QN(_31526_));
 DFF_X1 _64973_ (.D(_06002_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [507]),
    .QN(_31527_));
 DFF_X1 _64974_ (.D(_06003_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [508]),
    .QN(_31528_));
 DFF_X1 _64975_ (.D(_06004_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [509]),
    .QN(_31529_));
 DFF_X1 _64976_ (.D(_06006_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [510]),
    .QN(_31530_));
 DFF_X1 _64977_ (.D(_06007_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [511]),
    .QN(_31531_));
 DFF_X1 _64978_ (.D(_06008_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [512]),
    .QN(_31532_));
 DFF_X1 _64979_ (.D(_06009_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [513]),
    .QN(_31533_));
 DFF_X1 _64980_ (.D(_06010_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [514]),
    .QN(_31534_));
 DFF_X1 _64981_ (.D(_06011_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [515]),
    .QN(_31535_));
 DFF_X1 _64982_ (.D(_06012_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [516]),
    .QN(_31536_));
 DFF_X1 _64983_ (.D(_06013_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [517]),
    .QN(_31537_));
 DFF_X1 _64984_ (.D(_06014_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [518]),
    .QN(_31538_));
 DFF_X1 _64985_ (.D(_06015_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [519]),
    .QN(_31539_));
 DFF_X1 _64986_ (.D(_06017_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [520]),
    .QN(_31540_));
 DFF_X1 _64987_ (.D(_06018_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [521]),
    .QN(_31541_));
 DFF_X1 _64988_ (.D(_06019_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [522]),
    .QN(_31542_));
 DFF_X1 _64989_ (.D(_06020_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [524]),
    .QN(_31543_));
 DFF_X1 _64990_ (.D(_06021_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [525]),
    .QN(_31544_));
 DFF_X1 _64991_ (.D(_06022_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [526]),
    .QN(_31545_));
 DFF_X1 _64992_ (.D(_06023_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [527]),
    .QN(_31546_));
 DFF_X1 _64993_ (.D(_06024_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [528]),
    .QN(_31547_));
 DFF_X1 _64994_ (.D(_06025_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [529]),
    .QN(_31548_));
 DFF_X1 _64995_ (.D(_06027_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [530]),
    .QN(_31549_));
 DFF_X1 _64996_ (.D(_06028_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [531]),
    .QN(_31550_));
 DFF_X1 _64997_ (.D(_06029_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [532]),
    .QN(_31551_));
 DFF_X1 _64998_ (.D(_06030_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [533]),
    .QN(_31552_));
 DFF_X1 _64999_ (.D(_06031_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [534]),
    .QN(_31553_));
 DFF_X1 _65000_ (.D(_06032_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [535]),
    .QN(_31554_));
 DFF_X1 _65001_ (.D(_06033_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [536]),
    .QN(_31555_));
 DFF_X1 _65002_ (.D(_06034_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [537]),
    .QN(_31556_));
 DFF_X1 _65003_ (.D(_06035_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [538]),
    .QN(_31557_));
 DFF_X1 _65004_ (.D(_06036_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [539]),
    .QN(_31558_));
 DFF_X1 _65005_ (.D(_06038_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [540]),
    .QN(_31559_));
 DFF_X1 _65006_ (.D(_06039_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [541]),
    .QN(_31560_));
 DFF_X1 _65007_ (.D(_06040_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [542]),
    .QN(_31561_));
 DFF_X1 _65008_ (.D(_06041_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [543]),
    .QN(_31562_));
 DFF_X1 _65009_ (.D(_06042_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [544]),
    .QN(_31563_));
 DFF_X1 _65010_ (.D(_06043_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [545]),
    .QN(_31564_));
 DFF_X1 _65011_ (.D(_06044_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [546]),
    .QN(_31565_));
 DFF_X1 _65012_ (.D(_06045_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [547]),
    .QN(_31566_));
 DFF_X1 _65013_ (.D(_06046_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [548]),
    .QN(_31567_));
 DFF_X1 _65014_ (.D(_06047_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [549]),
    .QN(_31568_));
 DFF_X1 _65015_ (.D(_06049_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [550]),
    .QN(_31569_));
 DFF_X1 _65016_ (.D(_06050_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [551]),
    .QN(_31570_));
 DFF_X1 _65017_ (.D(_06051_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [552]),
    .QN(_31571_));
 DFF_X1 _65018_ (.D(_06052_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [553]),
    .QN(_31572_));
 DFF_X1 _65019_ (.D(_06053_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [554]),
    .QN(_31573_));
 DFF_X1 _65020_ (.D(_06054_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [555]),
    .QN(_31574_));
 DFF_X1 _65021_ (.D(_06055_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [556]),
    .QN(_31575_));
 DFF_X1 _65022_ (.D(_06056_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [557]),
    .QN(_31576_));
 DFF_X1 _65023_ (.D(_06057_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [558]),
    .QN(_31577_));
 DFF_X1 _65024_ (.D(_06058_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [559]),
    .QN(_31578_));
 DFF_X1 _65025_ (.D(_06060_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [560]),
    .QN(_31579_));
 DFF_X1 _65026_ (.D(_06061_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [561]),
    .QN(_31580_));
 DFF_X1 _65027_ (.D(_06062_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [562]),
    .QN(_31581_));
 DFF_X1 _65028_ (.D(_06063_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [563]),
    .QN(_31582_));
 DFF_X1 _65029_ (.D(_06064_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [564]),
    .QN(_31583_));
 DFF_X1 _65030_ (.D(_06065_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [565]),
    .QN(_31584_));
 DFF_X1 _65031_ (.D(_06066_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [566]),
    .QN(_31585_));
 DFF_X1 _65032_ (.D(_06067_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [567]),
    .QN(_31586_));
 DFF_X1 _65033_ (.D(_06068_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [568]),
    .QN(_31587_));
 DFF_X1 _65034_ (.D(_06069_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [569]),
    .QN(_31588_));
 DFF_X1 _65035_ (.D(_06071_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [570]),
    .QN(_31589_));
 DFF_X1 _65036_ (.D(_06072_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [571]),
    .QN(_31590_));
 DFF_X1 _65037_ (.D(_06073_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [572]),
    .QN(_31591_));
 DFF_X1 _65038_ (.D(_06074_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [573]),
    .QN(_31592_));
 DFF_X1 _65039_ (.D(_06075_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [574]),
    .QN(_31593_));
 DFF_X1 _65040_ (.D(_06076_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [575]),
    .QN(_31594_));
 DFF_X1 _65041_ (.D(_06077_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [576]),
    .QN(_31595_));
 DFF_X1 _65042_ (.D(_06078_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [577]),
    .QN(_31596_));
 DFF_X1 _65043_ (.D(_06079_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [578]),
    .QN(_31597_));
 DFF_X1 _65044_ (.D(_06080_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [579]),
    .QN(_31598_));
 DFF_X1 _65045_ (.D(_06082_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [580]),
    .QN(_31599_));
 DFF_X1 _65046_ (.D(_06083_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [581]),
    .QN(_31600_));
 DFF_X1 _65047_ (.D(_06084_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [582]),
    .QN(_31601_));
 DFF_X1 _65048_ (.D(_06085_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [583]),
    .QN(_31602_));
 DFF_X1 _65049_ (.D(_06086_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [584]),
    .QN(_31603_));
 DFF_X1 _65050_ (.D(_06087_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [585]),
    .QN(_31604_));
 DFF_X1 _65051_ (.D(_06088_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [586]),
    .QN(_31605_));
 DFF_X1 _65052_ (.D(_06089_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [587]),
    .QN(_31606_));
 DFF_X1 _65053_ (.D(_06090_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [588]),
    .QN(_31607_));
 DFF_X1 _65054_ (.D(_06091_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [589]),
    .QN(_31608_));
 DFF_X1 _65055_ (.D(_06093_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [590]),
    .QN(_31609_));
 DFF_X1 _65056_ (.D(_06094_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [591]),
    .QN(_31610_));
 DFF_X1 _65057_ (.D(_06095_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [592]),
    .QN(_31611_));
 DFF_X1 _65058_ (.D(_06096_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [593]),
    .QN(_31612_));
 DFF_X1 _65059_ (.D(_06097_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [594]),
    .QN(_31613_));
 DFF_X1 _65060_ (.D(_06098_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [595]),
    .QN(_31614_));
 DFF_X1 _65061_ (.D(_06099_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [596]),
    .QN(_31615_));
 DFF_X1 _65062_ (.D(_06100_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [597]),
    .QN(_31616_));
 DFF_X1 _65063_ (.D(_06101_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [598]),
    .QN(_31617_));
 DFF_X1 _65064_ (.D(_06102_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [599]),
    .QN(_31618_));
 DFF_X1 _65065_ (.D(_06104_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [600]),
    .QN(_31619_));
 DFF_X1 _65066_ (.D(_06105_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [601]),
    .QN(_31620_));
 DFF_X1 _65067_ (.D(_06106_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [602]),
    .QN(_31621_));
 DFF_X1 _65068_ (.D(_06107_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [603]),
    .QN(_31622_));
 DFF_X1 _65069_ (.D(_06108_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [604]),
    .QN(_31623_));
 DFF_X1 _65070_ (.D(_06109_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [605]),
    .QN(_31624_));
 DFF_X1 _65071_ (.D(_06110_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [606]),
    .QN(_31625_));
 DFF_X1 _65072_ (.D(_06111_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [607]),
    .QN(_31626_));
 DFF_X1 _65073_ (.D(_06112_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [608]),
    .QN(_31627_));
 DFF_X1 _65074_ (.D(_06113_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [609]),
    .QN(_31628_));
 DFF_X1 _65075_ (.D(_06115_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [610]),
    .QN(_31629_));
 DFF_X1 _65076_ (.D(_06116_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [611]),
    .QN(_31630_));
 DFF_X1 _65077_ (.D(_06117_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [612]),
    .QN(_31631_));
 DFF_X1 _65078_ (.D(_06118_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [613]),
    .QN(_31632_));
 DFF_X1 _65079_ (.D(_06119_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [614]),
    .QN(_31633_));
 DFF_X1 _65080_ (.D(_06120_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [615]),
    .QN(_31634_));
 DFF_X1 _65081_ (.D(_06121_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [616]),
    .QN(_31635_));
 DFF_X1 _65082_ (.D(_06122_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [617]),
    .QN(_31636_));
 DFF_X1 _65083_ (.D(_06123_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [618]),
    .QN(_31637_));
 DFF_X1 _65084_ (.D(_06124_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [619]),
    .QN(_31638_));
 DFF_X1 _65085_ (.D(_06126_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [620]),
    .QN(_31639_));
 DFF_X1 _65086_ (.D(_06127_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [621]),
    .QN(_31640_));
 DFF_X1 _65087_ (.D(_06128_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [622]),
    .QN(_31641_));
 DFF_X1 _65088_ (.D(_06129_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [623]),
    .QN(_31642_));
 DFF_X1 _65089_ (.D(_06130_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [624]),
    .QN(_31643_));
 DFF_X1 _65090_ (.D(_06131_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [625]),
    .QN(_31644_));
 DFF_X1 _65091_ (.D(_06132_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [626]),
    .QN(_31645_));
 DFF_X1 _65092_ (.D(_06133_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [627]),
    .QN(_31646_));
 DFF_X1 _65093_ (.D(_06134_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [628]),
    .QN(_31647_));
 DFF_X1 _65094_ (.D(_06135_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [629]),
    .QN(_31648_));
 DFF_X1 _65095_ (.D(_06137_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [630]),
    .QN(_31649_));
 DFF_X1 _65096_ (.D(_06138_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [631]),
    .QN(_31650_));
 DFF_X1 _65097_ (.D(_06139_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [632]),
    .QN(_31651_));
 DFF_X1 _65098_ (.D(_06140_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [633]),
    .QN(_31652_));
 DFF_X1 _65099_ (.D(_06141_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [634]),
    .QN(_31653_));
 DFF_X1 _65100_ (.D(_06142_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [635]),
    .QN(_31654_));
 DFF_X1 _65101_ (.D(_06143_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [636]),
    .QN(_31655_));
 DFF_X1 _65102_ (.D(_06144_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [637]),
    .QN(_31656_));
 DFF_X1 _65103_ (.D(_06145_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [638]),
    .QN(_31657_));
 DFF_X1 _65104_ (.D(_06146_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [639]),
    .QN(_31658_));
 DFF_X1 _65105_ (.D(_06148_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [640]),
    .QN(_31659_));
 DFF_X1 _65106_ (.D(_06149_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [641]),
    .QN(_31660_));
 DFF_X1 _65107_ (.D(_06150_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [642]),
    .QN(_31661_));
 DFF_X1 _65108_ (.D(_06151_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [643]),
    .QN(_31662_));
 DFF_X1 _65109_ (.D(_06152_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [644]),
    .QN(_31663_));
 DFF_X1 _65110_ (.D(_06153_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [645]),
    .QN(_31664_));
 DFF_X1 _65111_ (.D(_06154_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [646]),
    .QN(_31665_));
 DFF_X1 _65112_ (.D(_06155_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [647]),
    .QN(_31666_));
 DFF_X1 _65113_ (.D(_06156_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [648]),
    .QN(_31667_));
 DFF_X1 _65114_ (.D(_06157_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [649]),
    .QN(_31668_));
 DFF_X1 _65115_ (.D(_06159_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [650]),
    .QN(_31669_));
 DFF_X1 _65116_ (.D(_06160_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [651]),
    .QN(_31670_));
 DFF_X1 _65117_ (.D(_06161_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [652]),
    .QN(_31671_));
 DFF_X1 _65118_ (.D(_06162_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [653]),
    .QN(_31672_));
 DFF_X1 _65119_ (.D(_06163_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [654]),
    .QN(_31673_));
 DFF_X1 _65120_ (.D(_06164_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [655]),
    .QN(_31674_));
 DFF_X1 _65121_ (.D(_06165_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [656]),
    .QN(_31675_));
 DFF_X1 _65122_ (.D(_06166_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [657]),
    .QN(_31676_));
 DFF_X1 _65123_ (.D(_06167_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [658]),
    .QN(_31677_));
 DFF_X1 _65124_ (.D(_06168_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [659]),
    .QN(_31678_));
 DFF_X1 _65125_ (.D(_06170_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [660]),
    .QN(_31679_));
 DFF_X1 _65126_ (.D(_06171_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [661]),
    .QN(_31680_));
 DFF_X1 _65127_ (.D(_06172_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [662]),
    .QN(_31681_));
 DFF_X1 _65128_ (.D(_06173_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [663]),
    .QN(_31682_));
 DFF_X1 _65129_ (.D(_06174_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [664]),
    .QN(_31683_));
 DFF_X1 _65130_ (.D(_06175_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [665]),
    .QN(_31684_));
 DFF_X1 _65131_ (.D(_06176_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [666]),
    .QN(_31685_));
 DFF_X1 _65132_ (.D(_06177_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [667]),
    .QN(_31686_));
 DFF_X1 _65133_ (.D(_06178_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [668]),
    .QN(_31687_));
 DFF_X1 _65134_ (.D(_06179_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [669]),
    .QN(_31688_));
 DFF_X1 _65135_ (.D(_06181_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [670]),
    .QN(_31689_));
 DFF_X1 _65136_ (.D(_06182_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [671]),
    .QN(_31690_));
 DFF_X1 _65137_ (.D(_06183_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [672]),
    .QN(_31691_));
 DFF_X1 _65138_ (.D(_06184_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [673]),
    .QN(_31692_));
 DFF_X1 _65139_ (.D(_06185_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [674]),
    .QN(_31693_));
 DFF_X1 _65140_ (.D(_06186_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [675]),
    .QN(_31694_));
 DFF_X1 _65141_ (.D(_06187_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [676]),
    .QN(_31695_));
 DFF_X1 _65142_ (.D(_06188_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [677]),
    .QN(_31696_));
 DFF_X1 _65143_ (.D(_06189_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [678]),
    .QN(_31697_));
 DFF_X1 _65144_ (.D(_06190_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [679]),
    .QN(_31698_));
 DFF_X1 _65145_ (.D(_06192_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [680]),
    .QN(_31699_));
 DFF_X1 _65146_ (.D(_06193_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [681]),
    .QN(_31700_));
 DFF_X1 _65147_ (.D(_06194_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [682]),
    .QN(_31701_));
 DFF_X1 _65148_ (.D(_06195_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [683]),
    .QN(_31702_));
 DFF_X1 _65149_ (.D(_06196_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [684]),
    .QN(_31703_));
 DFF_X1 _65150_ (.D(_06197_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [685]),
    .QN(_31704_));
 DFF_X1 _65151_ (.D(_06198_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [686]),
    .QN(_31705_));
 DFF_X1 _65152_ (.D(_06199_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [687]),
    .QN(_31706_));
 DFF_X1 _65153_ (.D(_06200_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [688]),
    .QN(_31707_));
 DFF_X1 _65154_ (.D(_06201_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [689]),
    .QN(_31708_));
 DFF_X1 _65155_ (.D(_06203_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [690]),
    .QN(_31709_));
 DFF_X1 _65156_ (.D(_06204_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [691]),
    .QN(_31710_));
 DFF_X1 _65157_ (.D(_06205_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [692]),
    .QN(_31711_));
 DFF_X1 _65158_ (.D(_06206_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [693]),
    .QN(_31712_));
 DFF_X1 _65159_ (.D(_06207_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [694]),
    .QN(_31713_));
 DFF_X1 _65160_ (.D(_06208_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [695]),
    .QN(_31714_));
 DFF_X1 _65161_ (.D(_06209_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [696]),
    .QN(_31715_));
 DFF_X1 _65162_ (.D(_06210_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [697]),
    .QN(_31716_));
 DFF_X1 _65163_ (.D(_06211_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [698]),
    .QN(_31717_));
 DFF_X1 _65164_ (.D(_06212_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [699]),
    .QN(_31718_));
 DFF_X1 _65165_ (.D(_06215_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [700]),
    .QN(_31719_));
 DFF_X1 _65166_ (.D(_06216_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [701]),
    .QN(_31720_));
 DFF_X1 _65167_ (.D(_06217_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [702]),
    .QN(_31721_));
 DFF_X1 _65168_ (.D(_06218_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [703]),
    .QN(_31722_));
 DFF_X1 _65169_ (.D(_06219_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [704]),
    .QN(_31723_));
 DFF_X1 _65170_ (.D(_06220_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [705]),
    .QN(_31724_));
 DFF_X1 _65171_ (.D(_06221_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [706]),
    .QN(_31725_));
 DFF_X1 _65172_ (.D(_06222_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [707]),
    .QN(_31726_));
 DFF_X1 _65173_ (.D(_06223_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [708]),
    .QN(_31727_));
 DFF_X1 _65174_ (.D(_06224_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [709]),
    .QN(_31728_));
 DFF_X1 _65175_ (.D(_06226_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [710]),
    .QN(_31729_));
 DFF_X1 _65176_ (.D(_06227_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [711]),
    .QN(_31730_));
 DFF_X1 _65177_ (.D(_06228_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [712]),
    .QN(_31731_));
 DFF_X1 _65178_ (.D(_06229_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [713]),
    .QN(_31732_));
 DFF_X1 _65179_ (.D(_06230_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [714]),
    .QN(_31733_));
 DFF_X1 _65180_ (.D(_06231_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [715]),
    .QN(_31734_));
 DFF_X1 _65181_ (.D(_06232_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [716]),
    .QN(_31735_));
 DFF_X1 _65182_ (.D(_06233_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [717]),
    .QN(_31736_));
 DFF_X1 _65183_ (.D(_06234_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [718]),
    .QN(_31737_));
 DFF_X1 _65184_ (.D(_06235_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [719]),
    .QN(_31738_));
 DFF_X1 _65185_ (.D(_06237_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [720]),
    .QN(_31739_));
 DFF_X1 _65186_ (.D(_06238_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [721]),
    .QN(_31740_));
 DFF_X1 _65187_ (.D(_06239_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [722]),
    .QN(_31741_));
 DFF_X1 _65188_ (.D(_06240_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [723]),
    .QN(_31742_));
 DFF_X1 _65189_ (.D(_06241_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [724]),
    .QN(_31743_));
 DFF_X1 _65190_ (.D(_06242_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [725]),
    .QN(_31744_));
 DFF_X1 _65191_ (.D(_06243_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [726]),
    .QN(_31745_));
 DFF_X1 _65192_ (.D(_06244_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [727]),
    .QN(_31746_));
 DFF_X1 _65193_ (.D(_06245_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [728]),
    .QN(_31747_));
 DFF_X1 _65194_ (.D(_06246_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [729]),
    .QN(_31748_));
 DFF_X1 _65195_ (.D(_06248_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [730]),
    .QN(_31749_));
 DFF_X1 _65196_ (.D(_06249_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [731]),
    .QN(_31750_));
 DFF_X1 _65197_ (.D(_06250_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [732]),
    .QN(_31751_));
 DFF_X1 _65198_ (.D(_06251_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [733]),
    .QN(_31752_));
 DFF_X1 _65199_ (.D(_06252_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [734]),
    .QN(_31753_));
 DFF_X1 _65200_ (.D(_06253_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [735]),
    .QN(_31754_));
 DFF_X1 _65201_ (.D(_06254_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [736]),
    .QN(_31755_));
 DFF_X1 _65202_ (.D(_06255_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [737]),
    .QN(_31756_));
 DFF_X1 _65203_ (.D(_06256_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [738]),
    .QN(_31757_));
 DFF_X1 _65204_ (.D(_06257_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [739]),
    .QN(_31758_));
 DFF_X1 _65205_ (.D(_06259_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [740]),
    .QN(_31759_));
 DFF_X1 _65206_ (.D(_06260_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [741]),
    .QN(_31760_));
 DFF_X1 _65207_ (.D(_06261_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [742]),
    .QN(_31761_));
 DFF_X1 _65208_ (.D(_06262_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [743]),
    .QN(_31762_));
 DFF_X1 _65209_ (.D(_06263_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [744]),
    .QN(_31763_));
 DFF_X1 _65210_ (.D(_06264_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [745]),
    .QN(_31764_));
 DFF_X1 _65211_ (.D(_06265_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [746]),
    .QN(_31765_));
 DFF_X1 _65212_ (.D(_06266_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [747]),
    .QN(_31766_));
 DFF_X1 _65213_ (.D(_06267_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [748]),
    .QN(_31767_));
 DFF_X1 _65214_ (.D(_06268_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [749]),
    .QN(_31768_));
 DFF_X1 _65215_ (.D(_06270_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [750]),
    .QN(_31769_));
 DFF_X1 _65216_ (.D(_06271_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [751]),
    .QN(_31770_));
 DFF_X1 _65217_ (.D(_06272_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [752]),
    .QN(_31771_));
 DFF_X1 _65218_ (.D(_06273_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [753]),
    .QN(_31772_));
 DFF_X1 _65219_ (.D(_06274_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [754]),
    .QN(_31773_));
 DFF_X1 _65220_ (.D(_06275_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [755]),
    .QN(_31774_));
 DFF_X1 _65221_ (.D(_06276_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [756]),
    .QN(_31775_));
 DFF_X1 _65222_ (.D(_06277_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [757]),
    .QN(_31776_));
 DFF_X1 _65223_ (.D(_06278_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [758]),
    .QN(_31777_));
 DFF_X1 _65224_ (.D(_06279_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [759]),
    .QN(_31778_));
 DFF_X1 _65225_ (.D(_06281_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [760]),
    .QN(_31779_));
 DFF_X1 _65226_ (.D(_06282_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [761]),
    .QN(_31780_));
 DFF_X1 _65227_ (.D(_06283_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [762]),
    .QN(_31781_));
 DFF_X1 _65228_ (.D(_06284_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [763]),
    .QN(_31782_));
 DFF_X1 _65229_ (.D(_06285_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [764]),
    .QN(_31783_));
 DFF_X1 _65230_ (.D(_06286_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [765]),
    .QN(_31784_));
 DFF_X1 _65231_ (.D(_06287_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [766]),
    .QN(_31785_));
 DFF_X1 _65232_ (.D(_06288_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [767]),
    .QN(_31786_));
 DFF_X1 _65233_ (.D(_06289_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [768]),
    .QN(_31787_));
 DFF_X1 _65234_ (.D(_06290_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [769]),
    .QN(_31788_));
 DFF_X1 _65235_ (.D(_06292_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [770]),
    .QN(_31789_));
 DFF_X1 _65236_ (.D(_06293_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [771]),
    .QN(_31790_));
 DFF_X1 _65237_ (.D(_06294_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [772]),
    .QN(_31791_));
 DFF_X1 _65238_ (.D(_06295_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [773]),
    .QN(_31792_));
 DFF_X1 _65239_ (.D(_06296_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [774]),
    .QN(_31793_));
 DFF_X1 _65240_ (.D(_06297_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [775]),
    .QN(_31794_));
 DFF_X1 _65241_ (.D(_06298_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [776]),
    .QN(_31795_));
 DFF_X1 _65242_ (.D(_06299_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [777]),
    .QN(_31796_));
 DFF_X1 _65243_ (.D(_06300_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [778]),
    .QN(_31797_));
 DFF_X1 _65244_ (.D(_06301_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [779]),
    .QN(_31798_));
 DFF_X1 _65245_ (.D(_06303_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [780]),
    .QN(_31799_));
 DFF_X1 _65246_ (.D(_06304_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [781]),
    .QN(_31800_));
 DFF_X1 _65247_ (.D(_06305_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [782]),
    .QN(_31801_));
 DFF_X1 _65248_ (.D(_06306_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [783]),
    .QN(_31802_));
 DFF_X1 _65249_ (.D(_06307_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [784]),
    .QN(_31803_));
 DFF_X1 _65250_ (.D(_06308_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [785]),
    .QN(_31804_));
 DFF_X1 _65251_ (.D(_06309_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [786]),
    .QN(_31805_));
 DFF_X1 _65252_ (.D(_06310_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [787]),
    .QN(_31806_));
 DFF_X1 _65253_ (.D(_06311_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [788]),
    .QN(_31807_));
 DFF_X1 _65254_ (.D(_06312_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [789]),
    .QN(_31808_));
 DFF_X1 _65255_ (.D(_06314_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [790]),
    .QN(_31809_));
 DFF_X1 _65256_ (.D(_06315_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [791]),
    .QN(_31810_));
 DFF_X1 _65257_ (.D(_06316_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [792]),
    .QN(_31811_));
 DFF_X1 _65258_ (.D(_06317_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [793]),
    .QN(_31812_));
 DFF_X1 _65259_ (.D(_06318_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [794]),
    .QN(_31813_));
 DFF_X1 _65260_ (.D(_06319_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [795]),
    .QN(_31814_));
 DFF_X1 _65261_ (.D(_06320_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [796]),
    .QN(_31815_));
 DFF_X1 _65262_ (.D(_06321_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [797]),
    .QN(_31816_));
 DFF_X1 _65263_ (.D(_06322_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [798]),
    .QN(_31817_));
 DFF_X1 _65264_ (.D(_06323_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [799]),
    .QN(_31818_));
 DFF_X1 _65265_ (.D(_06326_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [800]),
    .QN(_31819_));
 DFF_X1 _65266_ (.D(_06327_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [801]),
    .QN(_31820_));
 DFF_X1 _65267_ (.D(_06328_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [802]),
    .QN(_31821_));
 DFF_X1 _65268_ (.D(_06329_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [803]),
    .QN(_31822_));
 DFF_X1 _65269_ (.D(_06330_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [804]),
    .QN(_31823_));
 DFF_X1 _65270_ (.D(_06331_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [805]),
    .QN(_31824_));
 DFF_X1 _65271_ (.D(_06332_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [806]),
    .QN(_31825_));
 DFF_X1 _65272_ (.D(_06333_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [807]),
    .QN(_31826_));
 DFF_X1 _65273_ (.D(_06334_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [808]),
    .QN(_31827_));
 DFF_X1 _65274_ (.D(_06335_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [809]),
    .QN(_31828_));
 DFF_X1 _65275_ (.D(_06337_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [810]),
    .QN(_31829_));
 DFF_X1 _65276_ (.D(_06338_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [811]),
    .QN(_31830_));
 DFF_X1 _65277_ (.D(_06339_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [812]),
    .QN(_31831_));
 DFF_X1 _65278_ (.D(_06340_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [813]),
    .QN(_31832_));
 DFF_X1 _65279_ (.D(_06341_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [814]),
    .QN(_31833_));
 DFF_X1 _65280_ (.D(_06342_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [815]),
    .QN(_31834_));
 DFF_X1 _65281_ (.D(_06343_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [816]),
    .QN(_31835_));
 DFF_X1 _65282_ (.D(_06344_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [817]),
    .QN(_31836_));
 DFF_X1 _65283_ (.D(_06345_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [818]),
    .QN(_31837_));
 DFF_X1 _65284_ (.D(_06346_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [819]),
    .QN(_31838_));
 DFF_X1 _65285_ (.D(_06348_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [820]),
    .QN(_31839_));
 DFF_X1 _65286_ (.D(_06349_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [821]),
    .QN(_31840_));
 DFF_X1 _65287_ (.D(_06350_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [822]),
    .QN(_31841_));
 DFF_X1 _65288_ (.D(_06351_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [823]),
    .QN(_31842_));
 DFF_X1 _65289_ (.D(_06352_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [824]),
    .QN(_31843_));
 DFF_X1 _65290_ (.D(_06353_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [825]),
    .QN(_31844_));
 DFF_X1 _65291_ (.D(_06354_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [826]),
    .QN(_31845_));
 DFF_X1 _65292_ (.D(_06355_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [827]),
    .QN(_31846_));
 DFF_X1 _65293_ (.D(_06356_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [828]),
    .QN(_31847_));
 DFF_X1 _65294_ (.D(_06357_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [829]),
    .QN(_31848_));
 DFF_X1 _65295_ (.D(_06359_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [830]),
    .QN(_31849_));
 DFF_X1 _65296_ (.D(_06360_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [831]),
    .QN(_31850_));
 DFF_X1 _65297_ (.D(_06361_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [832]),
    .QN(_31851_));
 DFF_X1 _65298_ (.D(_06362_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [833]),
    .QN(_31852_));
 DFF_X1 _65299_ (.D(_06363_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [834]),
    .QN(_31853_));
 DFF_X1 _65300_ (.D(_06364_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [835]),
    .QN(_31854_));
 DFF_X1 _65301_ (.D(_06365_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [836]),
    .QN(_31855_));
 DFF_X1 _65302_ (.D(_06366_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [837]),
    .QN(_31856_));
 DFF_X1 _65303_ (.D(_06367_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [838]),
    .QN(_31857_));
 DFF_X1 _65304_ (.D(_06368_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [839]),
    .QN(_31858_));
 DFF_X1 _65305_ (.D(_06370_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [840]),
    .QN(_31859_));
 DFF_X1 _65306_ (.D(_06371_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [841]),
    .QN(_31860_));
 DFF_X1 _65307_ (.D(_06372_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [842]),
    .QN(_31861_));
 DFF_X1 _65308_ (.D(_06373_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [843]),
    .QN(_31862_));
 DFF_X1 _65309_ (.D(_06374_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [844]),
    .QN(_31863_));
 DFF_X1 _65310_ (.D(_06375_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [845]),
    .QN(_31864_));
 DFF_X1 _65311_ (.D(_06376_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [846]),
    .QN(_31865_));
 DFF_X1 _65312_ (.D(_06377_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [847]),
    .QN(_31866_));
 DFF_X1 _65313_ (.D(_06378_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [848]),
    .QN(_31867_));
 DFF_X1 _65314_ (.D(_06379_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [849]),
    .QN(_31868_));
 DFF_X1 _65315_ (.D(_06381_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [850]),
    .QN(_31869_));
 DFF_X1 _65316_ (.D(_06382_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [851]),
    .QN(_31870_));
 DFF_X1 _65317_ (.D(_06383_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [852]),
    .QN(_31871_));
 DFF_X1 _65318_ (.D(_06384_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [853]),
    .QN(_31872_));
 DFF_X1 _65319_ (.D(_06385_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [854]),
    .QN(_31873_));
 DFF_X1 _65320_ (.D(_06386_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [855]),
    .QN(_31874_));
 DFF_X1 _65321_ (.D(_06387_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [856]),
    .QN(_31875_));
 DFF_X1 _65322_ (.D(_06388_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [857]),
    .QN(_31876_));
 DFF_X1 _65323_ (.D(_06389_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [858]),
    .QN(_31877_));
 DFF_X1 _65324_ (.D(_06390_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [859]),
    .QN(_31878_));
 DFF_X1 _65325_ (.D(_06392_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [860]),
    .QN(_31879_));
 DFF_X1 _65326_ (.D(_06393_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [861]),
    .QN(_31880_));
 DFF_X1 _65327_ (.D(_06394_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [862]),
    .QN(_31881_));
 DFF_X1 _65328_ (.D(_06395_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [863]),
    .QN(_31882_));
 DFF_X1 _65329_ (.D(_06396_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [864]),
    .QN(_31883_));
 DFF_X1 _65330_ (.D(_06397_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [865]),
    .QN(_31884_));
 DFF_X1 _65331_ (.D(_06398_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [866]),
    .QN(_31885_));
 DFF_X1 _65332_ (.D(_06399_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [867]),
    .QN(_31886_));
 DFF_X1 _65333_ (.D(_06400_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [868]),
    .QN(_31887_));
 DFF_X1 _65334_ (.D(_06401_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [869]),
    .QN(_31888_));
 DFF_X1 _65335_ (.D(_06403_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [870]),
    .QN(_31889_));
 DFF_X1 _65336_ (.D(_06404_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [871]),
    .QN(_31890_));
 DFF_X1 _65337_ (.D(_06405_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [872]),
    .QN(_31891_));
 DFF_X1 _65338_ (.D(_06406_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [873]),
    .QN(_31892_));
 DFF_X1 _65339_ (.D(_06407_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [874]),
    .QN(_31893_));
 DFF_X1 _65340_ (.D(_06408_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [875]),
    .QN(_31894_));
 DFF_X1 _65341_ (.D(_06409_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [876]),
    .QN(_31895_));
 DFF_X1 _65342_ (.D(_06410_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [877]),
    .QN(_31896_));
 DFF_X1 _65343_ (.D(_06411_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [878]),
    .QN(_31897_));
 DFF_X1 _65344_ (.D(_06412_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [879]),
    .QN(_31898_));
 DFF_X1 _65345_ (.D(_06414_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [880]),
    .QN(_31899_));
 DFF_X1 _65346_ (.D(_06415_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [881]),
    .QN(_31900_));
 DFF_X1 _65347_ (.D(_06416_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [882]),
    .QN(_31901_));
 DFF_X1 _65348_ (.D(_06417_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [883]),
    .QN(_31902_));
 DFF_X1 _65349_ (.D(_06418_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [884]),
    .QN(_31903_));
 DFF_X1 _65350_ (.D(_06419_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [885]),
    .QN(_31904_));
 DFF_X1 _65351_ (.D(_06420_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [886]),
    .QN(_31905_));
 DFF_X1 _65352_ (.D(_06421_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [887]),
    .QN(_31906_));
 DFF_X1 _65353_ (.D(_06422_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [888]),
    .QN(_31907_));
 DFF_X1 _65354_ (.D(_06423_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [889]),
    .QN(_31908_));
 DFF_X1 _65355_ (.D(_06425_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [890]),
    .QN(_31909_));
 DFF_X1 _65356_ (.D(_06426_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [891]),
    .QN(_31910_));
 DFF_X1 _65357_ (.D(_06427_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [892]),
    .QN(_31911_));
 DFF_X1 _65358_ (.D(_06428_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [893]),
    .QN(_31912_));
 DFF_X1 _65359_ (.D(_06429_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [894]),
    .QN(_31913_));
 DFF_X1 _65360_ (.D(_06430_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [895]),
    .QN(_31914_));
 DFF_X1 _65361_ (.D(_06431_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [896]),
    .QN(_31915_));
 DFF_X1 _65362_ (.D(_06432_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [897]),
    .QN(_31916_));
 DFF_X1 _65363_ (.D(_06433_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [898]),
    .QN(_31917_));
 DFF_X1 _65364_ (.D(_06434_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [899]),
    .QN(_31918_));
 DFF_X1 _65365_ (.D(_06437_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [900]),
    .QN(_31919_));
 DFF_X1 _65366_ (.D(_06438_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [901]),
    .QN(_31920_));
 DFF_X1 _65367_ (.D(_06439_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [902]),
    .QN(_31921_));
 DFF_X1 _65368_ (.D(_06440_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [903]),
    .QN(_31922_));
 DFF_X1 _65369_ (.D(_06441_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [904]),
    .QN(_31923_));
 DFF_X1 _65370_ (.D(_06442_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [905]),
    .QN(_31924_));
 DFF_X1 _65371_ (.D(_06443_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [906]),
    .QN(_31925_));
 DFF_X1 _65372_ (.D(_06444_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [907]),
    .QN(_31926_));
 DFF_X1 _65373_ (.D(_06445_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [908]),
    .QN(_31927_));
 DFF_X1 _65374_ (.D(_06446_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [909]),
    .QN(_31928_));
 DFF_X1 _65375_ (.D(_06448_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [910]),
    .QN(_31929_));
 DFF_X1 _65376_ (.D(_06449_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [911]),
    .QN(_31930_));
 DFF_X1 _65377_ (.D(_06450_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [912]),
    .QN(_31931_));
 DFF_X1 _65378_ (.D(_06451_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [913]),
    .QN(_31932_));
 DFF_X1 _65379_ (.D(_06452_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [914]),
    .QN(_31933_));
 DFF_X1 _65380_ (.D(_06453_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [915]),
    .QN(_31934_));
 DFF_X1 _65381_ (.D(_06454_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [916]),
    .QN(_31935_));
 DFF_X1 _65382_ (.D(_06455_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [917]),
    .QN(_31936_));
 DFF_X1 _65383_ (.D(_06456_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [918]),
    .QN(_31937_));
 DFF_X1 _65384_ (.D(_06457_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [919]),
    .QN(_31938_));
 DFF_X1 _65385_ (.D(_06459_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [920]),
    .QN(_31939_));
 DFF_X1 _65386_ (.D(_06460_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [921]),
    .QN(_31940_));
 DFF_X1 _65387_ (.D(_06461_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [922]),
    .QN(_31941_));
 DFF_X1 _65388_ (.D(_06462_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [923]),
    .QN(_31942_));
 DFF_X1 _65389_ (.D(_06463_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [924]),
    .QN(_31943_));
 DFF_X1 _65390_ (.D(_06464_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [925]),
    .QN(_31944_));
 DFF_X1 _65391_ (.D(_06465_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [926]),
    .QN(_31945_));
 DFF_X1 _65392_ (.D(_06466_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [927]),
    .QN(_31946_));
 DFF_X1 _65393_ (.D(_06467_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [928]),
    .QN(_31947_));
 DFF_X1 _65394_ (.D(_06468_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [929]),
    .QN(_31948_));
 DFF_X1 _65395_ (.D(_06470_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [930]),
    .QN(_31949_));
 DFF_X1 _65396_ (.D(_06471_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [931]),
    .QN(_31950_));
 DFF_X1 _65397_ (.D(_06472_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [932]),
    .QN(_31951_));
 DFF_X1 _65398_ (.D(_06473_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [933]),
    .QN(_31952_));
 DFF_X1 _65399_ (.D(_06474_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [934]),
    .QN(_31953_));
 DFF_X1 _65400_ (.D(_06475_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [935]),
    .QN(_31954_));
 DFF_X1 _65401_ (.D(_06476_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [936]),
    .QN(_31955_));
 DFF_X1 _65402_ (.D(_06477_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [937]),
    .QN(_31956_));
 DFF_X1 _65403_ (.D(_06478_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [938]),
    .QN(_31957_));
 DFF_X1 _65404_ (.D(_06479_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [939]),
    .QN(_31958_));
 DFF_X1 _65405_ (.D(_06481_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [940]),
    .QN(_31959_));
 DFF_X1 _65406_ (.D(_06482_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [941]),
    .QN(_31960_));
 DFF_X1 _65407_ (.D(_06483_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [942]),
    .QN(_31961_));
 DFF_X1 _65408_ (.D(_06484_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [943]),
    .QN(_31962_));
 DFF_X1 _65409_ (.D(_06485_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [944]),
    .QN(_31963_));
 DFF_X1 _65410_ (.D(_06486_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [945]),
    .QN(_31964_));
 DFF_X1 _65411_ (.D(_06487_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [946]),
    .QN(_31965_));
 DFF_X1 _65412_ (.D(_06488_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [947]),
    .QN(_31966_));
 DFF_X1 _65413_ (.D(_06489_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [948]),
    .QN(_31967_));
 DFF_X1 _65414_ (.D(_06490_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [949]),
    .QN(_31968_));
 DFF_X1 _65415_ (.D(_06492_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [950]),
    .QN(_31969_));
 DFF_X1 _65416_ (.D(_06493_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [951]),
    .QN(_31970_));
 DFF_X1 _65417_ (.D(_06494_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [952]),
    .QN(_31971_));
 DFF_X1 _65418_ (.D(_06495_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [953]),
    .QN(_31972_));
 DFF_X1 _65419_ (.D(_06496_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [954]),
    .QN(_31973_));
 DFF_X1 _65420_ (.D(_06497_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [955]),
    .QN(_31974_));
 DFF_X1 _65421_ (.D(_06498_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [956]),
    .QN(_31975_));
 DFF_X1 _65422_ (.D(_06499_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [957]),
    .QN(_31976_));
 DFF_X1 _65423_ (.D(_06500_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [958]),
    .QN(_31977_));
 DFF_X1 _65424_ (.D(_06501_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [959]),
    .QN(_31978_));
 DFF_X1 _65425_ (.D(_06503_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [960]),
    .QN(_31979_));
 DFF_X1 _65426_ (.D(_06504_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [961]),
    .QN(_31980_));
 DFF_X1 _65427_ (.D(_06505_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [962]),
    .QN(_31981_));
 DFF_X1 _65428_ (.D(_06506_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [963]),
    .QN(_31982_));
 DFF_X1 _65429_ (.D(_06507_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [964]),
    .QN(_31983_));
 DFF_X1 _65430_ (.D(_06508_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [965]),
    .QN(_31984_));
 DFF_X1 _65431_ (.D(_06509_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [966]),
    .QN(_31985_));
 DFF_X1 _65432_ (.D(_06510_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [967]),
    .QN(_31986_));
 DFF_X1 _65433_ (.D(_06511_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [968]),
    .QN(_31987_));
 DFF_X1 _65434_ (.D(_06512_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [969]),
    .QN(_31988_));
 DFF_X1 _65435_ (.D(_06514_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [970]),
    .QN(_31989_));
 DFF_X1 _65436_ (.D(_06515_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [971]),
    .QN(_31990_));
 DFF_X1 _65437_ (.D(_06516_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [972]),
    .QN(_31991_));
 DFF_X1 _65438_ (.D(_06517_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [973]),
    .QN(_31992_));
 DFF_X1 _65439_ (.D(_06518_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [974]),
    .QN(_31993_));
 DFF_X1 _65440_ (.D(_06519_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [975]),
    .QN(_31994_));
 DFF_X1 _65441_ (.D(_06520_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [976]),
    .QN(_31995_));
 DFF_X1 _65442_ (.D(_06521_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [977]),
    .QN(_31996_));
 DFF_X1 _65443_ (.D(_06522_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [978]),
    .QN(_31997_));
 DFF_X1 _65444_ (.D(_06523_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [979]),
    .QN(_31998_));
 DFF_X1 _65445_ (.D(_06525_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [980]),
    .QN(_31999_));
 DFF_X1 _65446_ (.D(_06526_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [981]),
    .QN(_32000_));
 DFF_X1 _65447_ (.D(_06527_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [982]),
    .QN(_32001_));
 DFF_X1 _65448_ (.D(_06528_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [983]),
    .QN(_32002_));
 DFF_X1 _65449_ (.D(_06529_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [984]),
    .QN(_32003_));
 DFF_X1 _65450_ (.D(_06530_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [985]),
    .QN(_32004_));
 DFF_X1 _65451_ (.D(_06531_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [986]),
    .QN(_32005_));
 DFF_X1 _65452_ (.D(_06532_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [987]),
    .QN(_32006_));
 DFF_X1 _65453_ (.D(_06533_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [988]),
    .QN(_32007_));
 DFF_X1 _65454_ (.D(_06534_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [989]),
    .QN(_32008_));
 DFF_X1 _65455_ (.D(_06536_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [990]),
    .QN(_32009_));
 DFF_X1 _65456_ (.D(_06537_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [991]),
    .QN(_32010_));
 DFF_X1 _65457_ (.D(_06538_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [992]),
    .QN(_32011_));
 DFF_X1 _65458_ (.D(_06539_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [993]),
    .QN(_32012_));
 DFF_X1 _65459_ (.D(_06540_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [994]),
    .QN(_32013_));
 DFF_X1 _65460_ (.D(_06541_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [995]),
    .QN(_32014_));
 DFF_X1 _65461_ (.D(_06542_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [996]),
    .QN(_32015_));
 DFF_X1 _65462_ (.D(_06543_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [997]),
    .QN(_32016_));
 DFF_X1 _65463_ (.D(_06544_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [998]),
    .QN(_32017_));
 DFF_X1 _65464_ (.D(_06545_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [999]),
    .QN(_32018_));
 DFF_X1 _65465_ (.D(_05515_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1000]),
    .QN(_32019_));
 DFF_X1 _65466_ (.D(_05516_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1001]),
    .QN(_32020_));
 DFF_X1 _65467_ (.D(_05517_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1002]),
    .QN(_32021_));
 DFF_X1 _65468_ (.D(_05518_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1003]),
    .QN(_32022_));
 DFF_X1 _65469_ (.D(_05519_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1004]),
    .QN(_32023_));
 DFF_X1 _65470_ (.D(_05520_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1005]),
    .QN(_32024_));
 DFF_X1 _65471_ (.D(_05521_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1006]),
    .QN(_32025_));
 DFF_X1 _65472_ (.D(_05522_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1007]),
    .QN(_32026_));
 DFF_X1 _65473_ (.D(_05523_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1008]),
    .QN(_32027_));
 DFF_X1 _65474_ (.D(_05524_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1009]),
    .QN(_32028_));
 DFF_X1 _65475_ (.D(_05526_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1010]),
    .QN(_32029_));
 DFF_X1 _65476_ (.D(_05527_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1011]),
    .QN(_32030_));
 DFF_X1 _65477_ (.D(_05528_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1012]),
    .QN(_32031_));
 DFF_X1 _65478_ (.D(_05529_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1013]),
    .QN(_32032_));
 DFF_X1 _65479_ (.D(_05530_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1014]),
    .QN(_32033_));
 DFF_X1 _65480_ (.D(_05531_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1015]),
    .QN(_32034_));
 DFF_X1 _65481_ (.D(_05532_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1016]),
    .QN(_32035_));
 DFF_X1 _65482_ (.D(_05533_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1017]),
    .QN(_32036_));
 DFF_X1 _65483_ (.D(_05534_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1018]),
    .QN(_32037_));
 DFF_X1 _65484_ (.D(_05535_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1019]),
    .QN(_32038_));
 DFF_X1 _65485_ (.D(_05537_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1020]),
    .QN(_32039_));
 DFF_X1 _65486_ (.D(_05538_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1021]),
    .QN(_32040_));
 DFF_X1 _65487_ (.D(_05539_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1022]),
    .QN(_32041_));
 DFF_X1 _65488_ (.D(_05540_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1023]),
    .QN(_32042_));
 DFF_X1 _65489_ (.D(_05541_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1024]),
    .QN(_32043_));
 DFF_X1 _65490_ (.D(_05542_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1025]),
    .QN(_32044_));
 DFF_X1 _65491_ (.D(_05543_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1026]),
    .QN(_32045_));
 DFF_X1 _65492_ (.D(_05544_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1027]),
    .QN(_32046_));
 DFF_X1 _65493_ (.D(_05545_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1028]),
    .QN(_32047_));
 DFF_X1 _65494_ (.D(_05546_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1029]),
    .QN(_32048_));
 DFF_X1 _65495_ (.D(_05548_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1030]),
    .QN(_32049_));
 DFF_X1 _65496_ (.D(_05549_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1031]),
    .QN(_32050_));
 DFF_X1 _65497_ (.D(_05550_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1032]),
    .QN(_32051_));
 DFF_X1 _65498_ (.D(_05551_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1033]),
    .QN(_32052_));
 DFF_X1 _65499_ (.D(_05552_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1034]),
    .QN(_32053_));
 DFF_X1 _65500_ (.D(_05553_),
    .CK(clk_i),
    .Q(\icache.lce.lce_data_cmd.rv_adapter.mem_1r1w.synth.mem [1035]),
    .QN(_32054_));
 DFF_X1 _65501_ (.D(N8),
    .CK(clk_i),
    .Q(itlb_fill_r),
    .QN(_00004_));
 DFF_X1 _65502_ (.D(_03958_),
    .CK(clk_i),
    .Q(\icache.addr_tv_r [0]),
    .QN(_32055_));
 DFF_X1 _65503_ (.D(_03969_),
    .CK(clk_i),
    .Q(\icache.addr_tv_r [1]),
    .QN(_32056_));
 DFF_X1 _65504_ (.D(_03980_),
    .CK(clk_i),
    .Q(\icache.N12 ),
    .QN(_32057_));
 DFF_X1 _65505_ (.D(_03990_),
    .CK(clk_i),
    .Q(\icache.addr_tv_r [3]),
    .QN(_32058_));
 DFF_X1 _65506_ (.D(_03991_),
    .CK(clk_i),
    .Q(\icache.addr_tv_r [4]),
    .QN(_32059_));
 DFF_X1 _65507_ (.D(_03992_),
    .CK(clk_i),
    .Q(\icache.addr_tv_r [5]),
    .QN(_32060_));
 DFF_X1 _65508_ (.D(_03993_),
    .CK(clk_i),
    .Q(\icache.addr_tv_r [6]),
    .QN(_32061_));
 DFF_X1 _65509_ (.D(_03994_),
    .CK(clk_i),
    .Q(\icache.addr_tv_r [7]),
    .QN(_32062_));
 DFF_X1 _65510_ (.D(_03995_),
    .CK(clk_i),
    .Q(\icache.addr_tv_r [8]),
    .QN(_32063_));
 DFF_X1 _65511_ (.D(_03996_),
    .CK(clk_i),
    .Q(\icache.addr_tv_r [9]),
    .QN(_32064_));
 DFF_X1 _65512_ (.D(_03959_),
    .CK(clk_i),
    .Q(\icache.addr_tv_r [10]),
    .QN(_32065_));
 DFF_X1 _65513_ (.D(_03960_),
    .CK(clk_i),
    .Q(\icache.addr_tv_r [11]),
    .QN(_32066_));
 DFF_X1 _65514_ (.D(_03961_),
    .CK(clk_i),
    .Q(\icache.addr_tv_r [12]),
    .QN(_32067_));
 DFF_X1 _65515_ (.D(_03962_),
    .CK(clk_i),
    .Q(\icache.addr_tv_r [13]),
    .QN(_32068_));
 DFF_X1 _65516_ (.D(_03963_),
    .CK(clk_i),
    .Q(\icache.addr_tv_r [14]),
    .QN(_32069_));
 DFF_X1 _65517_ (.D(_03964_),
    .CK(clk_i),
    .Q(\icache.addr_tv_r [15]),
    .QN(_32070_));
 DFF_X1 _65518_ (.D(_03965_),
    .CK(clk_i),
    .Q(\icache.addr_tv_r [16]),
    .QN(_32071_));
 DFF_X1 _65519_ (.D(_03966_),
    .CK(clk_i),
    .Q(\icache.addr_tv_r [17]),
    .QN(_32072_));
 DFF_X1 _65520_ (.D(_03967_),
    .CK(clk_i),
    .Q(\icache.addr_tv_r [18]),
    .QN(_32073_));
 DFF_X1 _65521_ (.D(_03968_),
    .CK(clk_i),
    .Q(\icache.addr_tv_r [19]),
    .QN(_32074_));
 DFF_X1 _65522_ (.D(_03970_),
    .CK(clk_i),
    .Q(\icache.addr_tv_r [20]),
    .QN(_32075_));
 DFF_X1 _65523_ (.D(_03971_),
    .CK(clk_i),
    .Q(\icache.addr_tv_r [21]),
    .QN(_32076_));
 DFF_X1 _65524_ (.D(_03972_),
    .CK(clk_i),
    .Q(\icache.addr_tv_r [22]),
    .QN(_32077_));
 DFF_X1 _65525_ (.D(_03973_),
    .CK(clk_i),
    .Q(\icache.addr_tv_r [23]),
    .QN(_32078_));
 DFF_X1 _65526_ (.D(_03974_),
    .CK(clk_i),
    .Q(\icache.addr_tv_r [24]),
    .QN(_32079_));
 DFF_X1 _65527_ (.D(_03975_),
    .CK(clk_i),
    .Q(\icache.addr_tv_r [25]),
    .QN(_32080_));
 DFF_X1 _65528_ (.D(_03976_),
    .CK(clk_i),
    .Q(\icache.addr_tv_r [26]),
    .QN(_32081_));
 DFF_X1 _65529_ (.D(_03977_),
    .CK(clk_i),
    .Q(\icache.addr_tv_r [27]),
    .QN(_32082_));
 DFF_X1 _65530_ (.D(_03978_),
    .CK(clk_i),
    .Q(\icache.addr_tv_r [28]),
    .QN(_32083_));
 DFF_X1 _65531_ (.D(_03979_),
    .CK(clk_i),
    .Q(\icache.addr_tv_r [29]),
    .QN(_32084_));
 DFF_X1 _65532_ (.D(_03981_),
    .CK(clk_i),
    .Q(\icache.addr_tv_r [30]),
    .QN(_32085_));
 DFF_X1 _65533_ (.D(_03982_),
    .CK(clk_i),
    .Q(\icache.addr_tv_r [31]),
    .QN(_32086_));
 DFF_X1 _65534_ (.D(_03983_),
    .CK(clk_i),
    .Q(\icache.addr_tv_r [32]),
    .QN(_32087_));
 DFF_X1 _65535_ (.D(_03984_),
    .CK(clk_i),
    .Q(\icache.addr_tv_r [33]),
    .QN(_32088_));
 DFF_X1 _65536_ (.D(_03985_),
    .CK(clk_i),
    .Q(\icache.addr_tv_r [34]),
    .QN(_32089_));
 DFF_X1 _65537_ (.D(_03986_),
    .CK(clk_i),
    .Q(\icache.addr_tv_r [35]),
    .QN(_32090_));
 DFF_X1 _65538_ (.D(_03987_),
    .CK(clk_i),
    .Q(\icache.addr_tv_r [36]),
    .QN(_32091_));
 DFF_X1 _65539_ (.D(_03988_),
    .CK(clk_i),
    .Q(\icache.addr_tv_r [37]),
    .QN(_32092_));
 DFF_X1 _65540_ (.D(_03989_),
    .CK(clk_i),
    .Q(\icache.addr_tv_r [38]),
    .QN(_32093_));
 DFF_X1 _65541_ (.D(_04783_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [64]),
    .QN(_00096_));
 DFF_X1 _65542_ (.D(_04794_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [65]),
    .QN(_00112_));
 DFF_X1 _65543_ (.D(_04805_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [66]),
    .QN(_00128_));
 DFF_X1 _65544_ (.D(_04816_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [67]),
    .QN(_00144_));
 DFF_X1 _65545_ (.D(_04827_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [68]),
    .QN(_00160_));
 DFF_X1 _65546_ (.D(_04838_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [69]),
    .QN(_00176_));
 DFF_X1 _65547_ (.D(_04843_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [70]),
    .QN(_00192_));
 DFF_X1 _65548_ (.D(_04844_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [71]),
    .QN(_00208_));
 DFF_X1 _65549_ (.D(_04845_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [72]),
    .QN(_00224_));
 DFF_X1 _65550_ (.D(_04846_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [73]),
    .QN(_00240_));
 DFF_X1 _65551_ (.D(_04784_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [74]),
    .QN(_00256_));
 DFF_X1 _65552_ (.D(_04785_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [75]),
    .QN(_00272_));
 DFF_X1 _65553_ (.D(_04786_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [76]),
    .QN(_00288_));
 DFF_X1 _65554_ (.D(_04787_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [77]),
    .QN(_00304_));
 DFF_X1 _65555_ (.D(_04788_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [78]),
    .QN(_00320_));
 DFF_X1 _65556_ (.D(_04789_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [79]),
    .QN(_00336_));
 DFF_X1 _65557_ (.D(_04790_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [80]),
    .QN(_00352_));
 DFF_X1 _65558_ (.D(_04791_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [81]),
    .QN(_00368_));
 DFF_X1 _65559_ (.D(_04792_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [82]),
    .QN(_00384_));
 DFF_X1 _65560_ (.D(_04793_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [83]),
    .QN(_00400_));
 DFF_X1 _65561_ (.D(_04795_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [84]),
    .QN(_00416_));
 DFF_X1 _65562_ (.D(_04796_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [85]),
    .QN(_00432_));
 DFF_X1 _65563_ (.D(_04797_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [86]),
    .QN(_00448_));
 DFF_X1 _65564_ (.D(_04798_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [87]),
    .QN(_00464_));
 DFF_X1 _65565_ (.D(_04799_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [88]),
    .QN(_00480_));
 DFF_X1 _65566_ (.D(_04800_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [89]),
    .QN(_00496_));
 DFF_X1 _65567_ (.D(_04801_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [90]),
    .QN(_00512_));
 DFF_X1 _65568_ (.D(_04802_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [91]),
    .QN(_00528_));
 DFF_X1 _65569_ (.D(_04803_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [92]),
    .QN(_00544_));
 DFF_X1 _65570_ (.D(_04804_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [93]),
    .QN(_00560_));
 DFF_X1 _65571_ (.D(_04806_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [94]),
    .QN(_32094_));
 DFF_X1 _65572_ (.D(_04807_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [95]),
    .QN(_32095_));
 DFF_X1 _65573_ (.D(_04808_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [96]),
    .QN(_00104_));
 DFF_X1 _65574_ (.D(_04809_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [97]),
    .QN(_00120_));
 DFF_X1 _65575_ (.D(_04810_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [98]),
    .QN(_00136_));
 DFF_X1 _65576_ (.D(_04811_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [99]),
    .QN(_00152_));
 DFF_X1 _65577_ (.D(_04812_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [100]),
    .QN(_00168_));
 DFF_X1 _65578_ (.D(_04813_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [101]),
    .QN(_00184_));
 DFF_X1 _65579_ (.D(_04814_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [102]),
    .QN(_00200_));
 DFF_X1 _65580_ (.D(_04815_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [103]),
    .QN(_00216_));
 DFF_X1 _65581_ (.D(_04817_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [104]),
    .QN(_00232_));
 DFF_X1 _65582_ (.D(_04818_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [105]),
    .QN(_00248_));
 DFF_X1 _65583_ (.D(_04819_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [106]),
    .QN(_00264_));
 DFF_X1 _65584_ (.D(_04820_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [107]),
    .QN(_00280_));
 DFF_X1 _65585_ (.D(_04821_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [108]),
    .QN(_00296_));
 DFF_X1 _65586_ (.D(_04822_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [109]),
    .QN(_00312_));
 DFF_X1 _65587_ (.D(_04823_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [110]),
    .QN(_00328_));
 DFF_X1 _65588_ (.D(_04824_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [111]),
    .QN(_00344_));
 DFF_X1 _65589_ (.D(_04825_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [112]),
    .QN(_00360_));
 DFF_X1 _65590_ (.D(_04826_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [113]),
    .QN(_00376_));
 DFF_X1 _65591_ (.D(_04828_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [114]),
    .QN(_00392_));
 DFF_X1 _65592_ (.D(_04829_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [115]),
    .QN(_00408_));
 DFF_X1 _65593_ (.D(_04830_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [116]),
    .QN(_00424_));
 DFF_X1 _65594_ (.D(_04831_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [117]),
    .QN(_00440_));
 DFF_X1 _65595_ (.D(_04832_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [118]),
    .QN(_00456_));
 DFF_X1 _65596_ (.D(_04833_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [119]),
    .QN(_00472_));
 DFF_X1 _65597_ (.D(_04834_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [120]),
    .QN(_00488_));
 DFF_X1 _65598_ (.D(_04835_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [121]),
    .QN(_00504_));
 DFF_X1 _65599_ (.D(_04836_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [122]),
    .QN(_00520_));
 DFF_X1 _65600_ (.D(_04837_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [123]),
    .QN(_00536_));
 DFF_X1 _65601_ (.D(_04839_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [124]),
    .QN(_00552_));
 DFF_X1 _65602_ (.D(_04840_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [125]),
    .QN(_00568_));
 DFF_X1 _65603_ (.D(_04841_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [126]),
    .QN(_32096_));
 DFF_X1 _65604_ (.D(_04842_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.data_i [127]),
    .QN(_32097_));
 DFF_X1 _65605_ (.D(_04036_),
    .CK(clk_i),
    .Q(\icache.read_mux_butterfly.mux_stage_0__mux_swap_0__swap_inst.N0 ),
    .QN(_32098_));
 DFF_X1 _65606_ (.D(_04037_),
    .CK(clk_i),
    .Q(\icache.read_mux_butterfly.mux_stage_1__mux_swap_0__swap_inst.N0 ),
    .QN(_32099_));
 DFF_X1 _65607_ (.D(_04038_),
    .CK(clk_i),
    .Q(\icache.read_mux_butterfly.mux_stage_2__mux_swap_0__swap_inst.N0 ),
    .QN(_32100_));
 DFF_X1 _65608_ (.D(_04551_),
    .CK(clk_i),
    .Q(\icache.state_tv_r [0]),
    .QN(_32101_));
 DFF_X1 _65609_ (.D(_04558_),
    .CK(clk_i),
    .Q(\icache.state_tv_r [1]),
    .QN(_32102_));
 DFF_X1 _65610_ (.D(_04559_),
    .CK(clk_i),
    .Q(\icache.state_tv_r [2]),
    .QN(_32103_));
 DFF_X1 _65611_ (.D(_04560_),
    .CK(clk_i),
    .Q(\icache.state_tv_r [3]),
    .QN(_32104_));
 DFF_X1 _65612_ (.D(_04561_),
    .CK(clk_i),
    .Q(\icache.state_tv_r [4]),
    .QN(_32105_));
 DFF_X1 _65613_ (.D(_04562_),
    .CK(clk_i),
    .Q(\icache.state_tv_r [5]),
    .QN(_32106_));
 DFF_X1 _65614_ (.D(_04563_),
    .CK(clk_i),
    .Q(\icache.state_tv_r [6]),
    .QN(_32107_));
 DFF_X1 _65615_ (.D(_04564_),
    .CK(clk_i),
    .Q(\icache.state_tv_r [7]),
    .QN(_32108_));
 DFF_X1 _65616_ (.D(_04565_),
    .CK(clk_i),
    .Q(\icache.state_tv_r [8]),
    .QN(_32109_));
 DFF_X1 _65617_ (.D(_04566_),
    .CK(clk_i),
    .Q(\icache.state_tv_r [9]),
    .QN(_32110_));
 DFF_X1 _65618_ (.D(_04552_),
    .CK(clk_i),
    .Q(\icache.state_tv_r [10]),
    .QN(_32111_));
 DFF_X1 _65619_ (.D(_04553_),
    .CK(clk_i),
    .Q(\icache.state_tv_r [11]),
    .QN(_32112_));
 DFF_X1 _65620_ (.D(_04554_),
    .CK(clk_i),
    .Q(\icache.state_tv_r [12]),
    .QN(_32113_));
 DFF_X1 _65621_ (.D(_04555_),
    .CK(clk_i),
    .Q(\icache.state_tv_r [13]),
    .QN(_32114_));
 DFF_X1 _65622_ (.D(_04556_),
    .CK(clk_i),
    .Q(\icache.state_tv_r [14]),
    .QN(_32115_));
 DFF_X1 _65623_ (.D(_04557_),
    .CK(clk_i),
    .Q(\icache.state_tv_r [15]),
    .QN(_32116_));
 DFF_X1 _65624_ (.D(_04567_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [0]),
    .QN(_32117_));
 DFF_X1 _65625_ (.D(_04678_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [1]),
    .QN(_32118_));
 DFF_X1 _65626_ (.D(_04705_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [2]),
    .QN(_32119_));
 DFF_X1 _65627_ (.D(_04716_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [3]),
    .QN(_32120_));
 DFF_X1 _65628_ (.D(_04727_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [4]),
    .QN(_32121_));
 DFF_X1 _65629_ (.D(_04738_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [5]),
    .QN(_32122_));
 DFF_X1 _65630_ (.D(_04749_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [6]),
    .QN(_32123_));
 DFF_X1 _65631_ (.D(_04760_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [7]),
    .QN(_32124_));
 DFF_X1 _65632_ (.D(_04771_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [8]),
    .QN(_32125_));
 DFF_X1 _65633_ (.D(_04782_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [9]),
    .QN(_32126_));
 DFF_X1 _65634_ (.D(_04578_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [10]),
    .QN(_32127_));
 DFF_X1 _65635_ (.D(_04589_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [11]),
    .QN(_32128_));
 DFF_X1 _65636_ (.D(_04600_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [12]),
    .QN(_32129_));
 DFF_X1 _65637_ (.D(_04611_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [13]),
    .QN(_32130_));
 DFF_X1 _65638_ (.D(_04622_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [14]),
    .QN(_32131_));
 DFF_X1 _65639_ (.D(_04633_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [15]),
    .QN(_32132_));
 DFF_X1 _65640_ (.D(_04644_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [16]),
    .QN(_32133_));
 DFF_X1 _65641_ (.D(_04655_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [17]),
    .QN(_32134_));
 DFF_X1 _65642_ (.D(_04666_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [18]),
    .QN(_32135_));
 DFF_X1 _65643_ (.D(_04677_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [19]),
    .QN(_32136_));
 DFF_X1 _65644_ (.D(_04689_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [20]),
    .QN(_32137_));
 DFF_X1 _65645_ (.D(_04696_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [21]),
    .QN(_32138_));
 DFF_X1 _65646_ (.D(_04697_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [22]),
    .QN(_32139_));
 DFF_X1 _65647_ (.D(_04698_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [23]),
    .QN(_32140_));
 DFF_X1 _65648_ (.D(_04699_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [24]),
    .QN(_32141_));
 DFF_X1 _65649_ (.D(_04700_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [25]),
    .QN(_32142_));
 DFF_X1 _65650_ (.D(_04701_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [26]),
    .QN(_32143_));
 DFF_X1 _65651_ (.D(_04702_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [27]),
    .QN(_32144_));
 DFF_X1 _65652_ (.D(_04703_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [28]),
    .QN(_32145_));
 DFF_X1 _65653_ (.D(_04704_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [29]),
    .QN(_32146_));
 DFF_X1 _65654_ (.D(_04706_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [30]),
    .QN(_32147_));
 DFF_X1 _65655_ (.D(_04707_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [31]),
    .QN(_32148_));
 DFF_X1 _65656_ (.D(_04708_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [32]),
    .QN(_32149_));
 DFF_X1 _65657_ (.D(_04709_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [33]),
    .QN(_32150_));
 DFF_X1 _65658_ (.D(_04710_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [34]),
    .QN(_32151_));
 DFF_X1 _65659_ (.D(_04711_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [35]),
    .QN(_32152_));
 DFF_X1 _65660_ (.D(_04712_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [36]),
    .QN(_32153_));
 DFF_X1 _65661_ (.D(_04713_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [37]),
    .QN(_32154_));
 DFF_X1 _65662_ (.D(_04714_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [38]),
    .QN(_32155_));
 DFF_X1 _65663_ (.D(_04715_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [39]),
    .QN(_32156_));
 DFF_X1 _65664_ (.D(_04717_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [40]),
    .QN(_32157_));
 DFF_X1 _65665_ (.D(_04718_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [41]),
    .QN(_32158_));
 DFF_X1 _65666_ (.D(_04719_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [42]),
    .QN(_32159_));
 DFF_X1 _65667_ (.D(_04720_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [43]),
    .QN(_32160_));
 DFF_X1 _65668_ (.D(_04721_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [44]),
    .QN(_32161_));
 DFF_X1 _65669_ (.D(_04722_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [45]),
    .QN(_32162_));
 DFF_X1 _65670_ (.D(_04723_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [46]),
    .QN(_32163_));
 DFF_X1 _65671_ (.D(_04724_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [47]),
    .QN(_32164_));
 DFF_X1 _65672_ (.D(_04725_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [48]),
    .QN(_32165_));
 DFF_X1 _65673_ (.D(_04726_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [49]),
    .QN(_32166_));
 DFF_X1 _65674_ (.D(_04728_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [50]),
    .QN(_32167_));
 DFF_X1 _65675_ (.D(_04729_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [51]),
    .QN(_32168_));
 DFF_X1 _65676_ (.D(_04730_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [52]),
    .QN(_32169_));
 DFF_X1 _65677_ (.D(_04731_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [53]),
    .QN(_32170_));
 DFF_X1 _65678_ (.D(_04732_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [54]),
    .QN(_32171_));
 DFF_X1 _65679_ (.D(_04733_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [55]),
    .QN(_32172_));
 DFF_X1 _65680_ (.D(_04734_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [56]),
    .QN(_32173_));
 DFF_X1 _65681_ (.D(_04735_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [57]),
    .QN(_32174_));
 DFF_X1 _65682_ (.D(_04736_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [58]),
    .QN(_32175_));
 DFF_X1 _65683_ (.D(_04737_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [59]),
    .QN(_32176_));
 DFF_X1 _65684_ (.D(_04739_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [60]),
    .QN(_32177_));
 DFF_X1 _65685_ (.D(_04740_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [61]),
    .QN(_32178_));
 DFF_X1 _65686_ (.D(_04741_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [62]),
    .QN(_32179_));
 DFF_X1 _65687_ (.D(_04742_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [63]),
    .QN(_32180_));
 DFF_X1 _65688_ (.D(_04743_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [64]),
    .QN(_32181_));
 DFF_X1 _65689_ (.D(_04744_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [65]),
    .QN(_32182_));
 DFF_X1 _65690_ (.D(_04745_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [66]),
    .QN(_32183_));
 DFF_X1 _65691_ (.D(_04746_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [67]),
    .QN(_32184_));
 DFF_X1 _65692_ (.D(_04747_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [68]),
    .QN(_32185_));
 DFF_X1 _65693_ (.D(_04748_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [69]),
    .QN(_32186_));
 DFF_X1 _65694_ (.D(_04750_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [70]),
    .QN(_32187_));
 DFF_X1 _65695_ (.D(_04751_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [71]),
    .QN(_32188_));
 DFF_X1 _65696_ (.D(_04752_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [72]),
    .QN(_32189_));
 DFF_X1 _65697_ (.D(_04753_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [73]),
    .QN(_32190_));
 DFF_X1 _65698_ (.D(_04754_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [74]),
    .QN(_32191_));
 DFF_X1 _65699_ (.D(_04755_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [75]),
    .QN(_32192_));
 DFF_X1 _65700_ (.D(_04756_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [76]),
    .QN(_32193_));
 DFF_X1 _65701_ (.D(_04757_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [77]),
    .QN(_32194_));
 DFF_X1 _65702_ (.D(_04758_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [78]),
    .QN(_32195_));
 DFF_X1 _65703_ (.D(_04759_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [79]),
    .QN(_32196_));
 DFF_X1 _65704_ (.D(_04761_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [80]),
    .QN(_32197_));
 DFF_X1 _65705_ (.D(_04762_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [81]),
    .QN(_32198_));
 DFF_X1 _65706_ (.D(_04763_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [82]),
    .QN(_32199_));
 DFF_X1 _65707_ (.D(_04764_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [83]),
    .QN(_32200_));
 DFF_X1 _65708_ (.D(_04765_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [84]),
    .QN(_32201_));
 DFF_X1 _65709_ (.D(_04766_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [85]),
    .QN(_32202_));
 DFF_X1 _65710_ (.D(_04767_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [86]),
    .QN(_32203_));
 DFF_X1 _65711_ (.D(_04768_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [87]),
    .QN(_32204_));
 DFF_X1 _65712_ (.D(_04769_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [88]),
    .QN(_32205_));
 DFF_X1 _65713_ (.D(_04770_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [89]),
    .QN(_32206_));
 DFF_X1 _65714_ (.D(_04772_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [90]),
    .QN(_32207_));
 DFF_X1 _65715_ (.D(_04773_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [91]),
    .QN(_32208_));
 DFF_X1 _65716_ (.D(_04774_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [92]),
    .QN(_32209_));
 DFF_X1 _65717_ (.D(_04775_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [93]),
    .QN(_32210_));
 DFF_X1 _65718_ (.D(_04776_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [94]),
    .QN(_32211_));
 DFF_X1 _65719_ (.D(_04777_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [95]),
    .QN(_32212_));
 DFF_X1 _65720_ (.D(_04778_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [96]),
    .QN(_32213_));
 DFF_X1 _65721_ (.D(_04779_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [97]),
    .QN(_32214_));
 DFF_X1 _65722_ (.D(_04780_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [98]),
    .QN(_32215_));
 DFF_X1 _65723_ (.D(_04781_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [99]),
    .QN(_32216_));
 DFF_X1 _65724_ (.D(_04568_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [100]),
    .QN(_32217_));
 DFF_X1 _65725_ (.D(_04569_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [101]),
    .QN(_32218_));
 DFF_X1 _65726_ (.D(_04570_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [102]),
    .QN(_32219_));
 DFF_X1 _65727_ (.D(_04571_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [103]),
    .QN(_32220_));
 DFF_X1 _65728_ (.D(_04572_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [104]),
    .QN(_32221_));
 DFF_X1 _65729_ (.D(_04573_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [105]),
    .QN(_32222_));
 DFF_X1 _65730_ (.D(_04574_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [106]),
    .QN(_32223_));
 DFF_X1 _65731_ (.D(_04575_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [107]),
    .QN(_32224_));
 DFF_X1 _65732_ (.D(_04576_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [108]),
    .QN(_32225_));
 DFF_X1 _65733_ (.D(_04577_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [109]),
    .QN(_32226_));
 DFF_X1 _65734_ (.D(_04579_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [110]),
    .QN(_32227_));
 DFF_X1 _65735_ (.D(_04580_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [111]),
    .QN(_32228_));
 DFF_X1 _65736_ (.D(_04581_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [112]),
    .QN(_32229_));
 DFF_X1 _65737_ (.D(_04582_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [113]),
    .QN(_32230_));
 DFF_X1 _65738_ (.D(_04583_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [114]),
    .QN(_32231_));
 DFF_X1 _65739_ (.D(_04584_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [115]),
    .QN(_32232_));
 DFF_X1 _65740_ (.D(_04585_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [116]),
    .QN(_32233_));
 DFF_X1 _65741_ (.D(_04586_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [117]),
    .QN(_32234_));
 DFF_X1 _65742_ (.D(_04587_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [118]),
    .QN(_32235_));
 DFF_X1 _65743_ (.D(_04588_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [119]),
    .QN(_32236_));
 DFF_X1 _65744_ (.D(_04590_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [120]),
    .QN(_32237_));
 DFF_X1 _65745_ (.D(_04591_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [121]),
    .QN(_32238_));
 DFF_X1 _65746_ (.D(_04592_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [122]),
    .QN(_32239_));
 DFF_X1 _65747_ (.D(_04593_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [123]),
    .QN(_32240_));
 DFF_X1 _65748_ (.D(_04594_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [124]),
    .QN(_32241_));
 DFF_X1 _65749_ (.D(_04595_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [125]),
    .QN(_32242_));
 DFF_X1 _65750_ (.D(_04596_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [126]),
    .QN(_32243_));
 DFF_X1 _65751_ (.D(_04597_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [127]),
    .QN(_32244_));
 DFF_X1 _65752_ (.D(_04598_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [128]),
    .QN(_32245_));
 DFF_X1 _65753_ (.D(_04599_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [129]),
    .QN(_32246_));
 DFF_X1 _65754_ (.D(_04601_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [130]),
    .QN(_32247_));
 DFF_X1 _65755_ (.D(_04602_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [131]),
    .QN(_32248_));
 DFF_X1 _65756_ (.D(_04603_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [132]),
    .QN(_32249_));
 DFF_X1 _65757_ (.D(_04604_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [133]),
    .QN(_32250_));
 DFF_X1 _65758_ (.D(_04605_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [134]),
    .QN(_32251_));
 DFF_X1 _65759_ (.D(_04606_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [135]),
    .QN(_32252_));
 DFF_X1 _65760_ (.D(_04607_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [136]),
    .QN(_32253_));
 DFF_X1 _65761_ (.D(_04608_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [137]),
    .QN(_32254_));
 DFF_X1 _65762_ (.D(_04609_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [138]),
    .QN(_32255_));
 DFF_X1 _65763_ (.D(_04610_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [139]),
    .QN(_32256_));
 DFF_X1 _65764_ (.D(_04612_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [140]),
    .QN(_32257_));
 DFF_X1 _65765_ (.D(_04613_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [141]),
    .QN(_32258_));
 DFF_X1 _65766_ (.D(_04614_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [142]),
    .QN(_32259_));
 DFF_X1 _65767_ (.D(_04615_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [143]),
    .QN(_32260_));
 DFF_X1 _65768_ (.D(_04616_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [144]),
    .QN(_32261_));
 DFF_X1 _65769_ (.D(_04617_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [145]),
    .QN(_32262_));
 DFF_X1 _65770_ (.D(_04618_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [146]),
    .QN(_32263_));
 DFF_X1 _65771_ (.D(_04619_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [147]),
    .QN(_32264_));
 DFF_X1 _65772_ (.D(_04620_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [148]),
    .QN(_32265_));
 DFF_X1 _65773_ (.D(_04621_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [149]),
    .QN(_32266_));
 DFF_X1 _65774_ (.D(_04623_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [150]),
    .QN(_32267_));
 DFF_X1 _65775_ (.D(_04624_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [151]),
    .QN(_32268_));
 DFF_X1 _65776_ (.D(_04625_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [152]),
    .QN(_32269_));
 DFF_X1 _65777_ (.D(_04626_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [153]),
    .QN(_32270_));
 DFF_X1 _65778_ (.D(_04627_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [154]),
    .QN(_32271_));
 DFF_X1 _65779_ (.D(_04628_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [155]),
    .QN(_32272_));
 DFF_X1 _65780_ (.D(_04629_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [156]),
    .QN(_32273_));
 DFF_X1 _65781_ (.D(_04630_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [157]),
    .QN(_32274_));
 DFF_X1 _65782_ (.D(_04631_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [158]),
    .QN(_32275_));
 DFF_X1 _65783_ (.D(_04632_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [159]),
    .QN(_32276_));
 DFF_X1 _65784_ (.D(_04634_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [160]),
    .QN(_32277_));
 DFF_X1 _65785_ (.D(_04635_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [161]),
    .QN(_32278_));
 DFF_X1 _65786_ (.D(_04636_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [162]),
    .QN(_32279_));
 DFF_X1 _65787_ (.D(_04637_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [163]),
    .QN(_32280_));
 DFF_X1 _65788_ (.D(_04638_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [164]),
    .QN(_32281_));
 DFF_X1 _65789_ (.D(_04639_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [165]),
    .QN(_32282_));
 DFF_X1 _65790_ (.D(_04640_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [166]),
    .QN(_32283_));
 DFF_X1 _65791_ (.D(_04641_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [167]),
    .QN(_32284_));
 DFF_X1 _65792_ (.D(_04642_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [168]),
    .QN(_32285_));
 DFF_X1 _65793_ (.D(_04643_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [169]),
    .QN(_32286_));
 DFF_X1 _65794_ (.D(_04645_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [170]),
    .QN(_32287_));
 DFF_X1 _65795_ (.D(_04646_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [171]),
    .QN(_32288_));
 DFF_X1 _65796_ (.D(_04647_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [172]),
    .QN(_32289_));
 DFF_X1 _65797_ (.D(_04648_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [173]),
    .QN(_32290_));
 DFF_X1 _65798_ (.D(_04649_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [174]),
    .QN(_32291_));
 DFF_X1 _65799_ (.D(_04650_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [175]),
    .QN(_32292_));
 DFF_X1 _65800_ (.D(_04651_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [176]),
    .QN(_32293_));
 DFF_X1 _65801_ (.D(_04652_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [177]),
    .QN(_32294_));
 DFF_X1 _65802_ (.D(_04653_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [178]),
    .QN(_32295_));
 DFF_X1 _65803_ (.D(_04654_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [179]),
    .QN(_32296_));
 DFF_X1 _65804_ (.D(_04656_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [180]),
    .QN(_32297_));
 DFF_X1 _65805_ (.D(_04657_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [181]),
    .QN(_32298_));
 DFF_X1 _65806_ (.D(_04658_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [182]),
    .QN(_32299_));
 DFF_X1 _65807_ (.D(_04659_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [183]),
    .QN(_32300_));
 DFF_X1 _65808_ (.D(_04660_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [184]),
    .QN(_32301_));
 DFF_X1 _65809_ (.D(_04661_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [185]),
    .QN(_32302_));
 DFF_X1 _65810_ (.D(_04662_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [186]),
    .QN(_32303_));
 DFF_X1 _65811_ (.D(_04663_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [187]),
    .QN(_32304_));
 DFF_X1 _65812_ (.D(_04664_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [188]),
    .QN(_32305_));
 DFF_X1 _65813_ (.D(_04665_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [189]),
    .QN(_32306_));
 DFF_X1 _65814_ (.D(_04667_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [190]),
    .QN(_32307_));
 DFF_X1 _65815_ (.D(_04668_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [191]),
    .QN(_32308_));
 DFF_X1 _65816_ (.D(_04669_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [192]),
    .QN(_32309_));
 DFF_X1 _65817_ (.D(_04670_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [193]),
    .QN(_32310_));
 DFF_X1 _65818_ (.D(_04671_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [194]),
    .QN(_32311_));
 DFF_X1 _65819_ (.D(_04672_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [195]),
    .QN(_32312_));
 DFF_X1 _65820_ (.D(_04673_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [196]),
    .QN(_32313_));
 DFF_X1 _65821_ (.D(_04674_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [197]),
    .QN(_32314_));
 DFF_X1 _65822_ (.D(_04675_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [198]),
    .QN(_32315_));
 DFF_X1 _65823_ (.D(_04676_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [199]),
    .QN(_32316_));
 DFF_X1 _65824_ (.D(_04679_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [200]),
    .QN(_32317_));
 DFF_X1 _65825_ (.D(_04680_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [201]),
    .QN(_32318_));
 DFF_X1 _65826_ (.D(_04681_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [202]),
    .QN(_32319_));
 DFF_X1 _65827_ (.D(_04682_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [203]),
    .QN(_32320_));
 DFF_X1 _65828_ (.D(_04683_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [204]),
    .QN(_32321_));
 DFF_X1 _65829_ (.D(_04684_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [205]),
    .QN(_32322_));
 DFF_X1 _65830_ (.D(_04685_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [206]),
    .QN(_32323_));
 DFF_X1 _65831_ (.D(_04686_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [207]),
    .QN(_32324_));
 DFF_X1 _65832_ (.D(_04687_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [208]),
    .QN(_32325_));
 DFF_X1 _65833_ (.D(_04688_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [209]),
    .QN(_32326_));
 DFF_X1 _65834_ (.D(_04690_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [210]),
    .QN(_32327_));
 DFF_X1 _65835_ (.D(_04691_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [211]),
    .QN(_32328_));
 DFF_X1 _65836_ (.D(_04692_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [212]),
    .QN(_32329_));
 DFF_X1 _65837_ (.D(_04693_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [213]),
    .QN(_32330_));
 DFF_X1 _65838_ (.D(_04694_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [214]),
    .QN(_32331_));
 DFF_X1 _65839_ (.D(_04695_),
    .CK(clk_i),
    .Q(\icache.tag_tv_r [215]),
    .QN(_32332_));
 DFF_X1 _65840_ (.D(_04039_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [0]),
    .QN(_00097_));
 DFF_X1 _65841_ (.D(_04150_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [1]),
    .QN(_00113_));
 DFF_X1 _65842_ (.D(_04261_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [2]),
    .QN(_00129_));
 DFF_X1 _65843_ (.D(_04372_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [3]),
    .QN(_00145_));
 DFF_X1 _65844_ (.D(_04483_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [4]),
    .QN(_00161_));
 DFF_X1 _65845_ (.D(_04506_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [5]),
    .QN(_00177_));
 DFF_X1 _65846_ (.D(_04517_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [6]),
    .QN(_00193_));
 DFF_X1 _65847_ (.D(_04528_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [7]),
    .QN(_00209_));
 DFF_X1 _65848_ (.D(_04539_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [8]),
    .QN(_00225_));
 DFF_X1 _65849_ (.D(_04550_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [9]),
    .QN(_00241_));
 DFF_X1 _65850_ (.D(_04050_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [10]),
    .QN(_00257_));
 DFF_X1 _65851_ (.D(_04061_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [11]),
    .QN(_00273_));
 DFF_X1 _65852_ (.D(_04072_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [12]),
    .QN(_00289_));
 DFF_X1 _65853_ (.D(_04083_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [13]),
    .QN(_00305_));
 DFF_X1 _65854_ (.D(_04094_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [14]),
    .QN(_00321_));
 DFF_X1 _65855_ (.D(_04105_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [15]),
    .QN(_00337_));
 DFF_X1 _65856_ (.D(_04116_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [16]),
    .QN(_00353_));
 DFF_X1 _65857_ (.D(_04127_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [17]),
    .QN(_00369_));
 DFF_X1 _65858_ (.D(_04138_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [18]),
    .QN(_00385_));
 DFF_X1 _65859_ (.D(_04149_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [19]),
    .QN(_00401_));
 DFF_X1 _65860_ (.D(_04161_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [20]),
    .QN(_00417_));
 DFF_X1 _65861_ (.D(_04172_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [21]),
    .QN(_00433_));
 DFF_X1 _65862_ (.D(_04183_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [22]),
    .QN(_00449_));
 DFF_X1 _65863_ (.D(_04194_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [23]),
    .QN(_00465_));
 DFF_X1 _65864_ (.D(_04205_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [24]),
    .QN(_00481_));
 DFF_X1 _65865_ (.D(_04216_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [25]),
    .QN(_00497_));
 DFF_X1 _65866_ (.D(_04227_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [26]),
    .QN(_00513_));
 DFF_X1 _65867_ (.D(_04238_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [27]),
    .QN(_00529_));
 DFF_X1 _65868_ (.D(_04249_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [28]),
    .QN(_00545_));
 DFF_X1 _65869_ (.D(_04260_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [29]),
    .QN(_00561_));
 DFF_X1 _65870_ (.D(_04272_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [30]),
    .QN(_32333_));
 DFF_X1 _65871_ (.D(_04283_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [31]),
    .QN(_32334_));
 DFF_X1 _65872_ (.D(_04294_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [32]),
    .QN(_00105_));
 DFF_X1 _65873_ (.D(_04305_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [33]),
    .QN(_00121_));
 DFF_X1 _65874_ (.D(_04316_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [34]),
    .QN(_00137_));
 DFF_X1 _65875_ (.D(_04327_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [35]),
    .QN(_00153_));
 DFF_X1 _65876_ (.D(_04338_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [36]),
    .QN(_00169_));
 DFF_X1 _65877_ (.D(_04349_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [37]),
    .QN(_00185_));
 DFF_X1 _65878_ (.D(_04360_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [38]),
    .QN(_00201_));
 DFF_X1 _65879_ (.D(_04371_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [39]),
    .QN(_00217_));
 DFF_X1 _65880_ (.D(_04383_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [40]),
    .QN(_00233_));
 DFF_X1 _65881_ (.D(_04394_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [41]),
    .QN(_00249_));
 DFF_X1 _65882_ (.D(_04405_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [42]),
    .QN(_00265_));
 DFF_X1 _65883_ (.D(_04416_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [43]),
    .QN(_00281_));
 DFF_X1 _65884_ (.D(_04427_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [44]),
    .QN(_00297_));
 DFF_X1 _65885_ (.D(_04438_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [45]),
    .QN(_00313_));
 DFF_X1 _65886_ (.D(_04449_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [46]),
    .QN(_00329_));
 DFF_X1 _65887_ (.D(_04460_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [47]),
    .QN(_00345_));
 DFF_X1 _65888_ (.D(_04471_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [48]),
    .QN(_00361_));
 DFF_X1 _65889_ (.D(_04482_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [49]),
    .QN(_00377_));
 DFF_X1 _65890_ (.D(_04494_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [50]),
    .QN(_00393_));
 DFF_X1 _65891_ (.D(_04497_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [51]),
    .QN(_00409_));
 DFF_X1 _65892_ (.D(_04498_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [52]),
    .QN(_00425_));
 DFF_X1 _65893_ (.D(_04499_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [53]),
    .QN(_00441_));
 DFF_X1 _65894_ (.D(_04500_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [54]),
    .QN(_00457_));
 DFF_X1 _65895_ (.D(_04501_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [55]),
    .QN(_00473_));
 DFF_X1 _65896_ (.D(_04502_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [56]),
    .QN(_00489_));
 DFF_X1 _65897_ (.D(_04503_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [57]),
    .QN(_00505_));
 DFF_X1 _65898_ (.D(_04504_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [58]),
    .QN(_00521_));
 DFF_X1 _65899_ (.D(_04505_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [59]),
    .QN(_00537_));
 DFF_X1 _65900_ (.D(_04507_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [60]),
    .QN(_00553_));
 DFF_X1 _65901_ (.D(_04508_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [61]),
    .QN(_00569_));
 DFF_X1 _65902_ (.D(_04509_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [62]),
    .QN(_32335_));
 DFF_X1 _65903_ (.D(_04510_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [63]),
    .QN(_32336_));
 DFF_X1 _65904_ (.D(_04511_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [64]),
    .QN(_00098_));
 DFF_X1 _65905_ (.D(_04512_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [65]),
    .QN(_00114_));
 DFF_X1 _65906_ (.D(_04513_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [66]),
    .QN(_00130_));
 DFF_X1 _65907_ (.D(_04514_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [67]),
    .QN(_00146_));
 DFF_X1 _65908_ (.D(_04515_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [68]),
    .QN(_00162_));
 DFF_X1 _65909_ (.D(_04516_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [69]),
    .QN(_00178_));
 DFF_X1 _65910_ (.D(_04518_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [70]),
    .QN(_00194_));
 DFF_X1 _65911_ (.D(_04519_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [71]),
    .QN(_00210_));
 DFF_X1 _65912_ (.D(_04520_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [72]),
    .QN(_00226_));
 DFF_X1 _65913_ (.D(_04521_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [73]),
    .QN(_00242_));
 DFF_X1 _65914_ (.D(_04522_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [74]),
    .QN(_00258_));
 DFF_X1 _65915_ (.D(_04523_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [75]),
    .QN(_00274_));
 DFF_X1 _65916_ (.D(_04524_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [76]),
    .QN(_00290_));
 DFF_X1 _65917_ (.D(_04525_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [77]),
    .QN(_00306_));
 DFF_X1 _65918_ (.D(_04526_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [78]),
    .QN(_00322_));
 DFF_X1 _65919_ (.D(_04527_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [79]),
    .QN(_00338_));
 DFF_X1 _65920_ (.D(_04529_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [80]),
    .QN(_00354_));
 DFF_X1 _65921_ (.D(_04530_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [81]),
    .QN(_00370_));
 DFF_X1 _65922_ (.D(_04531_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [82]),
    .QN(_00386_));
 DFF_X1 _65923_ (.D(_04532_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [83]),
    .QN(_00402_));
 DFF_X1 _65924_ (.D(_04533_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [84]),
    .QN(_00418_));
 DFF_X1 _65925_ (.D(_04534_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [85]),
    .QN(_00434_));
 DFF_X1 _65926_ (.D(_04535_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [86]),
    .QN(_00450_));
 DFF_X1 _65927_ (.D(_04536_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [87]),
    .QN(_00466_));
 DFF_X1 _65928_ (.D(_04537_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [88]),
    .QN(_00482_));
 DFF_X1 _65929_ (.D(_04538_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [89]),
    .QN(_00498_));
 DFF_X1 _65930_ (.D(_04540_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [90]),
    .QN(_00514_));
 DFF_X1 _65931_ (.D(_04541_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [91]),
    .QN(_00530_));
 DFF_X1 _65932_ (.D(_04542_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [92]),
    .QN(_00546_));
 DFF_X1 _65933_ (.D(_04543_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [93]),
    .QN(_00562_));
 DFF_X1 _65934_ (.D(_04544_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [94]),
    .QN(_32337_));
 DFF_X1 _65935_ (.D(_04545_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [95]),
    .QN(_32338_));
 DFF_X1 _65936_ (.D(_04546_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [96]),
    .QN(_00106_));
 DFF_X1 _65937_ (.D(_04547_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [97]),
    .QN(_00122_));
 DFF_X1 _65938_ (.D(_04548_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [98]),
    .QN(_00138_));
 DFF_X1 _65939_ (.D(_04549_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [99]),
    .QN(_00154_));
 DFF_X1 _65940_ (.D(_04040_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [100]),
    .QN(_00170_));
 DFF_X1 _65941_ (.D(_04041_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [101]),
    .QN(_00186_));
 DFF_X1 _65942_ (.D(_04042_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [102]),
    .QN(_00202_));
 DFF_X1 _65943_ (.D(_04043_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [103]),
    .QN(_00218_));
 DFF_X1 _65944_ (.D(_04044_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [104]),
    .QN(_00234_));
 DFF_X1 _65945_ (.D(_04045_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [105]),
    .QN(_00250_));
 DFF_X1 _65946_ (.D(_04046_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [106]),
    .QN(_00266_));
 DFF_X1 _65947_ (.D(_04047_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [107]),
    .QN(_00282_));
 DFF_X1 _65948_ (.D(_04048_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [108]),
    .QN(_00298_));
 DFF_X1 _65949_ (.D(_04049_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [109]),
    .QN(_00314_));
 DFF_X1 _65950_ (.D(_04051_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [110]),
    .QN(_00330_));
 DFF_X1 _65951_ (.D(_04052_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [111]),
    .QN(_00346_));
 DFF_X1 _65952_ (.D(_04053_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [112]),
    .QN(_00362_));
 DFF_X1 _65953_ (.D(_04054_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [113]),
    .QN(_00378_));
 DFF_X1 _65954_ (.D(_04055_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [114]),
    .QN(_00394_));
 DFF_X1 _65955_ (.D(_04056_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [115]),
    .QN(_00410_));
 DFF_X1 _65956_ (.D(_04057_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [116]),
    .QN(_00426_));
 DFF_X1 _65957_ (.D(_04058_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [117]),
    .QN(_00442_));
 DFF_X1 _65958_ (.D(_04059_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [118]),
    .QN(_00458_));
 DFF_X1 _65959_ (.D(_04060_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [119]),
    .QN(_00474_));
 DFF_X1 _65960_ (.D(_04062_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [120]),
    .QN(_00490_));
 DFF_X1 _65961_ (.D(_04063_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [121]),
    .QN(_00506_));
 DFF_X1 _65962_ (.D(_04064_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [122]),
    .QN(_00522_));
 DFF_X1 _65963_ (.D(_04065_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [123]),
    .QN(_00538_));
 DFF_X1 _65964_ (.D(_04066_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [124]),
    .QN(_00554_));
 DFF_X1 _65965_ (.D(_04067_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [125]),
    .QN(_00570_));
 DFF_X1 _65966_ (.D(_04068_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [126]),
    .QN(_32339_));
 DFF_X1 _65967_ (.D(_04069_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [127]),
    .QN(_32340_));
 DFF_X1 _65968_ (.D(_04070_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [128]),
    .QN(_00099_));
 DFF_X1 _65969_ (.D(_04071_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [129]),
    .QN(_00115_));
 DFF_X1 _65970_ (.D(_04073_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [130]),
    .QN(_00131_));
 DFF_X1 _65971_ (.D(_04074_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [131]),
    .QN(_00147_));
 DFF_X1 _65972_ (.D(_04075_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [132]),
    .QN(_00163_));
 DFF_X1 _65973_ (.D(_04076_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [133]),
    .QN(_00179_));
 DFF_X1 _65974_ (.D(_04077_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [134]),
    .QN(_00195_));
 DFF_X1 _65975_ (.D(_04078_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [135]),
    .QN(_00211_));
 DFF_X1 _65976_ (.D(_04079_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [136]),
    .QN(_00227_));
 DFF_X1 _65977_ (.D(_04080_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [137]),
    .QN(_00243_));
 DFF_X1 _65978_ (.D(_04081_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [138]),
    .QN(_00259_));
 DFF_X1 _65979_ (.D(_04082_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [139]),
    .QN(_00275_));
 DFF_X1 _65980_ (.D(_04084_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [140]),
    .QN(_00291_));
 DFF_X1 _65981_ (.D(_04085_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [141]),
    .QN(_00307_));
 DFF_X1 _65982_ (.D(_04086_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [142]),
    .QN(_00323_));
 DFF_X1 _65983_ (.D(_04087_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [143]),
    .QN(_00339_));
 DFF_X1 _65984_ (.D(_04088_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [144]),
    .QN(_00355_));
 DFF_X1 _65985_ (.D(_04089_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [145]),
    .QN(_00371_));
 DFF_X1 _65986_ (.D(_04090_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [146]),
    .QN(_00387_));
 DFF_X1 _65987_ (.D(_04091_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [147]),
    .QN(_00403_));
 DFF_X1 _65988_ (.D(_04092_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [148]),
    .QN(_00419_));
 DFF_X1 _65989_ (.D(_04093_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [149]),
    .QN(_00435_));
 DFF_X1 _65990_ (.D(_04095_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [150]),
    .QN(_00451_));
 DFF_X1 _65991_ (.D(_04096_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [151]),
    .QN(_00467_));
 DFF_X1 _65992_ (.D(_04097_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [152]),
    .QN(_00483_));
 DFF_X1 _65993_ (.D(_04098_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [153]),
    .QN(_00499_));
 DFF_X1 _65994_ (.D(_04099_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [154]),
    .QN(_00515_));
 DFF_X1 _65995_ (.D(_04100_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [155]),
    .QN(_00531_));
 DFF_X1 _65996_ (.D(_04101_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [156]),
    .QN(_00547_));
 DFF_X1 _65997_ (.D(_04102_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [157]),
    .QN(_00563_));
 DFF_X1 _65998_ (.D(_04103_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [158]),
    .QN(_32341_));
 DFF_X1 _65999_ (.D(_04104_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [159]),
    .QN(_32342_));
 DFF_X1 _66000_ (.D(_04106_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [160]),
    .QN(_00107_));
 DFF_X1 _66001_ (.D(_04107_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [161]),
    .QN(_00123_));
 DFF_X1 _66002_ (.D(_04108_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [162]),
    .QN(_00139_));
 DFF_X1 _66003_ (.D(_04109_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [163]),
    .QN(_00155_));
 DFF_X1 _66004_ (.D(_04110_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [164]),
    .QN(_00171_));
 DFF_X1 _66005_ (.D(_04111_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [165]),
    .QN(_00187_));
 DFF_X1 _66006_ (.D(_04112_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [166]),
    .QN(_00203_));
 DFF_X1 _66007_ (.D(_04113_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [167]),
    .QN(_00219_));
 DFF_X1 _66008_ (.D(_04114_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [168]),
    .QN(_00235_));
 DFF_X1 _66009_ (.D(_04115_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [169]),
    .QN(_00251_));
 DFF_X1 _66010_ (.D(_04117_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [170]),
    .QN(_00267_));
 DFF_X1 _66011_ (.D(_04118_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [171]),
    .QN(_00283_));
 DFF_X1 _66012_ (.D(_04119_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [172]),
    .QN(_00299_));
 DFF_X1 _66013_ (.D(_04120_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [173]),
    .QN(_00315_));
 DFF_X1 _66014_ (.D(_04121_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [174]),
    .QN(_00331_));
 DFF_X1 _66015_ (.D(_04122_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [175]),
    .QN(_00347_));
 DFF_X1 _66016_ (.D(_04123_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [176]),
    .QN(_00363_));
 DFF_X1 _66017_ (.D(_04124_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [177]),
    .QN(_00379_));
 DFF_X1 _66018_ (.D(_04125_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [178]),
    .QN(_00395_));
 DFF_X1 _66019_ (.D(_04126_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [179]),
    .QN(_00411_));
 DFF_X1 _66020_ (.D(_04128_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [180]),
    .QN(_00427_));
 DFF_X1 _66021_ (.D(_04129_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [181]),
    .QN(_00443_));
 DFF_X1 _66022_ (.D(_04130_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [182]),
    .QN(_00459_));
 DFF_X1 _66023_ (.D(_04131_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [183]),
    .QN(_00475_));
 DFF_X1 _66024_ (.D(_04132_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [184]),
    .QN(_00491_));
 DFF_X1 _66025_ (.D(_04133_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [185]),
    .QN(_00507_));
 DFF_X1 _66026_ (.D(_04134_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [186]),
    .QN(_00523_));
 DFF_X1 _66027_ (.D(_04135_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [187]),
    .QN(_00539_));
 DFF_X1 _66028_ (.D(_04136_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [188]),
    .QN(_00555_));
 DFF_X1 _66029_ (.D(_04137_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [189]),
    .QN(_00571_));
 DFF_X1 _66030_ (.D(_04139_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [190]),
    .QN(_32343_));
 DFF_X1 _66031_ (.D(_04140_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [191]),
    .QN(_32344_));
 DFF_X1 _66032_ (.D(_04141_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [192]),
    .QN(_00100_));
 DFF_X1 _66033_ (.D(_04142_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [193]),
    .QN(_00116_));
 DFF_X1 _66034_ (.D(_04143_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [194]),
    .QN(_00132_));
 DFF_X1 _66035_ (.D(_04144_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [195]),
    .QN(_00148_));
 DFF_X1 _66036_ (.D(_04145_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [196]),
    .QN(_00164_));
 DFF_X1 _66037_ (.D(_04146_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [197]),
    .QN(_00180_));
 DFF_X1 _66038_ (.D(_04147_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [198]),
    .QN(_00196_));
 DFF_X1 _66039_ (.D(_04148_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [199]),
    .QN(_00212_));
 DFF_X1 _66040_ (.D(_04151_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [200]),
    .QN(_00228_));
 DFF_X1 _66041_ (.D(_04152_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [201]),
    .QN(_00244_));
 DFF_X1 _66042_ (.D(_04153_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [202]),
    .QN(_00260_));
 DFF_X1 _66043_ (.D(_04154_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [203]),
    .QN(_00276_));
 DFF_X1 _66044_ (.D(_04155_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [204]),
    .QN(_00292_));
 DFF_X1 _66045_ (.D(_04156_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [205]),
    .QN(_00308_));
 DFF_X1 _66046_ (.D(_04157_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [206]),
    .QN(_00324_));
 DFF_X1 _66047_ (.D(_04158_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [207]),
    .QN(_00340_));
 DFF_X1 _66048_ (.D(_04159_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [208]),
    .QN(_00356_));
 DFF_X1 _66049_ (.D(_04160_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [209]),
    .QN(_00372_));
 DFF_X1 _66050_ (.D(_04162_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [210]),
    .QN(_00388_));
 DFF_X1 _66051_ (.D(_04163_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [211]),
    .QN(_00404_));
 DFF_X1 _66052_ (.D(_04164_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [212]),
    .QN(_00420_));
 DFF_X1 _66053_ (.D(_04165_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [213]),
    .QN(_00436_));
 DFF_X1 _66054_ (.D(_04166_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [214]),
    .QN(_00452_));
 DFF_X1 _66055_ (.D(_04167_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [215]),
    .QN(_00468_));
 DFF_X1 _66056_ (.D(_04168_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [216]),
    .QN(_00484_));
 DFF_X1 _66057_ (.D(_04169_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [217]),
    .QN(_00500_));
 DFF_X1 _66058_ (.D(_04170_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [218]),
    .QN(_00516_));
 DFF_X1 _66059_ (.D(_04171_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [219]),
    .QN(_00532_));
 DFF_X1 _66060_ (.D(_04173_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [220]),
    .QN(_00548_));
 DFF_X1 _66061_ (.D(_04174_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [221]),
    .QN(_00564_));
 DFF_X1 _66062_ (.D(_04175_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [222]),
    .QN(_32345_));
 DFF_X1 _66063_ (.D(_04176_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [223]),
    .QN(_32346_));
 DFF_X1 _66064_ (.D(_04177_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [224]),
    .QN(_00108_));
 DFF_X1 _66065_ (.D(_04178_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [225]),
    .QN(_00124_));
 DFF_X1 _66066_ (.D(_04179_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [226]),
    .QN(_00140_));
 DFF_X1 _66067_ (.D(_04180_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [227]),
    .QN(_00156_));
 DFF_X1 _66068_ (.D(_04181_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [228]),
    .QN(_00172_));
 DFF_X1 _66069_ (.D(_04182_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [229]),
    .QN(_00188_));
 DFF_X1 _66070_ (.D(_04184_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [230]),
    .QN(_00204_));
 DFF_X1 _66071_ (.D(_04185_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [231]),
    .QN(_00220_));
 DFF_X1 _66072_ (.D(_04186_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [232]),
    .QN(_00236_));
 DFF_X1 _66073_ (.D(_04187_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [233]),
    .QN(_00252_));
 DFF_X1 _66074_ (.D(_04188_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [234]),
    .QN(_00268_));
 DFF_X1 _66075_ (.D(_04189_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [235]),
    .QN(_00284_));
 DFF_X1 _66076_ (.D(_04190_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [236]),
    .QN(_00300_));
 DFF_X1 _66077_ (.D(_04191_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [237]),
    .QN(_00316_));
 DFF_X1 _66078_ (.D(_04192_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [238]),
    .QN(_00332_));
 DFF_X1 _66079_ (.D(_04193_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [239]),
    .QN(_00348_));
 DFF_X1 _66080_ (.D(_04195_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [240]),
    .QN(_00364_));
 DFF_X1 _66081_ (.D(_04196_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [241]),
    .QN(_00380_));
 DFF_X1 _66082_ (.D(_04197_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [242]),
    .QN(_00396_));
 DFF_X1 _66083_ (.D(_04198_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [243]),
    .QN(_00412_));
 DFF_X1 _66084_ (.D(_04199_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [244]),
    .QN(_00428_));
 DFF_X1 _66085_ (.D(_04200_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [245]),
    .QN(_00444_));
 DFF_X1 _66086_ (.D(_04201_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [246]),
    .QN(_00460_));
 DFF_X1 _66087_ (.D(_04202_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [247]),
    .QN(_00476_));
 DFF_X1 _66088_ (.D(_04203_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [248]),
    .QN(_00492_));
 DFF_X1 _66089_ (.D(_04204_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [249]),
    .QN(_00508_));
 DFF_X1 _66090_ (.D(_04206_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [250]),
    .QN(_00524_));
 DFF_X1 _66091_ (.D(_04207_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [251]),
    .QN(_00540_));
 DFF_X1 _66092_ (.D(_04208_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [252]),
    .QN(_00556_));
 DFF_X1 _66093_ (.D(_04209_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [253]),
    .QN(_00572_));
 DFF_X1 _66094_ (.D(_04210_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [254]),
    .QN(_32347_));
 DFF_X1 _66095_ (.D(_04211_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [255]),
    .QN(_32348_));
 DFF_X1 _66096_ (.D(_04212_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [256]),
    .QN(_00101_));
 DFF_X1 _66097_ (.D(_04213_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [257]),
    .QN(_00117_));
 DFF_X1 _66098_ (.D(_04214_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [258]),
    .QN(_00133_));
 DFF_X1 _66099_ (.D(_04215_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [259]),
    .QN(_00149_));
 DFF_X1 _66100_ (.D(_04217_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [260]),
    .QN(_00165_));
 DFF_X1 _66101_ (.D(_04218_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [261]),
    .QN(_00181_));
 DFF_X1 _66102_ (.D(_04219_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [262]),
    .QN(_00197_));
 DFF_X1 _66103_ (.D(_04220_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [263]),
    .QN(_00213_));
 DFF_X1 _66104_ (.D(_04221_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [264]),
    .QN(_00229_));
 DFF_X1 _66105_ (.D(_04222_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [265]),
    .QN(_00245_));
 DFF_X1 _66106_ (.D(_04223_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [266]),
    .QN(_00261_));
 DFF_X1 _66107_ (.D(_04224_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [267]),
    .QN(_00277_));
 DFF_X1 _66108_ (.D(_04225_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [268]),
    .QN(_00293_));
 DFF_X1 _66109_ (.D(_04226_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [269]),
    .QN(_00309_));
 DFF_X1 _66110_ (.D(_04228_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [270]),
    .QN(_00325_));
 DFF_X1 _66111_ (.D(_04229_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [271]),
    .QN(_00341_));
 DFF_X1 _66112_ (.D(_04230_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [272]),
    .QN(_00357_));
 DFF_X1 _66113_ (.D(_04231_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [273]),
    .QN(_00373_));
 DFF_X1 _66114_ (.D(_04232_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [274]),
    .QN(_00389_));
 DFF_X1 _66115_ (.D(_04233_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [275]),
    .QN(_00405_));
 DFF_X1 _66116_ (.D(_04234_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [276]),
    .QN(_00421_));
 DFF_X1 _66117_ (.D(_04235_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [277]),
    .QN(_00437_));
 DFF_X1 _66118_ (.D(_04236_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [278]),
    .QN(_00453_));
 DFF_X1 _66119_ (.D(_04237_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [279]),
    .QN(_00469_));
 DFF_X1 _66120_ (.D(_04239_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [280]),
    .QN(_00485_));
 DFF_X1 _66121_ (.D(_04240_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [281]),
    .QN(_00501_));
 DFF_X1 _66122_ (.D(_04241_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [282]),
    .QN(_00517_));
 DFF_X1 _66123_ (.D(_04242_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [283]),
    .QN(_00533_));
 DFF_X1 _66124_ (.D(_04243_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [284]),
    .QN(_00549_));
 DFF_X1 _66125_ (.D(_04244_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [285]),
    .QN(_00565_));
 DFF_X1 _66126_ (.D(_04245_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [286]),
    .QN(_32349_));
 DFF_X1 _66127_ (.D(_04246_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [287]),
    .QN(_32350_));
 DFF_X1 _66128_ (.D(_04247_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [288]),
    .QN(_00109_));
 DFF_X1 _66129_ (.D(_04248_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [289]),
    .QN(_00125_));
 DFF_X1 _66130_ (.D(_04250_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [290]),
    .QN(_00141_));
 DFF_X1 _66131_ (.D(_04251_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [291]),
    .QN(_00157_));
 DFF_X1 _66132_ (.D(_04252_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [292]),
    .QN(_00173_));
 DFF_X1 _66133_ (.D(_04253_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [293]),
    .QN(_00189_));
 DFF_X1 _66134_ (.D(_04254_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [294]),
    .QN(_00205_));
 DFF_X1 _66135_ (.D(_04255_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [295]),
    .QN(_00221_));
 DFF_X1 _66136_ (.D(_04256_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [296]),
    .QN(_00237_));
 DFF_X1 _66137_ (.D(_04257_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [297]),
    .QN(_00253_));
 DFF_X1 _66138_ (.D(_04258_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [298]),
    .QN(_00269_));
 DFF_X1 _66139_ (.D(_04259_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [299]),
    .QN(_00285_));
 DFF_X1 _66140_ (.D(_04262_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [300]),
    .QN(_00301_));
 DFF_X1 _66141_ (.D(_04263_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [301]),
    .QN(_00317_));
 DFF_X1 _66142_ (.D(_04264_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [302]),
    .QN(_00333_));
 DFF_X1 _66143_ (.D(_04265_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [303]),
    .QN(_00349_));
 DFF_X1 _66144_ (.D(_04266_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [304]),
    .QN(_00365_));
 DFF_X1 _66145_ (.D(_04267_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [305]),
    .QN(_00381_));
 DFF_X1 _66146_ (.D(_04268_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [306]),
    .QN(_00397_));
 DFF_X1 _66147_ (.D(_04269_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [307]),
    .QN(_00413_));
 DFF_X1 _66148_ (.D(_04270_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [308]),
    .QN(_00429_));
 DFF_X1 _66149_ (.D(_04271_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [309]),
    .QN(_00445_));
 DFF_X1 _66150_ (.D(_04273_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [310]),
    .QN(_00461_));
 DFF_X1 _66151_ (.D(_04274_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [311]),
    .QN(_00477_));
 DFF_X1 _66152_ (.D(_04275_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [312]),
    .QN(_00493_));
 DFF_X1 _66153_ (.D(_04276_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [313]),
    .QN(_00509_));
 DFF_X1 _66154_ (.D(_04277_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [314]),
    .QN(_00525_));
 DFF_X1 _66155_ (.D(_04278_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [315]),
    .QN(_00541_));
 DFF_X1 _66156_ (.D(_04279_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [316]),
    .QN(_00557_));
 DFF_X1 _66157_ (.D(_04280_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [317]),
    .QN(_00573_));
 DFF_X1 _66158_ (.D(_04281_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [318]),
    .QN(_32351_));
 DFF_X1 _66159_ (.D(_04282_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [319]),
    .QN(_32352_));
 DFF_X1 _66160_ (.D(_04284_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [320]),
    .QN(_00102_));
 DFF_X1 _66161_ (.D(_04285_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [321]),
    .QN(_00118_));
 DFF_X1 _66162_ (.D(_04286_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [322]),
    .QN(_00134_));
 DFF_X1 _66163_ (.D(_04287_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [323]),
    .QN(_00150_));
 DFF_X1 _66164_ (.D(_04288_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [324]),
    .QN(_00166_));
 DFF_X1 _66165_ (.D(_04289_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [325]),
    .QN(_00182_));
 DFF_X1 _66166_ (.D(_04290_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [326]),
    .QN(_00198_));
 DFF_X1 _66167_ (.D(_04291_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [327]),
    .QN(_00214_));
 DFF_X1 _66168_ (.D(_04292_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [328]),
    .QN(_00230_));
 DFF_X1 _66169_ (.D(_04293_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [329]),
    .QN(_00246_));
 DFF_X1 _66170_ (.D(_04295_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [330]),
    .QN(_00262_));
 DFF_X1 _66171_ (.D(_04296_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [331]),
    .QN(_00278_));
 DFF_X1 _66172_ (.D(_04297_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [332]),
    .QN(_00294_));
 DFF_X1 _66173_ (.D(_04298_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [333]),
    .QN(_00310_));
 DFF_X1 _66174_ (.D(_04299_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [334]),
    .QN(_00326_));
 DFF_X1 _66175_ (.D(_04300_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [335]),
    .QN(_00342_));
 DFF_X1 _66176_ (.D(_04301_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [336]),
    .QN(_00358_));
 DFF_X1 _66177_ (.D(_04302_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [337]),
    .QN(_00374_));
 DFF_X1 _66178_ (.D(_04303_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [338]),
    .QN(_00390_));
 DFF_X1 _66179_ (.D(_04304_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [339]),
    .QN(_00406_));
 DFF_X1 _66180_ (.D(_04306_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [340]),
    .QN(_00422_));
 DFF_X1 _66181_ (.D(_04307_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [341]),
    .QN(_00438_));
 DFF_X1 _66182_ (.D(_04308_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [342]),
    .QN(_00454_));
 DFF_X1 _66183_ (.D(_04309_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [343]),
    .QN(_00470_));
 DFF_X1 _66184_ (.D(_04310_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [344]),
    .QN(_00486_));
 DFF_X1 _66185_ (.D(_04311_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [345]),
    .QN(_00502_));
 DFF_X1 _66186_ (.D(_04312_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [346]),
    .QN(_00518_));
 DFF_X1 _66187_ (.D(_04313_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [347]),
    .QN(_00534_));
 DFF_X1 _66188_ (.D(_04314_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [348]),
    .QN(_00550_));
 DFF_X1 _66189_ (.D(_04315_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [349]),
    .QN(_00566_));
 DFF_X1 _66190_ (.D(_04317_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [350]),
    .QN(_32353_));
 DFF_X1 _66191_ (.D(_04318_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [351]),
    .QN(_32354_));
 DFF_X1 _66192_ (.D(_04319_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [352]),
    .QN(_00110_));
 DFF_X1 _66193_ (.D(_04320_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [353]),
    .QN(_00126_));
 DFF_X1 _66194_ (.D(_04321_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [354]),
    .QN(_00142_));
 DFF_X1 _66195_ (.D(_04322_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [355]),
    .QN(_00158_));
 DFF_X1 _66196_ (.D(_04323_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [356]),
    .QN(_00174_));
 DFF_X1 _66197_ (.D(_04324_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [357]),
    .QN(_00190_));
 DFF_X1 _66198_ (.D(_04325_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [358]),
    .QN(_00206_));
 DFF_X1 _66199_ (.D(_04326_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [359]),
    .QN(_00222_));
 DFF_X1 _66200_ (.D(_04328_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [360]),
    .QN(_00238_));
 DFF_X1 _66201_ (.D(_04329_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [361]),
    .QN(_00254_));
 DFF_X1 _66202_ (.D(_04330_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [362]),
    .QN(_00270_));
 DFF_X1 _66203_ (.D(_04331_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [363]),
    .QN(_00286_));
 DFF_X1 _66204_ (.D(_04332_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [364]),
    .QN(_00302_));
 DFF_X1 _66205_ (.D(_04333_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [365]),
    .QN(_00318_));
 DFF_X1 _66206_ (.D(_04334_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [366]),
    .QN(_00334_));
 DFF_X1 _66207_ (.D(_04335_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [367]),
    .QN(_00350_));
 DFF_X1 _66208_ (.D(_04336_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [368]),
    .QN(_00366_));
 DFF_X1 _66209_ (.D(_04337_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [369]),
    .QN(_00382_));
 DFF_X1 _66210_ (.D(_04339_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [370]),
    .QN(_00398_));
 DFF_X1 _66211_ (.D(_04340_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [371]),
    .QN(_00414_));
 DFF_X1 _66212_ (.D(_04341_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [372]),
    .QN(_00430_));
 DFF_X1 _66213_ (.D(_04342_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [373]),
    .QN(_00446_));
 DFF_X1 _66214_ (.D(_04343_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [374]),
    .QN(_00462_));
 DFF_X1 _66215_ (.D(_04344_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [375]),
    .QN(_00478_));
 DFF_X1 _66216_ (.D(_04345_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [376]),
    .QN(_00494_));
 DFF_X1 _66217_ (.D(_04346_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [377]),
    .QN(_00510_));
 DFF_X1 _66218_ (.D(_04347_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [378]),
    .QN(_00526_));
 DFF_X1 _66219_ (.D(_04348_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [379]),
    .QN(_00542_));
 DFF_X1 _66220_ (.D(_04350_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [380]),
    .QN(_00558_));
 DFF_X1 _66221_ (.D(_04351_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [381]),
    .QN(_00574_));
 DFF_X1 _66222_ (.D(_04352_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [382]),
    .QN(_32355_));
 DFF_X1 _66223_ (.D(_04353_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [383]),
    .QN(_32356_));
 DFF_X1 _66224_ (.D(_04354_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [384]),
    .QN(_00103_));
 DFF_X1 _66225_ (.D(_04355_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [385]),
    .QN(_00119_));
 DFF_X1 _66226_ (.D(_04356_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [386]),
    .QN(_00135_));
 DFF_X1 _66227_ (.D(_04357_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [387]),
    .QN(_00151_));
 DFF_X1 _66228_ (.D(_04358_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [388]),
    .QN(_00167_));
 DFF_X1 _66229_ (.D(_04359_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [389]),
    .QN(_00183_));
 DFF_X1 _66230_ (.D(_04361_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [390]),
    .QN(_00199_));
 DFF_X1 _66231_ (.D(_04362_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [391]),
    .QN(_00215_));
 DFF_X1 _66232_ (.D(_04363_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [392]),
    .QN(_00231_));
 DFF_X1 _66233_ (.D(_04364_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [393]),
    .QN(_00247_));
 DFF_X1 _66234_ (.D(_04365_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [394]),
    .QN(_00263_));
 DFF_X1 _66235_ (.D(_04366_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [395]),
    .QN(_00279_));
 DFF_X1 _66236_ (.D(_04367_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [396]),
    .QN(_00295_));
 DFF_X1 _66237_ (.D(_04368_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [397]),
    .QN(_00311_));
 DFF_X1 _66238_ (.D(_04369_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [398]),
    .QN(_00327_));
 DFF_X1 _66239_ (.D(_04370_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [399]),
    .QN(_00343_));
 DFF_X1 _66240_ (.D(_04373_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [400]),
    .QN(_00359_));
 DFF_X1 _66241_ (.D(_04374_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [401]),
    .QN(_00375_));
 DFF_X1 _66242_ (.D(_04375_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [402]),
    .QN(_00391_));
 DFF_X1 _66243_ (.D(_04376_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [403]),
    .QN(_00407_));
 DFF_X1 _66244_ (.D(_04377_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [404]),
    .QN(_00423_));
 DFF_X1 _66245_ (.D(_04378_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [405]),
    .QN(_00439_));
 DFF_X1 _66246_ (.D(_04379_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [406]),
    .QN(_00455_));
 DFF_X1 _66247_ (.D(_04380_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [407]),
    .QN(_00471_));
 DFF_X1 _66248_ (.D(_04381_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [408]),
    .QN(_00487_));
 DFF_X1 _66249_ (.D(_04382_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [409]),
    .QN(_00503_));
 DFF_X1 _66250_ (.D(_04384_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [410]),
    .QN(_00519_));
 DFF_X1 _66251_ (.D(_04385_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [411]),
    .QN(_00535_));
 DFF_X1 _66252_ (.D(_04386_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [412]),
    .QN(_00551_));
 DFF_X1 _66253_ (.D(_04387_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [413]),
    .QN(_00567_));
 DFF_X1 _66254_ (.D(_04388_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [414]),
    .QN(_32357_));
 DFF_X1 _66255_ (.D(_04389_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [415]),
    .QN(_32358_));
 DFF_X1 _66256_ (.D(_04390_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [416]),
    .QN(_00111_));
 DFF_X1 _66257_ (.D(_04391_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [417]),
    .QN(_00127_));
 DFF_X1 _66258_ (.D(_04392_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [418]),
    .QN(_00143_));
 DFF_X1 _66259_ (.D(_04393_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [419]),
    .QN(_00159_));
 DFF_X1 _66260_ (.D(_04395_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [420]),
    .QN(_00175_));
 DFF_X1 _66261_ (.D(_04396_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [421]),
    .QN(_00191_));
 DFF_X1 _66262_ (.D(_04397_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [422]),
    .QN(_00207_));
 DFF_X1 _66263_ (.D(_04398_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [423]),
    .QN(_00223_));
 DFF_X1 _66264_ (.D(_04399_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [424]),
    .QN(_00239_));
 DFF_X1 _66265_ (.D(_04400_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [425]),
    .QN(_00255_));
 DFF_X1 _66266_ (.D(_04401_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [426]),
    .QN(_00271_));
 DFF_X1 _66267_ (.D(_04402_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [427]),
    .QN(_00287_));
 DFF_X1 _66268_ (.D(_04403_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [428]),
    .QN(_00303_));
 DFF_X1 _66269_ (.D(_04404_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [429]),
    .QN(_00319_));
 DFF_X1 _66270_ (.D(_04406_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [430]),
    .QN(_00335_));
 DFF_X1 _66271_ (.D(_04407_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [431]),
    .QN(_00351_));
 DFF_X1 _66272_ (.D(_04408_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [432]),
    .QN(_00367_));
 DFF_X1 _66273_ (.D(_04409_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [433]),
    .QN(_00383_));
 DFF_X1 _66274_ (.D(_04410_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [434]),
    .QN(_00399_));
 DFF_X1 _66275_ (.D(_04411_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [435]),
    .QN(_00415_));
 DFF_X1 _66276_ (.D(_04412_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [436]),
    .QN(_00431_));
 DFF_X1 _66277_ (.D(_04413_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [437]),
    .QN(_00447_));
 DFF_X1 _66278_ (.D(_04414_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [438]),
    .QN(_00463_));
 DFF_X1 _66279_ (.D(_04415_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [439]),
    .QN(_00479_));
 DFF_X1 _66280_ (.D(_04417_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [440]),
    .QN(_00495_));
 DFF_X1 _66281_ (.D(_04418_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [441]),
    .QN(_00511_));
 DFF_X1 _66282_ (.D(_04419_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [442]),
    .QN(_00527_));
 DFF_X1 _66283_ (.D(_04420_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [443]),
    .QN(_00543_));
 DFF_X1 _66284_ (.D(_04421_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [444]),
    .QN(_00559_));
 DFF_X1 _66285_ (.D(_04422_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [445]),
    .QN(_00575_));
 DFF_X1 _66286_ (.D(_04423_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [446]),
    .QN(_32359_));
 DFF_X1 _66287_ (.D(_04424_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [447]),
    .QN(_32360_));
 DFF_X1 _66288_ (.D(_04425_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [448]),
    .QN(_32361_));
 DFF_X1 _66289_ (.D(_04426_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [449]),
    .QN(_32362_));
 DFF_X1 _66290_ (.D(_04428_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [450]),
    .QN(_32363_));
 DFF_X1 _66291_ (.D(_04429_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [451]),
    .QN(_32364_));
 DFF_X1 _66292_ (.D(_04430_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [452]),
    .QN(_32365_));
 DFF_X1 _66293_ (.D(_04431_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [453]),
    .QN(_32366_));
 DFF_X1 _66294_ (.D(_04432_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [454]),
    .QN(_32367_));
 DFF_X1 _66295_ (.D(_04433_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [455]),
    .QN(_32368_));
 DFF_X1 _66296_ (.D(_04434_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [456]),
    .QN(_32369_));
 DFF_X1 _66297_ (.D(_04435_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [457]),
    .QN(_32370_));
 DFF_X1 _66298_ (.D(_04436_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [458]),
    .QN(_32371_));
 DFF_X1 _66299_ (.D(_04437_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [459]),
    .QN(_32372_));
 DFF_X1 _66300_ (.D(_04439_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [460]),
    .QN(_32373_));
 DFF_X1 _66301_ (.D(_04440_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [461]),
    .QN(_32374_));
 DFF_X1 _66302_ (.D(_04441_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [462]),
    .QN(_32375_));
 DFF_X1 _66303_ (.D(_04442_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [463]),
    .QN(_32376_));
 DFF_X1 _66304_ (.D(_04443_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [464]),
    .QN(_32377_));
 DFF_X1 _66305_ (.D(_04444_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [465]),
    .QN(_32378_));
 DFF_X1 _66306_ (.D(_04445_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [466]),
    .QN(_32379_));
 DFF_X1 _66307_ (.D(_04446_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [467]),
    .QN(_32380_));
 DFF_X1 _66308_ (.D(_04447_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [468]),
    .QN(_32381_));
 DFF_X1 _66309_ (.D(_04448_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [469]),
    .QN(_32382_));
 DFF_X1 _66310_ (.D(_04450_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [470]),
    .QN(_32383_));
 DFF_X1 _66311_ (.D(_04451_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [471]),
    .QN(_32384_));
 DFF_X1 _66312_ (.D(_04452_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [472]),
    .QN(_32385_));
 DFF_X1 _66313_ (.D(_04453_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [473]),
    .QN(_32386_));
 DFF_X1 _66314_ (.D(_04454_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [474]),
    .QN(_32387_));
 DFF_X1 _66315_ (.D(_04455_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [475]),
    .QN(_32388_));
 DFF_X1 _66316_ (.D(_04456_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [476]),
    .QN(_32389_));
 DFF_X1 _66317_ (.D(_04457_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [477]),
    .QN(_32390_));
 DFF_X1 _66318_ (.D(_04458_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [478]),
    .QN(_32391_));
 DFF_X1 _66319_ (.D(_04459_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [479]),
    .QN(_32392_));
 DFF_X1 _66320_ (.D(_04461_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [480]),
    .QN(_32393_));
 DFF_X1 _66321_ (.D(_04462_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [481]),
    .QN(_32394_));
 DFF_X1 _66322_ (.D(_04463_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [482]),
    .QN(_32395_));
 DFF_X1 _66323_ (.D(_04464_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [483]),
    .QN(_32396_));
 DFF_X1 _66324_ (.D(_04465_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [484]),
    .QN(_32397_));
 DFF_X1 _66325_ (.D(_04466_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [485]),
    .QN(_32398_));
 DFF_X1 _66326_ (.D(_04467_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [486]),
    .QN(_32399_));
 DFF_X1 _66327_ (.D(_04468_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [487]),
    .QN(_32400_));
 DFF_X1 _66328_ (.D(_04469_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [488]),
    .QN(_32401_));
 DFF_X1 _66329_ (.D(_04470_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [489]),
    .QN(_32402_));
 DFF_X1 _66330_ (.D(_04472_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [490]),
    .QN(_32403_));
 DFF_X1 _66331_ (.D(_04473_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [491]),
    .QN(_32404_));
 DFF_X1 _66332_ (.D(_04474_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [492]),
    .QN(_32405_));
 DFF_X1 _66333_ (.D(_04475_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [493]),
    .QN(_32406_));
 DFF_X1 _66334_ (.D(_04476_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [494]),
    .QN(_32407_));
 DFF_X1 _66335_ (.D(_04477_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [495]),
    .QN(_32408_));
 DFF_X1 _66336_ (.D(_04478_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [496]),
    .QN(_32409_));
 DFF_X1 _66337_ (.D(_04479_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [497]),
    .QN(_32410_));
 DFF_X1 _66338_ (.D(_04480_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [498]),
    .QN(_32411_));
 DFF_X1 _66339_ (.D(_04481_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [499]),
    .QN(_32412_));
 DFF_X1 _66340_ (.D(_04484_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [500]),
    .QN(_32413_));
 DFF_X1 _66341_ (.D(_04485_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [501]),
    .QN(_32414_));
 DFF_X1 _66342_ (.D(_04486_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [502]),
    .QN(_32415_));
 DFF_X1 _66343_ (.D(_04487_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [503]),
    .QN(_32416_));
 DFF_X1 _66344_ (.D(_04488_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [504]),
    .QN(_32417_));
 DFF_X1 _66345_ (.D(_04489_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [505]),
    .QN(_32418_));
 DFF_X1 _66346_ (.D(_04490_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [506]),
    .QN(_32419_));
 DFF_X1 _66347_ (.D(_04491_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [507]),
    .QN(_32420_));
 DFF_X1 _66348_ (.D(_04492_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [508]),
    .QN(_32421_));
 DFF_X1 _66349_ (.D(_04493_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [509]),
    .QN(_32422_));
 DFF_X1 _66350_ (.D(_04495_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [510]),
    .QN(_32423_));
 DFF_X1 _66351_ (.D(_04496_),
    .CK(clk_i),
    .Q(\icache.data_set_select_mux.data_i [511]),
    .QN(_32424_));
 DFF_X1 _66352_ (.D(_04847_),
    .CK(clk_i),
    .Q(\icache.final_data_mux.N0 ),
    .QN(_00003_));
 DFF_X1 _66353_ (.D(_04848_),
    .CK(clk_i),
    .Q(\icache.N8 ),
    .QN(_32425_));
 DFF_X1 _66354_ (.D(\icache.N29 ),
    .CK(clk_i),
    .Q(\icache.N10 ),
    .QN(_00000_));
 DFF_X1 _66355_ (.D(_04849_),
    .CK(clk_i),
    .Q(\icache.vaddr_tl_r [0]),
    .QN(_32426_));
 DFF_X1 _66356_ (.D(_04860_),
    .CK(clk_i),
    .Q(\icache.vaddr_tl_r [1]),
    .QN(_32427_));
 DFF_X1 _66357_ (.D(_04871_),
    .CK(clk_i),
    .Q(\icache.vaddr_tl_r [2]),
    .QN(_32428_));
 DFF_X1 _66358_ (.D(_04881_),
    .CK(clk_i),
    .Q(\icache.vaddr_tl_r [3]),
    .QN(_32429_));
 DFF_X1 _66359_ (.D(_04882_),
    .CK(clk_i),
    .Q(\icache.vaddr_tl_r [4]),
    .QN(_32430_));
 DFF_X1 _66360_ (.D(_04883_),
    .CK(clk_i),
    .Q(\icache.vaddr_tl_r [5]),
    .QN(_32431_));
 DFF_X1 _66361_ (.D(_04884_),
    .CK(clk_i),
    .Q(\icache.vaddr_tl_r [6]),
    .QN(_32432_));
 DFF_X1 _66362_ (.D(_04885_),
    .CK(clk_i),
    .Q(\icache.vaddr_tl_r [7]),
    .QN(_32433_));
 DFF_X1 _66363_ (.D(_04886_),
    .CK(clk_i),
    .Q(\icache.vaddr_tl_r [8]),
    .QN(_32434_));
 DFF_X1 _66364_ (.D(_04887_),
    .CK(clk_i),
    .Q(\icache.vaddr_tl_r [9]),
    .QN(_32435_));
 DFF_X1 _66365_ (.D(_04850_),
    .CK(clk_i),
    .Q(\icache.vaddr_tl_r [10]),
    .QN(_32436_));
 DFF_X1 _66366_ (.D(_04851_),
    .CK(clk_i),
    .Q(\icache.vaddr_tl_r [11]),
    .QN(_32437_));
 DFF_X1 _66367_ (.D(_04852_),
    .CK(clk_i),
    .Q(\icache.vaddr_tl_r [12]),
    .QN(_32438_));
 DFF_X1 _66368_ (.D(_04853_),
    .CK(clk_i),
    .Q(\icache.vaddr_tl_r [13]),
    .QN(_32439_));
 DFF_X1 _66369_ (.D(_04854_),
    .CK(clk_i),
    .Q(\icache.vaddr_tl_r [14]),
    .QN(_32440_));
 DFF_X1 _66370_ (.D(_04855_),
    .CK(clk_i),
    .Q(\icache.vaddr_tl_r [15]),
    .QN(_32441_));
 DFF_X1 _66371_ (.D(_04856_),
    .CK(clk_i),
    .Q(\icache.vaddr_tl_r [16]),
    .QN(_32442_));
 DFF_X1 _66372_ (.D(_04857_),
    .CK(clk_i),
    .Q(\icache.vaddr_tl_r [17]),
    .QN(_32443_));
 DFF_X1 _66373_ (.D(_04858_),
    .CK(clk_i),
    .Q(\icache.vaddr_tl_r [18]),
    .QN(_32444_));
 DFF_X1 _66374_ (.D(_04859_),
    .CK(clk_i),
    .Q(\icache.vaddr_tl_r [19]),
    .QN(_32445_));
 DFF_X1 _66375_ (.D(_04861_),
    .CK(clk_i),
    .Q(\icache.vaddr_tl_r [20]),
    .QN(_32446_));
 DFF_X1 _66376_ (.D(_04862_),
    .CK(clk_i),
    .Q(\icache.vaddr_tl_r [21]),
    .QN(_32447_));
 DFF_X1 _66377_ (.D(_04863_),
    .CK(clk_i),
    .Q(\icache.vaddr_tl_r [22]),
    .QN(_32448_));
 DFF_X1 _66378_ (.D(_04864_),
    .CK(clk_i),
    .Q(\icache.vaddr_tl_r [23]),
    .QN(_32449_));
 DFF_X1 _66379_ (.D(_04865_),
    .CK(clk_i),
    .Q(\icache.vaddr_tl_r [24]),
    .QN(_32450_));
 DFF_X1 _66380_ (.D(_04866_),
    .CK(clk_i),
    .Q(\icache.vaddr_tl_r [25]),
    .QN(_32451_));
 DFF_X1 _66381_ (.D(_04867_),
    .CK(clk_i),
    .Q(\icache.vaddr_tl_r [26]),
    .QN(_32452_));
 DFF_X1 _66382_ (.D(_04868_),
    .CK(clk_i),
    .Q(\icache.vaddr_tl_r [27]),
    .QN(_32453_));
 DFF_X1 _66383_ (.D(_04869_),
    .CK(clk_i),
    .Q(\icache.vaddr_tl_r [28]),
    .QN(_32454_));
 DFF_X1 _66384_ (.D(_04870_),
    .CK(clk_i),
    .Q(\icache.vaddr_tl_r [29]),
    .QN(_32455_));
 DFF_X1 _66385_ (.D(_04872_),
    .CK(clk_i),
    .Q(\icache.vaddr_tl_r [30]),
    .QN(_32456_));
 DFF_X1 _66386_ (.D(_04873_),
    .CK(clk_i),
    .Q(\icache.vaddr_tl_r [31]),
    .QN(_32457_));
 DFF_X1 _66387_ (.D(_04874_),
    .CK(clk_i),
    .Q(\icache.vaddr_tl_r [32]),
    .QN(_32458_));
 DFF_X1 _66388_ (.D(_04875_),
    .CK(clk_i),
    .Q(\icache.vaddr_tl_r [33]),
    .QN(_32459_));
 DFF_X1 _66389_ (.D(_04876_),
    .CK(clk_i),
    .Q(\icache.vaddr_tl_r [34]),
    .QN(_32460_));
 DFF_X1 _66390_ (.D(_04877_),
    .CK(clk_i),
    .Q(\icache.vaddr_tl_r [35]),
    .QN(_32461_));
 DFF_X1 _66391_ (.D(_04878_),
    .CK(clk_i),
    .Q(\icache.vaddr_tl_r [36]),
    .QN(_32462_));
 DFF_X1 _66392_ (.D(_04879_),
    .CK(clk_i),
    .Q(\icache.vaddr_tl_r [37]),
    .QN(_32463_));
 DFF_X1 _66393_ (.D(_04880_),
    .CK(clk_i),
    .Q(\icache.vaddr_tl_r [38]),
    .QN(_32464_));
 DFF_X1 _66394_ (.D(\icache.N25 ),
    .CK(clk_i),
    .Q(\icache.itlb_icache_data_resp_ready_o ),
    .QN(_32465_));
 DFF_X1 _66395_ (.D(_03997_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.icache_pc_gen_i [0]),
    .QN(_32466_));
 DFF_X1 _66396_ (.D(_04008_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.icache_pc_gen_i [1]),
    .QN(_32467_));
 DFF_X1 _66397_ (.D(_04019_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [11]),
    .QN(_32468_));
 DFF_X1 _66398_ (.D(_04029_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [12]),
    .QN(_32469_));
 DFF_X1 _66399_ (.D(_04030_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [13]),
    .QN(_32470_));
 DFF_X1 _66400_ (.D(_04031_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [14]),
    .QN(_32471_));
 DFF_X1 _66401_ (.D(_04032_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [15]),
    .QN(_32472_));
 DFF_X1 _66402_ (.D(_04033_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [16]),
    .QN(_32473_));
 DFF_X1 _66403_ (.D(_04034_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [17]),
    .QN(_32474_));
 DFF_X1 _66404_ (.D(_04035_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [18]),
    .QN(_32475_));
 DFF_X1 _66405_ (.D(_03998_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [19]),
    .QN(_32476_));
 DFF_X1 _66406_ (.D(_03999_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [20]),
    .QN(_32477_));
 DFF_X1 _66407_ (.D(_04000_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [21]),
    .QN(_32478_));
 DFF_X1 _66408_ (.D(_04001_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [22]),
    .QN(_32479_));
 DFF_X1 _66409_ (.D(_04002_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [23]),
    .QN(_32480_));
 DFF_X1 _66410_ (.D(_04003_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [24]),
    .QN(_32481_));
 DFF_X1 _66411_ (.D(_04004_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [25]),
    .QN(_32482_));
 DFF_X1 _66412_ (.D(_04005_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.branch_metadata_fwd_reg.data_i [26]),
    .QN(_32483_));
 DFF_X1 _66413_ (.D(_04006_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.icache_pc_gen_i [18]),
    .QN(_32484_));
 DFF_X1 _66414_ (.D(_04007_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.icache_pc_gen_i [19]),
    .QN(_32485_));
 DFF_X1 _66415_ (.D(_04009_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.icache_pc_gen_i [20]),
    .QN(_32486_));
 DFF_X1 _66416_ (.D(_04010_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.icache_pc_gen_i [21]),
    .QN(_32487_));
 DFF_X1 _66417_ (.D(_04011_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.icache_pc_gen_i [22]),
    .QN(_32488_));
 DFF_X1 _66418_ (.D(_04012_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.icache_pc_gen_i [23]),
    .QN(_32489_));
 DFF_X1 _66419_ (.D(_04013_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.icache_pc_gen_i [24]),
    .QN(_32490_));
 DFF_X1 _66420_ (.D(_04014_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.icache_pc_gen_i [25]),
    .QN(_32491_));
 DFF_X1 _66421_ (.D(_04015_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.icache_pc_gen_i [26]),
    .QN(_32492_));
 DFF_X1 _66422_ (.D(_04016_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.icache_pc_gen_i [27]),
    .QN(_32493_));
 DFF_X1 _66423_ (.D(_04017_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.icache_pc_gen_i [28]),
    .QN(_32494_));
 DFF_X1 _66424_ (.D(_04018_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.icache_pc_gen_i [29]),
    .QN(_32495_));
 DFF_X1 _66425_ (.D(_04020_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.icache_pc_gen_i [30]),
    .QN(_32496_));
 DFF_X1 _66426_ (.D(_04021_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.icache_pc_gen_i [31]),
    .QN(_32497_));
 DFF_X1 _66427_ (.D(_04022_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.icache_pc_gen_i [32]),
    .QN(_32498_));
 DFF_X1 _66428_ (.D(_04023_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.icache_pc_gen_i [33]),
    .QN(_32499_));
 DFF_X1 _66429_ (.D(_04024_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.icache_pc_gen_i [34]),
    .QN(_32500_));
 DFF_X1 _66430_ (.D(_04025_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.icache_pc_gen_i [35]),
    .QN(_32501_));
 DFF_X1 _66431_ (.D(_04026_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.icache_pc_gen_i [36]),
    .QN(_32502_));
 DFF_X1 _66432_ (.D(_04027_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.icache_pc_gen_i [37]),
    .QN(_32503_));
 DFF_X1 _66433_ (.D(_04028_),
    .CK(clk_i),
    .Q(\bp_fe_pc_gen_1.icache_pc_gen_i [38]),
    .QN(_32504_));
 BUF_X4 buffer1 (.A(_26016_),
    .Z(net1));
 BUF_X4 buffer10 (.A(_24775_),
    .Z(net10));
 BUF_X4 buffer100 (.A(net97),
    .Z(net100));
 BUF_X4 buffer1000 (.A(\icache.stat_mem.data_i [6]),
    .Z(net1000));
 BUF_X4 buffer1001 (.A(\icache.stat_mem.w_mask_i [5]),
    .Z(net1001));
 BUF_X4 buffer1002 (.A(net1001),
    .Z(net1002));
 BUF_X4 buffer1003 (.A(\icache.n_9_net_ ),
    .Z(net1003));
 BUF_X4 buffer1004 (.A(\icache.stat_mem.data_i [4]),
    .Z(net1004));
 BUF_X4 buffer1005 (.A(\icache.tag_mem.data_i [103]),
    .Z(net1005));
 BUF_X4 buffer1006 (.A(\icache.tag_mem.data_i [103]),
    .Z(net1006));
 BUF_X4 buffer1007 (.A(\icache.tag_mem.data_i [103]),
    .Z(net1007));
 BUF_X4 buffer1008 (.A(\icache.tag_mem.data_i [103]),
    .Z(net1008));
 BUF_X4 buffer1009 (.A(\icache.tag_mem.data_i [103]),
    .Z(net1009));
 BUF_X4 buffer101 (.A(net97),
    .Z(net101));
 BUF_X4 buffer1010 (.A(\icache.tag_mem.data_i [103]),
    .Z(net1010));
 BUF_X4 buffer1011 (.A(\icache.tag_mem.data_i [103]),
    .Z(net1011));
 BUF_X4 buffer1012 (.A(\icache.tag_mem.data_i [103]),
    .Z(net1012));
 BUF_X4 buffer1013 (.A(\icache.tag_mem.data_i [102]),
    .Z(net1013));
 BUF_X4 buffer1014 (.A(\icache.tag_mem.data_i [102]),
    .Z(net1014));
 BUF_X4 buffer1015 (.A(\icache.tag_mem.data_i [102]),
    .Z(net1015));
 BUF_X4 buffer1016 (.A(\icache.tag_mem.data_i [102]),
    .Z(net1016));
 BUF_X4 buffer1017 (.A(\icache.tag_mem.data_i [102]),
    .Z(net1017));
 BUF_X4 buffer1018 (.A(\icache.tag_mem.data_i [102]),
    .Z(net1018));
 BUF_X4 buffer1019 (.A(\icache.tag_mem.data_i [102]),
    .Z(net1019));
 BUF_X4 buffer102 (.A(net101),
    .Z(net102));
 BUF_X4 buffer1020 (.A(\icache.tag_mem.data_i [102]),
    .Z(net1020));
 BUF_X4 buffer1021 (.A(\icache.tag_mem.data_i [128]),
    .Z(net1021));
 BUF_X4 buffer1022 (.A(\icache.tag_mem.data_i [128]),
    .Z(net1022));
 BUF_X4 buffer1023 (.A(\icache.tag_mem.data_i [128]),
    .Z(net1023));
 BUF_X4 buffer1024 (.A(\icache.tag_mem.data_i [128]),
    .Z(net1024));
 BUF_X4 buffer1025 (.A(\icache.tag_mem.data_i [128]),
    .Z(net1025));
 BUF_X4 buffer1026 (.A(\icache.tag_mem.data_i [128]),
    .Z(net1026));
 BUF_X4 buffer1027 (.A(\icache.tag_mem.data_i [128]),
    .Z(net1027));
 BUF_X4 buffer1028 (.A(\icache.tag_mem.data_i [128]),
    .Z(net1028));
 BUF_X4 buffer1029 (.A(\icache.tag_mem.data_i [11]),
    .Z(net1029));
 BUF_X4 buffer103 (.A(net101),
    .Z(net103));
 BUF_X4 buffer1030 (.A(\icache.tag_mem.data_i [11]),
    .Z(net1030));
 BUF_X4 buffer1031 (.A(\icache.tag_mem.data_i [11]),
    .Z(net1031));
 BUF_X4 buffer1032 (.A(\icache.tag_mem.data_i [11]),
    .Z(net1032));
 BUF_X4 buffer1033 (.A(\icache.tag_mem.data_i [11]),
    .Z(net1033));
 BUF_X4 buffer1034 (.A(\icache.tag_mem.data_i [11]),
    .Z(net1034));
 BUF_X4 buffer1035 (.A(\icache.tag_mem.data_i [11]),
    .Z(net1035));
 BUF_X4 buffer1036 (.A(\icache.tag_mem.data_i [11]),
    .Z(net1036));
 BUF_X4 buffer1037 (.A(\icache.tag_mem.data_i [125]),
    .Z(net1037));
 BUF_X4 buffer1038 (.A(\icache.tag_mem.data_i [125]),
    .Z(net1038));
 BUF_X4 buffer1039 (.A(\icache.tag_mem.data_i [125]),
    .Z(net1039));
 BUF_X4 buffer104 (.A(_10772_),
    .Z(net104));
 BUF_X4 buffer1040 (.A(\icache.tag_mem.data_i [125]),
    .Z(net1040));
 BUF_X4 buffer1041 (.A(\icache.tag_mem.data_i [125]),
    .Z(net1041));
 BUF_X4 buffer1042 (.A(\icache.tag_mem.data_i [125]),
    .Z(net1042));
 BUF_X4 buffer1043 (.A(\icache.tag_mem.data_i [125]),
    .Z(net1043));
 BUF_X4 buffer1044 (.A(\icache.tag_mem.data_i [125]),
    .Z(net1044));
 BUF_X4 buffer1045 (.A(\icache.tag_mem.data_i [124]),
    .Z(net1045));
 BUF_X4 buffer1046 (.A(\icache.tag_mem.data_i [124]),
    .Z(net1046));
 BUF_X4 buffer1047 (.A(\icache.tag_mem.data_i [124]),
    .Z(net1047));
 BUF_X4 buffer1048 (.A(\icache.tag_mem.data_i [124]),
    .Z(net1048));
 BUF_X4 buffer1049 (.A(\icache.tag_mem.data_i [124]),
    .Z(net1049));
 BUF_X4 buffer105 (.A(net104),
    .Z(net105));
 BUF_X4 buffer1050 (.A(\icache.tag_mem.data_i [124]),
    .Z(net1050));
 BUF_X4 buffer1051 (.A(\icache.tag_mem.data_i [124]),
    .Z(net1051));
 BUF_X4 buffer1052 (.A(\icache.tag_mem.data_i [124]),
    .Z(net1052));
 BUF_X4 buffer1053 (.A(\icache.tag_mem.data_i [121]),
    .Z(net1053));
 BUF_X4 buffer1054 (.A(\icache.tag_mem.data_i [121]),
    .Z(net1054));
 BUF_X4 buffer1055 (.A(\icache.tag_mem.data_i [121]),
    .Z(net1055));
 BUF_X4 buffer1056 (.A(\icache.tag_mem.data_i [121]),
    .Z(net1056));
 BUF_X4 buffer1057 (.A(\icache.tag_mem.data_i [121]),
    .Z(net1057));
 BUF_X4 buffer1058 (.A(\icache.tag_mem.data_i [121]),
    .Z(net1058));
 BUF_X4 buffer1059 (.A(\icache.tag_mem.data_i [121]),
    .Z(net1059));
 BUF_X4 buffer106 (.A(net104),
    .Z(net106));
 BUF_X4 buffer1060 (.A(\icache.tag_mem.data_i [121]),
    .Z(net1060));
 BUF_X4 buffer1061 (.A(\icache.tag_mem.data_i [120]),
    .Z(net1061));
 BUF_X4 buffer1062 (.A(\icache.tag_mem.data_i [120]),
    .Z(net1062));
 BUF_X4 buffer1063 (.A(\icache.tag_mem.data_i [120]),
    .Z(net1063));
 BUF_X4 buffer1064 (.A(\icache.tag_mem.data_i [120]),
    .Z(net1064));
 BUF_X4 buffer1065 (.A(\icache.tag_mem.data_i [120]),
    .Z(net1065));
 BUF_X4 buffer1066 (.A(\icache.tag_mem.data_i [120]),
    .Z(net1066));
 BUF_X4 buffer1067 (.A(\icache.tag_mem.data_i [120]),
    .Z(net1067));
 BUF_X4 buffer1068 (.A(\icache.tag_mem.data_i [120]),
    .Z(net1068));
 BUF_X4 buffer1069 (.A(\icache.tag_mem.data_i [119]),
    .Z(net1069));
 BUF_X4 buffer107 (.A(net104),
    .Z(net107));
 BUF_X4 buffer1070 (.A(\icache.tag_mem.data_i [119]),
    .Z(net1070));
 BUF_X4 buffer1071 (.A(\icache.tag_mem.data_i [119]),
    .Z(net1071));
 BUF_X4 buffer1072 (.A(\icache.tag_mem.data_i [119]),
    .Z(net1072));
 BUF_X4 buffer1073 (.A(\icache.tag_mem.data_i [119]),
    .Z(net1073));
 BUF_X4 buffer1074 (.A(\icache.tag_mem.data_i [119]),
    .Z(net1074));
 BUF_X4 buffer1075 (.A(\icache.tag_mem.data_i [119]),
    .Z(net1075));
 BUF_X4 buffer1076 (.A(\icache.tag_mem.data_i [119]),
    .Z(net1076));
 BUF_X4 buffer1077 (.A(\icache.tag_mem.data_i [117]),
    .Z(net1077));
 BUF_X4 buffer1078 (.A(\icache.tag_mem.data_i [117]),
    .Z(net1078));
 BUF_X4 buffer1079 (.A(\icache.tag_mem.data_i [117]),
    .Z(net1079));
 BUF_X4 buffer108 (.A(net107),
    .Z(net108));
 BUF_X4 buffer1080 (.A(\icache.tag_mem.data_i [117]),
    .Z(net1080));
 BUF_X4 buffer1081 (.A(\icache.tag_mem.data_i [117]),
    .Z(net1081));
 BUF_X4 buffer1082 (.A(\icache.tag_mem.data_i [117]),
    .Z(net1082));
 BUF_X4 buffer1083 (.A(\icache.tag_mem.data_i [117]),
    .Z(net1083));
 BUF_X4 buffer1084 (.A(\icache.tag_mem.data_i [117]),
    .Z(net1084));
 BUF_X4 buffer1085 (.A(\icache.stat_mem.addr_i [5]),
    .Z(net1085));
 BUF_X4 buffer1086 (.A(\icache.stat_mem.addr_i [4]),
    .Z(net1086));
 BUF_X4 buffer1087 (.A(\icache.stat_mem.addr_i [3]),
    .Z(net1087));
 BUF_X4 buffer1088 (.A(\icache.stat_mem.addr_i [2]),
    .Z(net1088));
 BUF_X4 buffer1089 (.A(\icache.stat_mem.addr_i [1]),
    .Z(net1089));
 BUF_X4 buffer109 (.A(net107),
    .Z(net109));
 BUF_X4 buffer1090 (.A(\icache.stat_mem.addr_i [0]),
    .Z(net1090));
 BUF_X4 buffer1091 (.A(\icache.tag_mem.data_i [115]),
    .Z(net1091));
 BUF_X4 buffer1092 (.A(\icache.tag_mem.data_i [115]),
    .Z(net1092));
 BUF_X4 buffer1093 (.A(\icache.tag_mem.data_i [115]),
    .Z(net1093));
 BUF_X4 buffer1094 (.A(\icache.tag_mem.data_i [115]),
    .Z(net1094));
 BUF_X4 buffer1095 (.A(\icache.tag_mem.data_i [115]),
    .Z(net1095));
 BUF_X4 buffer1096 (.A(\icache.tag_mem.data_i [115]),
    .Z(net1096));
 BUF_X4 buffer1097 (.A(\icache.tag_mem.data_i [115]),
    .Z(net1097));
 BUF_X4 buffer1098 (.A(\icache.tag_mem.data_i [115]),
    .Z(net1098));
 BUF_X4 buffer1099 (.A(\icache.tag_mem.data_i [114]),
    .Z(net1099));
 BUF_X4 buffer11 (.A(_23283_),
    .Z(net11));
 BUF_X4 buffer110 (.A(_10756_),
    .Z(net110));
 BUF_X4 buffer1100 (.A(\icache.tag_mem.data_i [114]),
    .Z(net1100));
 BUF_X4 buffer1101 (.A(\icache.tag_mem.data_i [114]),
    .Z(net1101));
 BUF_X4 buffer1102 (.A(\icache.tag_mem.data_i [114]),
    .Z(net1102));
 BUF_X4 buffer1103 (.A(\icache.tag_mem.data_i [114]),
    .Z(net1103));
 BUF_X4 buffer1104 (.A(\icache.tag_mem.data_i [114]),
    .Z(net1104));
 BUF_X4 buffer1105 (.A(\icache.tag_mem.data_i [114]),
    .Z(net1105));
 BUF_X4 buffer1106 (.A(\icache.tag_mem.data_i [114]),
    .Z(net1106));
 BUF_X4 buffer1107 (.A(\icache.tag_mem.data_i [111]),
    .Z(net1107));
 BUF_X4 buffer1108 (.A(\icache.tag_mem.data_i [111]),
    .Z(net1108));
 BUF_X4 buffer1109 (.A(\icache.tag_mem.data_i [111]),
    .Z(net1109));
 BUF_X4 buffer111 (.A(_10756_),
    .Z(net111));
 BUF_X4 buffer1110 (.A(\icache.tag_mem.data_i [111]),
    .Z(net1110));
 BUF_X4 buffer1111 (.A(\icache.tag_mem.data_i [111]),
    .Z(net1111));
 BUF_X4 buffer1112 (.A(\icache.tag_mem.data_i [111]),
    .Z(net1112));
 BUF_X4 buffer1113 (.A(\icache.tag_mem.data_i [111]),
    .Z(net1113));
 BUF_X4 buffer1114 (.A(\icache.tag_mem.data_i [111]),
    .Z(net1114));
 BUF_X4 buffer1115 (.A(\icache.tag_mem.data_i [107]),
    .Z(net1115));
 BUF_X4 buffer1116 (.A(net1115),
    .Z(net1116));
 BUF_X4 buffer1117 (.A(net1115),
    .Z(net1117));
 BUF_X4 buffer1118 (.A(net1115),
    .Z(net1118));
 BUF_X4 buffer1119 (.A(net1115),
    .Z(net1119));
 BUF_X4 buffer112 (.A(_10756_),
    .Z(net112));
 BUF_X4 buffer1120 (.A(net1115),
    .Z(net1120));
 BUF_X4 buffer1121 (.A(net1115),
    .Z(net1121));
 BUF_X4 buffer1122 (.A(net1115),
    .Z(net1122));
 BUF_X4 buffer1123 (.A(net1115),
    .Z(net1123));
 BUF_X4 buffer1124 (.A(\icache.tag_mem.data_i [106]),
    .Z(net1124));
 BUF_X4 buffer1125 (.A(net1124),
    .Z(net1125));
 BUF_X4 buffer1126 (.A(net1124),
    .Z(net1126));
 BUF_X4 buffer1127 (.A(net1124),
    .Z(net1127));
 BUF_X4 buffer1128 (.A(net1124),
    .Z(net1128));
 BUF_X4 buffer1129 (.A(net1124),
    .Z(net1129));
 BUF_X4 buffer113 (.A(net112),
    .Z(net113));
 BUF_X4 buffer1130 (.A(net1124),
    .Z(net1130));
 BUF_X4 buffer1131 (.A(net1124),
    .Z(net1131));
 BUF_X4 buffer1132 (.A(net1124),
    .Z(net1132));
 BUF_X4 buffer1133 (.A(\icache.tag_mem.data_i [105]),
    .Z(net1133));
 BUF_X4 buffer1134 (.A(\icache.tag_mem.data_i [105]),
    .Z(net1134));
 BUF_X4 buffer1135 (.A(\icache.tag_mem.data_i [105]),
    .Z(net1135));
 BUF_X4 buffer1136 (.A(\icache.tag_mem.data_i [105]),
    .Z(net1136));
 BUF_X4 buffer1137 (.A(\icache.tag_mem.data_i [105]),
    .Z(net1137));
 BUF_X4 buffer1138 (.A(\icache.tag_mem.data_i [105]),
    .Z(net1138));
 BUF_X4 buffer1139 (.A(\icache.tag_mem.data_i [105]),
    .Z(net1139));
 BUF_X4 buffer114 (.A(\icache.data_mem_addr_li [0]),
    .Z(net114));
 BUF_X4 buffer1140 (.A(\icache.tag_mem.data_i [105]),
    .Z(net1140));
 BUF_X4 buffer1141 (.A(\icache.tag_mem.data_i [104]),
    .Z(net1141));
 BUF_X4 buffer1142 (.A(net1141),
    .Z(net1142));
 BUF_X4 buffer1143 (.A(net1141),
    .Z(net1143));
 BUF_X4 buffer1144 (.A(net1141),
    .Z(net1144));
 BUF_X4 buffer1145 (.A(net1141),
    .Z(net1145));
 BUF_X4 buffer1146 (.A(net1141),
    .Z(net1146));
 BUF_X4 buffer1147 (.A(net1141),
    .Z(net1147));
 BUF_X4 buffer1148 (.A(net1141),
    .Z(net1148));
 BUF_X4 buffer1149 (.A(net1141),
    .Z(net1149));
 BUF_X4 buffer115 (.A(net114),
    .Z(net115));
 BUF_X4 buffer1150 (.A(\icache.tag_mem.data_i [101]),
    .Z(net1150));
 BUF_X4 buffer1151 (.A(net1150),
    .Z(net1151));
 BUF_X4 buffer1152 (.A(net1150),
    .Z(net1152));
 BUF_X4 buffer1153 (.A(net1150),
    .Z(net1153));
 BUF_X4 buffer1154 (.A(net1150),
    .Z(net1154));
 BUF_X4 buffer1155 (.A(net1150),
    .Z(net1155));
 BUF_X4 buffer1156 (.A(net1150),
    .Z(net1156));
 BUF_X4 buffer1157 (.A(net1150),
    .Z(net1157));
 BUF_X4 buffer1158 (.A(net1150),
    .Z(net1158));
 BUF_X4 buffer1159 (.A(\icache.tag_mem.data_i [100]),
    .Z(net1159));
 BUF_X4 buffer116 (.A(net114),
    .Z(net116));
 BUF_X4 buffer1160 (.A(net1159),
    .Z(net1160));
 BUF_X4 buffer1161 (.A(net1159),
    .Z(net1161));
 BUF_X4 buffer1162 (.A(net1159),
    .Z(net1162));
 BUF_X4 buffer1163 (.A(net1159),
    .Z(net1163));
 BUF_X4 buffer1164 (.A(net1159),
    .Z(net1164));
 BUF_X4 buffer1165 (.A(net1159),
    .Z(net1165));
 BUF_X4 buffer1166 (.A(net1159),
    .Z(net1166));
 BUF_X4 buffer1167 (.A(net1159),
    .Z(net1167));
 BUF_X4 buffer1168 (.A(\icache.tag_mem.data_i [10]),
    .Z(net1168));
 BUF_X4 buffer1169 (.A(net1168),
    .Z(net1169));
 BUF_X4 buffer117 (.A(net114),
    .Z(net117));
 BUF_X4 buffer1170 (.A(net1168),
    .Z(net1170));
 BUF_X4 buffer1171 (.A(net1168),
    .Z(net1171));
 BUF_X4 buffer1172 (.A(net1168),
    .Z(net1172));
 BUF_X4 buffer1173 (.A(net1168),
    .Z(net1173));
 BUF_X4 buffer1174 (.A(net1168),
    .Z(net1174));
 BUF_X4 buffer1175 (.A(net1168),
    .Z(net1175));
 BUF_X4 buffer1176 (.A(net1168),
    .Z(net1176));
 BUF_X4 buffer1177 (.A(\icache.tag_mem.data_i [123]),
    .Z(net1177));
 BUF_X4 buffer1178 (.A(net1177),
    .Z(net1178));
 BUF_X4 buffer1179 (.A(net1177),
    .Z(net1179));
 BUF_X4 buffer118 (.A(net114),
    .Z(net118));
 BUF_X4 buffer1180 (.A(net1177),
    .Z(net1180));
 BUF_X4 buffer1181 (.A(net1177),
    .Z(net1181));
 BUF_X4 buffer1182 (.A(net1177),
    .Z(net1182));
 BUF_X4 buffer1183 (.A(net1177),
    .Z(net1183));
 BUF_X4 buffer1184 (.A(net1177),
    .Z(net1184));
 BUF_X4 buffer1185 (.A(net1177),
    .Z(net1185));
 BUF_X4 buffer1186 (.A(\icache.tag_mem.data_i [122]),
    .Z(net1186));
 BUF_X4 buffer1187 (.A(net1186),
    .Z(net1187));
 BUF_X4 buffer1188 (.A(net1186),
    .Z(net1188));
 BUF_X4 buffer1189 (.A(net1186),
    .Z(net1189));
 BUF_X4 buffer119 (.A(\icache.data_mem_addr_li [27]),
    .Z(net119));
 BUF_X4 buffer1190 (.A(net1186),
    .Z(net1190));
 BUF_X4 buffer1191 (.A(net1186),
    .Z(net1191));
 BUF_X4 buffer1192 (.A(net1186),
    .Z(net1192));
 BUF_X4 buffer1193 (.A(net1186),
    .Z(net1193));
 BUF_X4 buffer1194 (.A(net1186),
    .Z(net1194));
 BUF_X4 buffer1195 (.A(\icache.tag_mem.data_i [118]),
    .Z(net1195));
 BUF_X4 buffer1196 (.A(net1195),
    .Z(net1196));
 BUF_X4 buffer1197 (.A(net1195),
    .Z(net1197));
 BUF_X4 buffer1198 (.A(net1195),
    .Z(net1198));
 BUF_X4 buffer1199 (.A(net1195),
    .Z(net1199));
 BUF_X4 buffer12 (.A(_25953_),
    .Z(net12));
 BUF_X4 buffer120 (.A(net119),
    .Z(net120));
 BUF_X4 buffer1200 (.A(net1195),
    .Z(net1200));
 BUF_X4 buffer1201 (.A(net1195),
    .Z(net1201));
 BUF_X4 buffer1202 (.A(net1195),
    .Z(net1202));
 BUF_X4 buffer1203 (.A(net1195),
    .Z(net1203));
 BUF_X4 buffer1204 (.A(\icache.tag_mem.data_i [0]),
    .Z(net1204));
 BUF_X4 buffer1205 (.A(net1204),
    .Z(net1205));
 BUF_X4 buffer1206 (.A(net1204),
    .Z(net1206));
 BUF_X4 buffer1207 (.A(net1204),
    .Z(net1207));
 BUF_X4 buffer1208 (.A(net1204),
    .Z(net1208));
 BUF_X4 buffer1209 (.A(net1204),
    .Z(net1209));
 BUF_X4 buffer121 (.A(net119),
    .Z(net121));
 BUF_X4 buffer1210 (.A(net1204),
    .Z(net1210));
 BUF_X4 buffer1211 (.A(net1204),
    .Z(net1211));
 BUF_X4 buffer1212 (.A(net1204),
    .Z(net1212));
 BUF_X4 buffer1213 (.A(_07516_),
    .Z(net1213));
 BUF_X4 buffer1214 (.A(net1213),
    .Z(net1214));
 BUF_X4 buffer1215 (.A(net1214),
    .Z(net1215));
 BUF_X4 buffer1216 (.A(\icache.tag_mem.data_i [113]),
    .Z(net1216));
 BUF_X4 buffer1217 (.A(net1216),
    .Z(net1217));
 BUF_X4 buffer1218 (.A(net1216),
    .Z(net1218));
 BUF_X4 buffer1219 (.A(net1216),
    .Z(net1219));
 BUF_X4 buffer122 (.A(net119),
    .Z(net122));
 BUF_X4 buffer1220 (.A(net1216),
    .Z(net1220));
 BUF_X4 buffer1221 (.A(net1216),
    .Z(net1221));
 BUF_X4 buffer1222 (.A(net1216),
    .Z(net1222));
 BUF_X4 buffer1223 (.A(net1216),
    .Z(net1223));
 BUF_X4 buffer1224 (.A(net1216),
    .Z(net1224));
 BUF_X4 buffer1225 (.A(\icache.tag_mem.data_i [112]),
    .Z(net1225));
 BUF_X4 buffer1226 (.A(net1225),
    .Z(net1226));
 BUF_X4 buffer1227 (.A(net1225),
    .Z(net1227));
 BUF_X4 buffer1228 (.A(net1225),
    .Z(net1228));
 BUF_X4 buffer1229 (.A(net1225),
    .Z(net1229));
 BUF_X4 buffer123 (.A(net119),
    .Z(net123));
 BUF_X4 buffer1230 (.A(net1225),
    .Z(net1230));
 BUF_X4 buffer1231 (.A(net1225),
    .Z(net1231));
 BUF_X4 buffer1232 (.A(net1225),
    .Z(net1232));
 BUF_X4 buffer1233 (.A(net1225),
    .Z(net1233));
 BUF_X4 buffer1234 (.A(\icache.tag_mem.data_i [110]),
    .Z(net1234));
 BUF_X4 buffer1235 (.A(net1234),
    .Z(net1235));
 BUF_X4 buffer1236 (.A(net1234),
    .Z(net1236));
 BUF_X4 buffer1237 (.A(net1234),
    .Z(net1237));
 BUF_X4 buffer1238 (.A(net1234),
    .Z(net1238));
 BUF_X4 buffer1239 (.A(net1234),
    .Z(net1239));
 BUF_X4 buffer124 (.A(\icache.data_mem_addr_li [17]),
    .Z(net124));
 BUF_X4 buffer1240 (.A(net1234),
    .Z(net1240));
 BUF_X4 buffer1241 (.A(net1234),
    .Z(net1241));
 BUF_X4 buffer1242 (.A(net1234),
    .Z(net1242));
 BUF_X4 buffer1243 (.A(\icache.tag_mem.data_i [109]),
    .Z(net1243));
 BUF_X4 buffer1244 (.A(net1243),
    .Z(net1244));
 BUF_X4 buffer1245 (.A(net1243),
    .Z(net1245));
 BUF_X4 buffer1246 (.A(net1243),
    .Z(net1246));
 BUF_X4 buffer1247 (.A(net1243),
    .Z(net1247));
 BUF_X4 buffer1248 (.A(net1243),
    .Z(net1248));
 BUF_X4 buffer1249 (.A(net1243),
    .Z(net1249));
 BUF_X4 buffer125 (.A(net124),
    .Z(net125));
 BUF_X4 buffer1250 (.A(net1243),
    .Z(net1250));
 BUF_X4 buffer1251 (.A(net1243),
    .Z(net1251));
 BUF_X4 buffer1252 (.A(\icache.tag_mem.data_i [108]),
    .Z(net1252));
 BUF_X4 buffer1253 (.A(net1252),
    .Z(net1253));
 BUF_X4 buffer1254 (.A(net1252),
    .Z(net1254));
 BUF_X4 buffer1255 (.A(net1252),
    .Z(net1255));
 BUF_X4 buffer1256 (.A(net1252),
    .Z(net1256));
 BUF_X4 buffer1257 (.A(net1252),
    .Z(net1257));
 BUF_X4 buffer1258 (.A(net1252),
    .Z(net1258));
 BUF_X4 buffer1259 (.A(net1252),
    .Z(net1259));
 BUF_X4 buffer126 (.A(net124),
    .Z(net126));
 BUF_X4 buffer1260 (.A(net1252),
    .Z(net1260));
 BUF_X4 buffer1261 (.A(_07621_),
    .Z(net1261));
 BUF_X4 buffer1262 (.A(net1261),
    .Z(net1262));
 BUF_X4 buffer1263 (.A(\icache.final_data_mux.N0 ),
    .Z(net1263));
 BUF_X4 buffer1264 (.A(net1263),
    .Z(net1264));
 BUF_X4 buffer1265 (.A(\icache.data_set_select_mux.data_i [95]),
    .Z(net1265));
 BUF_X4 buffer1266 (.A(\icache.data_set_select_mux.data_i [94]),
    .Z(net1266));
 BUF_X4 buffer1267 (.A(\icache.tag_tv_r [138]),
    .Z(net1267));
 BUF_X4 buffer1268 (.A(\icache.tag_tv_r [137]),
    .Z(net1268));
 BUF_X4 buffer1269 (.A(\icache.tag_tv_r [136]),
    .Z(net1269));
 BUF_X4 buffer127 (.A(net124),
    .Z(net127));
 BUF_X4 buffer1270 (.A(\icache.tag_tv_r [135]),
    .Z(net1270));
 BUF_X4 buffer1271 (.A(\icache.tag_tv_r [134]),
    .Z(net1271));
 BUF_X4 buffer1272 (.A(\icache.tag_tv_r [133]),
    .Z(net1272));
 BUF_X4 buffer1273 (.A(\icache.tag_tv_r [132]),
    .Z(net1273));
 BUF_X4 buffer1274 (.A(\icache.tag_tv_r [130]),
    .Z(net1274));
 BUF_X4 buffer1275 (.A(\icache.tag_tv_r [129]),
    .Z(net1275));
 BUF_X4 buffer1276 (.A(\icache.tag_tv_r [128]),
    .Z(net1276));
 BUF_X4 buffer1277 (.A(\icache.tag_tv_r [127]),
    .Z(net1277));
 BUF_X4 buffer1278 (.A(\icache.tag_tv_r [126]),
    .Z(net1278));
 BUF_X4 buffer1279 (.A(\icache.tag_tv_r [125]),
    .Z(net1279));
 BUF_X4 buffer128 (.A(net124),
    .Z(net128));
 BUF_X4 buffer1280 (.A(\icache.tag_tv_r [124]),
    .Z(net1280));
 BUF_X4 buffer1281 (.A(net1280),
    .Z(net1281));
 BUF_X4 buffer1282 (.A(net1280),
    .Z(net1282));
 BUF_X4 buffer1283 (.A(\icache.tag_tv_r [123]),
    .Z(net1283));
 BUF_X4 buffer1284 (.A(\icache.tag_tv_r [122]),
    .Z(net1284));
 BUF_X4 buffer1285 (.A(net1284),
    .Z(net1285));
 BUF_X4 buffer1286 (.A(\icache.tag_tv_r [121]),
    .Z(net1286));
 BUF_X4 buffer1287 (.A(net1286),
    .Z(net1287));
 BUF_X4 buffer1288 (.A(\icache.tag_tv_r [120]),
    .Z(net1288));
 BUF_X4 buffer1289 (.A(\icache.tag_tv_r [119]),
    .Z(net1289));
 BUF_X4 buffer129 (.A(net124),
    .Z(net129));
 BUF_X4 buffer1290 (.A(\icache.tag_tv_r [118]),
    .Z(net1290));
 BUF_X4 buffer1291 (.A(\icache.tag_tv_r [117]),
    .Z(net1291));
 BUF_X4 buffer1292 (.A(\icache.tag_tv_r [116]),
    .Z(net1292));
 BUF_X4 buffer1293 (.A(\icache.tag_tv_r [115]),
    .Z(net1293));
 BUF_X4 buffer1294 (.A(net1293),
    .Z(net1294));
 BUF_X4 buffer1295 (.A(net1294),
    .Z(net1295));
 BUF_X4 buffer1296 (.A(\icache.tag_tv_r [114]),
    .Z(net1296));
 BUF_X4 buffer1297 (.A(\icache.tag_tv_r [113]),
    .Z(net1297));
 BUF_X4 buffer1298 (.A(net1297),
    .Z(net1298));
 BUF_X4 buffer1299 (.A(\icache.tag_tv_r [112]),
    .Z(net1299));
 BUF_X4 buffer13 (.A(_25814_),
    .Z(net13));
 BUF_X4 buffer130 (.A(net124),
    .Z(net130));
 BUF_X4 buffer1300 (.A(\icache.tag_tv_r [111]),
    .Z(net1300));
 BUF_X4 buffer1301 (.A(\icache.tag_tv_r [110]),
    .Z(net1301));
 BUF_X4 buffer1302 (.A(\icache.tag_tv_r [109]),
    .Z(net1302));
 BUF_X4 buffer1303 (.A(\icache.read_mux_butterfly.mux_stage_1__mux_swap_0__swap_inst.N0 ),
    .Z(net1303));
 BUF_X4 buffer1304 (.A(net1303),
    .Z(net1304));
 BUF_X4 buffer1305 (.A(net1303),
    .Z(net1305));
 BUF_X4 buffer1306 (.A(net1303),
    .Z(net1306));
 BUF_X4 buffer1307 (.A(\icache.read_mux_butterfly.mux_stage_0__mux_swap_0__swap_inst.N0 ),
    .Z(net1307));
 BUF_X4 buffer1308 (.A(net1307),
    .Z(net1308));
 BUF_X4 buffer1309 (.A(net1307),
    .Z(net1309));
 BUF_X4 buffer131 (.A(net124),
    .Z(net131));
 BUF_X4 buffer1310 (.A(net1307),
    .Z(net1310));
 BUF_X4 buffer1311 (.A(net1307),
    .Z(net1311));
 BUF_X4 buffer1312 (.A(net1307),
    .Z(net1312));
 BUF_X4 buffer1313 (.A(net1307),
    .Z(net1313));
 BUF_X4 buffer1314 (.A(\icache.addr_tv_r [38]),
    .Z(net1314));
 BUF_X4 buffer1315 (.A(net1314),
    .Z(net1315));
 BUF_X4 buffer1316 (.A(net1314),
    .Z(net1316));
 BUF_X4 buffer1317 (.A(\icache.addr_tv_r [37]),
    .Z(net1317));
 BUF_X4 buffer1318 (.A(net1317),
    .Z(net1318));
 BUF_X4 buffer1319 (.A(net1318),
    .Z(net1319));
 BUF_X4 buffer132 (.A(net124),
    .Z(net132));
 BUF_X4 buffer1320 (.A(net1318),
    .Z(net1320));
 BUF_X4 buffer1321 (.A(net1317),
    .Z(net1321));
 BUF_X4 buffer1322 (.A(net1317),
    .Z(net1322));
 BUF_X4 buffer1323 (.A(net1317),
    .Z(net1323));
 BUF_X4 buffer1324 (.A(net1317),
    .Z(net1324));
 BUF_X4 buffer1325 (.A(\icache.addr_tv_r [35]),
    .Z(net1325));
 BUF_X4 buffer1326 (.A(net1325),
    .Z(net1326));
 BUF_X4 buffer1327 (.A(net1325),
    .Z(net1327));
 BUF_X4 buffer1328 (.A(net1325),
    .Z(net1328));
 BUF_X4 buffer1329 (.A(net1325),
    .Z(net1329));
 BUF_X4 buffer133 (.A(\icache.data_mem_addr_li [16]),
    .Z(net133));
 BUF_X4 buffer1330 (.A(\icache.addr_tv_r [33]),
    .Z(net1330));
 BUF_X4 buffer1331 (.A(net1330),
    .Z(net1331));
 BUF_X4 buffer1332 (.A(net1330),
    .Z(net1332));
 BUF_X4 buffer1333 (.A(net1330),
    .Z(net1333));
 BUF_X4 buffer1334 (.A(net1330),
    .Z(net1334));
 BUF_X4 buffer1335 (.A(\icache.addr_tv_r [31]),
    .Z(net1335));
 BUF_X4 buffer1336 (.A(net1335),
    .Z(net1336));
 BUF_X4 buffer1337 (.A(net1335),
    .Z(net1337));
 BUF_X4 buffer1338 (.A(net1337),
    .Z(net1338));
 BUF_X4 buffer1339 (.A(\icache.addr_tv_r [30]),
    .Z(net1339));
 BUF_X4 buffer134 (.A(net133),
    .Z(net134));
 BUF_X4 buffer1340 (.A(\icache.addr_tv_r [30]),
    .Z(net1340));
 BUF_X4 buffer1341 (.A(net1340),
    .Z(net1341));
 BUF_X4 buffer1342 (.A(net1340),
    .Z(net1342));
 BUF_X4 buffer1343 (.A(net1342),
    .Z(net1343));
 BUF_X4 buffer1344 (.A(\icache.addr_tv_r [28]),
    .Z(net1344));
 BUF_X4 buffer1345 (.A(net1344),
    .Z(net1345));
 BUF_X4 buffer1346 (.A(net1345),
    .Z(net1346));
 BUF_X4 buffer1347 (.A(net1345),
    .Z(net1347));
 BUF_X4 buffer1348 (.A(net1345),
    .Z(net1348));
 BUF_X4 buffer1349 (.A(\icache.addr_tv_r [27]),
    .Z(net1349));
 BUF_X4 buffer135 (.A(net133),
    .Z(net135));
 BUF_X4 buffer1350 (.A(net1349),
    .Z(net1350));
 BUF_X4 buffer1351 (.A(\icache.addr_tv_r [24]),
    .Z(net1351));
 BUF_X4 buffer1352 (.A(net1351),
    .Z(net1352));
 BUF_X4 buffer1353 (.A(\icache.addr_tv_r [23]),
    .Z(net1353));
 BUF_X4 buffer1354 (.A(net1353),
    .Z(net1354));
 BUF_X4 buffer1355 (.A(net1354),
    .Z(net1355));
 BUF_X4 buffer1356 (.A(\icache.addr_tv_r [21]),
    .Z(net1356));
 BUF_X4 buffer1357 (.A(net1356),
    .Z(net1357));
 BUF_X4 buffer1358 (.A(net1356),
    .Z(net1358));
 BUF_X4 buffer1359 (.A(net1356),
    .Z(net1359));
 BUF_X4 buffer136 (.A(net133),
    .Z(net136));
 BUF_X4 buffer1360 (.A(net1359),
    .Z(net1360));
 BUF_X4 buffer1361 (.A(\icache.addr_tv_r [19]),
    .Z(net1361));
 BUF_X4 buffer1362 (.A(net1361),
    .Z(net1362));
 BUF_X4 buffer1363 (.A(net1361),
    .Z(net1363));
 BUF_X4 buffer1364 (.A(net1363),
    .Z(net1364));
 BUF_X4 buffer1365 (.A(net1363),
    .Z(net1365));
 BUF_X4 buffer1366 (.A(\icache.addr_tv_r [18]),
    .Z(net1366));
 BUF_X4 buffer1367 (.A(net1366),
    .Z(net1367));
 BUF_X4 buffer1368 (.A(net1366),
    .Z(net1368));
 BUF_X4 buffer1369 (.A(\icache.addr_tv_r [17]),
    .Z(net1369));
 BUF_X4 buffer137 (.A(net133),
    .Z(net137));
 BUF_X4 buffer1370 (.A(net1369),
    .Z(net1370));
 BUF_X4 buffer1371 (.A(net1369),
    .Z(net1371));
 BUF_X4 buffer1372 (.A(net1369),
    .Z(net1372));
 BUF_X4 buffer1373 (.A(net1372),
    .Z(net1373));
 BUF_X4 buffer1374 (.A(\icache.addr_tv_r [15]),
    .Z(net1374));
 BUF_X4 buffer1375 (.A(net1374),
    .Z(net1375));
 BUF_X4 buffer1376 (.A(\icache.addr_tv_r [14]),
    .Z(net1376));
 BUF_X4 buffer1377 (.A(net1376),
    .Z(net1377));
 BUF_X4 buffer1378 (.A(net1376),
    .Z(net1378));
 BUF_X4 buffer1379 (.A(net1376),
    .Z(net1379));
 BUF_X4 buffer138 (.A(net133),
    .Z(net138));
 BUF_X4 buffer1380 (.A(\icache.addr_tv_r [13]),
    .Z(net1380));
 BUF_X4 buffer1381 (.A(net1380),
    .Z(net1381));
 BUF_X4 buffer1382 (.A(net1380),
    .Z(net1382));
 BUF_X4 buffer1383 (.A(net1382),
    .Z(net1383));
 BUF_X4 buffer1384 (.A(net1383),
    .Z(net1384));
 BUF_X4 buffer1385 (.A(\icache.addr_tv_r [12]),
    .Z(net1385));
 BUF_X4 buffer1386 (.A(\icache.addr_tv_r [12]),
    .Z(net1386));
 BUF_X4 buffer1387 (.A(net1386),
    .Z(net1387));
 BUF_X4 buffer1388 (.A(net1386),
    .Z(net1388));
 BUF_X4 buffer1389 (.A(\icache.N12 ),
    .Z(net1389));
 BUF_X4 buffer139 (.A(net133),
    .Z(net139));
 BUF_X4 buffer1390 (.A(net1389),
    .Z(net1390));
 BUF_X4 buffer1391 (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [728]),
    .Z(net1391));
 BUF_X4 buffer1392 (.A(\bp_fe_pc_gen_1.btb.tag_mem.z_s1r1w_mem.synth.mem [696]),
    .Z(net1392));
 BUF_X4 buffer1393 (.A(\icache.lce.lce_data_cmd.rv_adapter.head_r ),
    .Z(net1393));
 BUF_X4 buffer1394 (.A(net1393),
    .Z(net1394));
 BUF_X4 buffer1395 (.A(net1393),
    .Z(net1395));
 BUF_X4 buffer1396 (.A(net1393),
    .Z(net1396));
 BUF_X4 buffer1397 (.A(\icache.lce.N14 ),
    .Z(net1397));
 BUF_X4 buffer1398 (.A(\bp_fe_pc_gen_1.btb.tag_mem.data_o [46]),
    .Z(net1398));
 BUF_X4 buffer1399 (.A(\bp_fe_pc_gen_1.btb.tag_mem.data_o [45]),
    .Z(net1399));
 BUF_X4 buffer14 (.A(_24113_),
    .Z(net14));
 BUF_X4 buffer140 (.A(net133),
    .Z(net140));
 BUF_X4 buffer1400 (.A(\bp_fe_pc_gen_1.btb.tag_mem.data_o [42]),
    .Z(net1400));
 BUF_X4 buffer1401 (.A(\bp_fe_pc_gen_1.btb.tag_mem.data_o [41]),
    .Z(net1401));
 BUF_X4 buffer1402 (.A(\bp_fe_pc_gen_1.btb.br_tgt_o [38]),
    .Z(net1402));
 BUF_X4 buffer1403 (.A(\bp_fe_pc_gen_1.btb.br_tgt_o [33]),
    .Z(net1403));
 BUF_X4 buffer1404 (.A(\bp_fe_pc_gen_1.btb.br_tgt_o [32]),
    .Z(net1404));
 BUF_X4 buffer1405 (.A(\bp_fe_pc_gen_1.btb.br_tgt_o [31]),
    .Z(net1405));
 BUF_X4 buffer1406 (.A(\bp_fe_pc_gen_1.btb.br_tgt_o [22]),
    .Z(net1406));
 BUF_X4 buffer1407 (.A(\bp_fe_pc_gen_1.btb.br_tgt_o [21]),
    .Z(net1407));
 BUF_X4 buffer1408 (.A(\bp_fe_pc_gen_1.btb.br_tgt_o [19]),
    .Z(net1408));
 BUF_X4 buffer1409 (.A(\bp_fe_pc_gen_1.btb.br_tgt_o [18]),
    .Z(net1409));
 BUF_X4 buffer141 (.A(net133),
    .Z(net141));
 BUF_X4 buffer1410 (.A(\bp_fe_pc_gen_1.btb.br_tgt_o [16]),
    .Z(net1410));
 BUF_X4 buffer1411 (.A(\bp_fe_pc_gen_1.btb.br_tgt_o [15]),
    .Z(net1411));
 BUF_X4 buffer1412 (.A(\bp_fe_pc_gen_1.btb.br_tgt_o [14]),
    .Z(net1412));
 BUF_X4 buffer1413 (.A(\bp_fe_pc_gen_1.btb.br_tgt_o [10]),
    .Z(net1413));
 BUF_X4 buffer1414 (.A(\bp_fe_pc_gen_1.btb.br_tgt_o [9]),
    .Z(net1414));
 BUF_X4 buffer1415 (.A(\bp_fe_pc_gen_1.btb.br_tgt_o [5]),
    .Z(net1415));
 BUF_X4 buffer1416 (.A(\bp_fe_pc_gen_1.btb.br_tgt_o [1]),
    .Z(net1416));
 BUF_X4 buffer1417 (.A(\bp_fe_pc_gen_1.btb.br_tgt_o [0]),
    .Z(net1417));
 BUF_X4 buffer1418 (.A(\icache.lce.lce_cmd_inst.N10 ),
    .Z(net1418));
 BUF_X4 buffer1419 (.A(net1418),
    .Z(net1419));
 BUF_X4 buffer142 (.A(\icache.data_mem_addr_li [15]),
    .Z(net142));
 BUF_X4 buffer143 (.A(net142),
    .Z(net143));
 BUF_X4 buffer144 (.A(net142),
    .Z(net144));
 BUF_X4 buffer145 (.A(net142),
    .Z(net145));
 BUF_X4 buffer146 (.A(net142),
    .Z(net146));
 BUF_X4 buffer147 (.A(net142),
    .Z(net147));
 BUF_X4 buffer148 (.A(net142),
    .Z(net148));
 BUF_X4 buffer149 (.A(net142),
    .Z(net149));
 BUF_X4 buffer15 (.A(_23960_),
    .Z(net15));
 BUF_X4 buffer150 (.A(net142),
    .Z(net150));
 BUF_X4 buffer151 (.A(\icache.data_mem_addr_li [14]),
    .Z(net151));
 BUF_X4 buffer152 (.A(net151),
    .Z(net152));
 BUF_X4 buffer153 (.A(net151),
    .Z(net153));
 BUF_X4 buffer154 (.A(net151),
    .Z(net154));
 BUF_X4 buffer155 (.A(net151),
    .Z(net155));
 BUF_X4 buffer156 (.A(net151),
    .Z(net156));
 BUF_X4 buffer157 (.A(net151),
    .Z(net157));
 BUF_X4 buffer158 (.A(net151),
    .Z(net158));
 BUF_X4 buffer159 (.A(net151),
    .Z(net159));
 BUF_X4 buffer16 (.A(_23450_),
    .Z(net16));
 BUF_X4 buffer160 (.A(\icache.data_mem_addr_li [11]),
    .Z(net160));
 BUF_X4 buffer161 (.A(net160),
    .Z(net161));
 BUF_X4 buffer162 (.A(net160),
    .Z(net162));
 BUF_X4 buffer163 (.A(net160),
    .Z(net163));
 BUF_X4 buffer164 (.A(net160),
    .Z(net164));
 BUF_X4 buffer165 (.A(\icache.data_mem_addr_li [10]),
    .Z(net165));
 BUF_X4 buffer166 (.A(net165),
    .Z(net166));
 BUF_X4 buffer167 (.A(net165),
    .Z(net167));
 BUF_X4 buffer168 (.A(net165),
    .Z(net168));
 BUF_X4 buffer169 (.A(net165),
    .Z(net169));
 BUF_X4 buffer17 (.A(_25782_),
    .Z(net17));
 BUF_X4 buffer170 (.A(\icache.data_mem_addr_li [19]),
    .Z(net170));
 BUF_X4 buffer171 (.A(net170),
    .Z(net171));
 BUF_X4 buffer172 (.A(net170),
    .Z(net172));
 BUF_X4 buffer173 (.A(net170),
    .Z(net173));
 BUF_X4 buffer174 (.A(net170),
    .Z(net174));
 BUF_X4 buffer175 (.A(\icache.data_mem_addr_li [38]),
    .Z(net175));
 BUF_X4 buffer176 (.A(net175),
    .Z(net176));
 BUF_X4 buffer177 (.A(net175),
    .Z(net177));
 BUF_X4 buffer178 (.A(net175),
    .Z(net178));
 BUF_X4 buffer179 (.A(net175),
    .Z(net179));
 BUF_X4 buffer18 (.A(_25742_),
    .Z(net18));
 BUF_X4 buffer180 (.A(\icache.tag_mem.addr_i [5]),
    .Z(net180));
 BUF_X4 buffer181 (.A(\icache.tag_mem.addr_i [5]),
    .Z(net181));
 BUF_X4 buffer182 (.A(\icache.tag_mem.addr_i [4]),
    .Z(net182));
 BUF_X4 buffer183 (.A(\icache.tag_mem.addr_i [4]),
    .Z(net183));
 BUF_X4 buffer184 (.A(\icache.tag_mem.addr_i [3]),
    .Z(net184));
 BUF_X4 buffer185 (.A(\icache.tag_mem.addr_i [3]),
    .Z(net185));
 BUF_X4 buffer186 (.A(\icache.tag_mem.addr_i [2]),
    .Z(net186));
 BUF_X4 buffer187 (.A(\icache.tag_mem.addr_i [2]),
    .Z(net187));
 BUF_X4 buffer188 (.A(\icache.data_mem_addr_li [13]),
    .Z(net188));
 BUF_X4 buffer189 (.A(net188),
    .Z(net189));
 BUF_X4 buffer19 (.A(_25618_),
    .Z(net19));
 BUF_X4 buffer190 (.A(net188),
    .Z(net190));
 BUF_X4 buffer191 (.A(net188),
    .Z(net191));
 BUF_X4 buffer192 (.A(net188),
    .Z(net192));
 BUF_X4 buffer193 (.A(net188),
    .Z(net193));
 BUF_X4 buffer194 (.A(net188),
    .Z(net194));
 BUF_X4 buffer195 (.A(net188),
    .Z(net195));
 BUF_X4 buffer196 (.A(net188),
    .Z(net196));
 BUF_X4 buffer197 (.A(\icache.data_mem_addr_li [12]),
    .Z(net197));
 BUF_X4 buffer198 (.A(net197),
    .Z(net198));
 BUF_X4 buffer199 (.A(net197),
    .Z(net199));
 BUF_X4 buffer2 (.A(_25579_),
    .Z(net2));
 BUF_X4 buffer20 (.A(_25616_),
    .Z(net20));
 BUF_X4 buffer200 (.A(net197),
    .Z(net200));
 BUF_X4 buffer201 (.A(net197),
    .Z(net201));
 BUF_X4 buffer202 (.A(net197),
    .Z(net202));
 BUF_X4 buffer203 (.A(net197),
    .Z(net203));
 BUF_X4 buffer204 (.A(net197),
    .Z(net204));
 BUF_X4 buffer205 (.A(net197),
    .Z(net205));
 BUF_X4 buffer206 (.A(\icache.tag_mem.addr_i [1]),
    .Z(net206));
 BUF_X4 buffer207 (.A(\icache.tag_mem.addr_i [1]),
    .Z(net207));
 BUF_X4 buffer208 (.A(\icache.tag_mem.addr_i [0]),
    .Z(net208));
 BUF_X4 buffer209 (.A(\icache.tag_mem.addr_i [0]),
    .Z(net209));
 BUF_X4 buffer21 (.A(_25499_),
    .Z(net21));
 BUF_X4 buffer210 (.A(_08848_),
    .Z(net210));
 BUF_X4 buffer211 (.A(net210),
    .Z(net211));
 BUF_X4 buffer212 (.A(_08800_),
    .Z(net212));
 BUF_X4 buffer213 (.A(\icache.data_mem_w_li ),
    .Z(net213));
 BUF_X4 buffer214 (.A(net213),
    .Z(net214));
 BUF_X4 buffer215 (.A(net213),
    .Z(net215));
 BUF_X4 buffer216 (.A(net213),
    .Z(net216));
 BUF_X4 buffer217 (.A(net213),
    .Z(net217));
 BUF_X4 buffer218 (.A(net213),
    .Z(net218));
 BUF_X4 buffer219 (.A(net213),
    .Z(net219));
 BUF_X4 buffer22 (.A(_24984_),
    .Z(net22));
 BUF_X4 buffer220 (.A(net213),
    .Z(net220));
 BUF_X4 buffer221 (.A(net213),
    .Z(net221));
 BUF_X4 buffer222 (.A(\icache.n_0_net_ ),
    .Z(net222));
 BUF_X4 buffer223 (.A(net222),
    .Z(net223));
 BUF_X4 buffer224 (.A(net222),
    .Z(net224));
 BUF_X4 buffer225 (.A(\icache.data_mems_0__data_mem.v_i ),
    .Z(net225));
 BUF_X4 buffer226 (.A(net225),
    .Z(net226));
 BUF_X4 buffer227 (.A(net225),
    .Z(net227));
 BUF_X4 buffer228 (.A(net225),
    .Z(net228));
 BUF_X4 buffer229 (.A(net225),
    .Z(net229));
 BUF_X4 buffer23 (.A(_24951_),
    .Z(net23));
 BUF_X4 buffer230 (.A(net225),
    .Z(net230));
 BUF_X4 buffer231 (.A(net225),
    .Z(net231));
 BUF_X4 buffer232 (.A(net225),
    .Z(net232));
 BUF_X4 buffer233 (.A(net225),
    .Z(net233));
 BUF_X4 buffer234 (.A(\icache.lce.lce_cmd_inst.tag_mem_pkt_yumi_i ),
    .Z(net234));
 BUF_X4 buffer235 (.A(net234),
    .Z(net235));
 BUF_X4 buffer236 (.A(net234),
    .Z(net236));
 BUF_X4 buffer237 (.A(net234),
    .Z(net237));
 BUF_X4 buffer238 (.A(\icache.data_mem_data_li [511]),
    .Z(net238));
 BUF_X4 buffer239 (.A(\icache.data_mem_data_li [510]),
    .Z(net239));
 BUF_X4 buffer24 (.A(_24885_),
    .Z(net24));
 BUF_X4 buffer240 (.A(\icache.data_mem_data_li [509]),
    .Z(net240));
 BUF_X4 buffer241 (.A(\icache.data_mem_data_li [508]),
    .Z(net241));
 BUF_X4 buffer242 (.A(\icache.data_mem_data_li [507]),
    .Z(net242));
 BUF_X4 buffer243 (.A(\icache.data_mem_data_li [506]),
    .Z(net243));
 BUF_X4 buffer244 (.A(\icache.data_mem_data_li [505]),
    .Z(net244));
 BUF_X4 buffer245 (.A(\icache.data_mem_data_li [504]),
    .Z(net245));
 BUF_X4 buffer246 (.A(\icache.data_mem_data_li [503]),
    .Z(net246));
 BUF_X4 buffer247 (.A(\icache.data_mem_data_li [502]),
    .Z(net247));
 BUF_X4 buffer248 (.A(\icache.data_mem_data_li [501]),
    .Z(net248));
 BUF_X4 buffer249 (.A(\icache.data_mem_data_li [500]),
    .Z(net249));
 BUF_X4 buffer25 (.A(_24768_),
    .Z(net25));
 BUF_X4 buffer250 (.A(\icache.data_mem_data_li [499]),
    .Z(net250));
 BUF_X4 buffer251 (.A(\icache.data_mem_data_li [498]),
    .Z(net251));
 BUF_X4 buffer252 (.A(\icache.data_mem_data_li [497]),
    .Z(net252));
 BUF_X4 buffer253 (.A(\icache.data_mem_data_li [496]),
    .Z(net253));
 BUF_X4 buffer254 (.A(\icache.data_mem_data_li [495]),
    .Z(net254));
 BUF_X4 buffer255 (.A(\icache.data_mem_data_li [494]),
    .Z(net255));
 BUF_X4 buffer256 (.A(\icache.data_mem_data_li [493]),
    .Z(net256));
 BUF_X4 buffer257 (.A(\icache.data_mem_data_li [492]),
    .Z(net257));
 BUF_X4 buffer258 (.A(\icache.data_mem_data_li [491]),
    .Z(net258));
 BUF_X4 buffer259 (.A(\icache.data_mem_data_li [490]),
    .Z(net259));
 BUF_X4 buffer26 (.A(_24711_),
    .Z(net26));
 BUF_X4 buffer260 (.A(\icache.data_mem_data_li [489]),
    .Z(net260));
 BUF_X4 buffer261 (.A(\icache.data_mem_data_li [488]),
    .Z(net261));
 BUF_X4 buffer262 (.A(\icache.data_mem_data_li [487]),
    .Z(net262));
 BUF_X4 buffer263 (.A(\icache.data_mem_data_li [486]),
    .Z(net263));
 BUF_X4 buffer264 (.A(\icache.data_mem_data_li [485]),
    .Z(net264));
 BUF_X4 buffer265 (.A(\icache.data_mem_data_li [484]),
    .Z(net265));
 BUF_X4 buffer266 (.A(\icache.data_mem_data_li [483]),
    .Z(net266));
 BUF_X4 buffer267 (.A(\icache.data_mem_data_li [482]),
    .Z(net267));
 BUF_X4 buffer268 (.A(\icache.data_mem_data_li [481]),
    .Z(net268));
 BUF_X4 buffer269 (.A(\icache.data_mem_data_li [480]),
    .Z(net269));
 BUF_X4 buffer27 (.A(_24603_),
    .Z(net27));
 BUF_X4 buffer270 (.A(\icache.data_mem_data_li [479]),
    .Z(net270));
 BUF_X4 buffer271 (.A(\icache.data_mem_data_li [478]),
    .Z(net271));
 BUF_X4 buffer272 (.A(\icache.data_mem_data_li [477]),
    .Z(net272));
 BUF_X4 buffer273 (.A(\icache.data_mem_data_li [476]),
    .Z(net273));
 BUF_X4 buffer274 (.A(\icache.data_mem_data_li [475]),
    .Z(net274));
 BUF_X4 buffer275 (.A(\icache.data_mem_data_li [474]),
    .Z(net275));
 BUF_X4 buffer276 (.A(\icache.data_mem_data_li [473]),
    .Z(net276));
 BUF_X4 buffer277 (.A(\icache.data_mem_data_li [472]),
    .Z(net277));
 BUF_X4 buffer278 (.A(\icache.data_mem_data_li [471]),
    .Z(net278));
 BUF_X4 buffer279 (.A(\icache.data_mem_data_li [470]),
    .Z(net279));
 BUF_X4 buffer28 (.A(_24527_),
    .Z(net28));
 BUF_X4 buffer280 (.A(\icache.data_mem_data_li [469]),
    .Z(net280));
 BUF_X4 buffer281 (.A(\icache.data_mem_data_li [468]),
    .Z(net281));
 BUF_X4 buffer282 (.A(\icache.data_mem_data_li [467]),
    .Z(net282));
 BUF_X4 buffer283 (.A(\icache.data_mem_data_li [466]),
    .Z(net283));
 BUF_X4 buffer284 (.A(\icache.data_mem_data_li [465]),
    .Z(net284));
 BUF_X4 buffer285 (.A(\icache.data_mem_data_li [464]),
    .Z(net285));
 BUF_X4 buffer286 (.A(\icache.data_mem_data_li [463]),
    .Z(net286));
 BUF_X4 buffer287 (.A(\icache.data_mem_data_li [462]),
    .Z(net287));
 BUF_X4 buffer288 (.A(\icache.data_mem_data_li [461]),
    .Z(net288));
 BUF_X4 buffer289 (.A(\icache.data_mem_data_li [460]),
    .Z(net289));
 BUF_X4 buffer29 (.A(_24524_),
    .Z(net29));
 BUF_X4 buffer290 (.A(\icache.data_mem_data_li [459]),
    .Z(net290));
 BUF_X4 buffer291 (.A(\icache.data_mem_data_li [458]),
    .Z(net291));
 BUF_X4 buffer292 (.A(\icache.data_mem_data_li [457]),
    .Z(net292));
 BUF_X4 buffer293 (.A(\icache.data_mem_data_li [456]),
    .Z(net293));
 BUF_X4 buffer294 (.A(\icache.data_mem_data_li [455]),
    .Z(net294));
 BUF_X4 buffer295 (.A(\icache.data_mem_data_li [454]),
    .Z(net295));
 BUF_X4 buffer296 (.A(\icache.data_mem_data_li [453]),
    .Z(net296));
 BUF_X4 buffer297 (.A(\icache.data_mem_data_li [452]),
    .Z(net297));
 BUF_X4 buffer298 (.A(\icache.data_mem_data_li [451]),
    .Z(net298));
 BUF_X4 buffer299 (.A(\icache.data_mem_data_li [450]),
    .Z(net299));
 BUF_X4 buffer3 (.A(_24809_),
    .Z(net3));
 BUF_X4 buffer30 (.A(_24370_),
    .Z(net30));
 BUF_X4 buffer300 (.A(\icache.data_mem_data_li [449]),
    .Z(net300));
 BUF_X4 buffer301 (.A(\icache.data_mem_data_li [448]),
    .Z(net301));
 BUF_X4 buffer302 (.A(\icache.data_mem_data_li [447]),
    .Z(net302));
 BUF_X4 buffer303 (.A(\icache.data_mem_data_li [446]),
    .Z(net303));
 BUF_X4 buffer304 (.A(\icache.data_mem_data_li [445]),
    .Z(net304));
 BUF_X4 buffer305 (.A(\icache.data_mem_data_li [444]),
    .Z(net305));
 BUF_X4 buffer306 (.A(\icache.data_mem_data_li [443]),
    .Z(net306));
 BUF_X4 buffer307 (.A(\icache.data_mem_data_li [442]),
    .Z(net307));
 BUF_X4 buffer308 (.A(\icache.data_mem_data_li [441]),
    .Z(net308));
 BUF_X4 buffer309 (.A(\icache.data_mem_data_li [440]),
    .Z(net309));
 BUF_X4 buffer31 (.A(_24271_),
    .Z(net31));
 BUF_X4 buffer310 (.A(\icache.data_mem_data_li [439]),
    .Z(net310));
 BUF_X4 buffer311 (.A(\icache.data_mem_data_li [438]),
    .Z(net311));
 BUF_X4 buffer312 (.A(\icache.data_mem_data_li [437]),
    .Z(net312));
 BUF_X4 buffer313 (.A(\icache.data_mem_data_li [436]),
    .Z(net313));
 BUF_X4 buffer314 (.A(\icache.data_mem_data_li [435]),
    .Z(net314));
 BUF_X4 buffer315 (.A(\icache.data_mem_data_li [434]),
    .Z(net315));
 BUF_X4 buffer316 (.A(\icache.data_mem_data_li [433]),
    .Z(net316));
 BUF_X4 buffer317 (.A(\icache.data_mem_data_li [432]),
    .Z(net317));
 BUF_X4 buffer318 (.A(\icache.data_mem_data_li [431]),
    .Z(net318));
 BUF_X4 buffer319 (.A(\icache.data_mem_data_li [430]),
    .Z(net319));
 BUF_X4 buffer32 (.A(_24230_),
    .Z(net32));
 BUF_X4 buffer320 (.A(\icache.data_mem_data_li [429]),
    .Z(net320));
 BUF_X4 buffer321 (.A(\icache.data_mem_data_li [428]),
    .Z(net321));
 BUF_X4 buffer322 (.A(\icache.data_mem_data_li [427]),
    .Z(net322));
 BUF_X4 buffer323 (.A(\icache.data_mem_data_li [426]),
    .Z(net323));
 BUF_X4 buffer324 (.A(\icache.data_mem_data_li [425]),
    .Z(net324));
 BUF_X4 buffer325 (.A(\icache.data_mem_data_li [424]),
    .Z(net325));
 BUF_X4 buffer326 (.A(\icache.data_mem_data_li [423]),
    .Z(net326));
 BUF_X4 buffer327 (.A(\icache.data_mem_data_li [422]),
    .Z(net327));
 BUF_X4 buffer328 (.A(\icache.data_mem_data_li [421]),
    .Z(net328));
 BUF_X4 buffer329 (.A(\icache.data_mem_data_li [420]),
    .Z(net329));
 BUF_X4 buffer33 (.A(_24195_),
    .Z(net33));
 BUF_X4 buffer330 (.A(\icache.data_mem_data_li [419]),
    .Z(net330));
 BUF_X4 buffer331 (.A(\icache.data_mem_data_li [418]),
    .Z(net331));
 BUF_X4 buffer332 (.A(\icache.data_mem_data_li [417]),
    .Z(net332));
 BUF_X4 buffer333 (.A(\icache.data_mem_data_li [416]),
    .Z(net333));
 BUF_X4 buffer334 (.A(\icache.data_mem_data_li [415]),
    .Z(net334));
 BUF_X4 buffer335 (.A(\icache.data_mem_data_li [414]),
    .Z(net335));
 BUF_X4 buffer336 (.A(\icache.data_mem_data_li [413]),
    .Z(net336));
 BUF_X4 buffer337 (.A(\icache.data_mem_data_li [412]),
    .Z(net337));
 BUF_X4 buffer338 (.A(\icache.data_mem_data_li [411]),
    .Z(net338));
 BUF_X4 buffer339 (.A(\icache.data_mem_data_li [410]),
    .Z(net339));
 BUF_X4 buffer34 (.A(_24121_),
    .Z(net34));
 BUF_X4 buffer340 (.A(\icache.data_mem_data_li [409]),
    .Z(net340));
 BUF_X4 buffer341 (.A(\icache.data_mem_data_li [408]),
    .Z(net341));
 BUF_X4 buffer342 (.A(\icache.data_mem_data_li [407]),
    .Z(net342));
 BUF_X4 buffer343 (.A(\icache.data_mem_data_li [406]),
    .Z(net343));
 BUF_X4 buffer344 (.A(\icache.data_mem_data_li [405]),
    .Z(net344));
 BUF_X4 buffer345 (.A(\icache.data_mem_data_li [404]),
    .Z(net345));
 BUF_X4 buffer346 (.A(\icache.data_mem_data_li [403]),
    .Z(net346));
 BUF_X4 buffer347 (.A(\icache.data_mem_data_li [402]),
    .Z(net347));
 BUF_X4 buffer348 (.A(\icache.data_mem_data_li [401]),
    .Z(net348));
 BUF_X4 buffer349 (.A(\icache.data_mem_data_li [400]),
    .Z(net349));
 BUF_X4 buffer35 (.A(_24117_),
    .Z(net35));
 BUF_X4 buffer350 (.A(\icache.data_mem_data_li [399]),
    .Z(net350));
 BUF_X4 buffer351 (.A(\icache.data_mem_data_li [398]),
    .Z(net351));
 BUF_X4 buffer352 (.A(\icache.data_mem_data_li [397]),
    .Z(net352));
 BUF_X4 buffer353 (.A(\icache.data_mem_data_li [396]),
    .Z(net353));
 BUF_X4 buffer354 (.A(\icache.data_mem_data_li [395]),
    .Z(net354));
 BUF_X4 buffer355 (.A(\icache.data_mem_data_li [394]),
    .Z(net355));
 BUF_X4 buffer356 (.A(\icache.data_mem_data_li [393]),
    .Z(net356));
 BUF_X4 buffer357 (.A(\icache.data_mem_data_li [392]),
    .Z(net357));
 BUF_X4 buffer358 (.A(\icache.data_mem_data_li [391]),
    .Z(net358));
 BUF_X4 buffer359 (.A(\icache.data_mem_data_li [390]),
    .Z(net359));
 BUF_X4 buffer36 (.A(_23874_),
    .Z(net36));
 BUF_X4 buffer360 (.A(\icache.data_mem_data_li [389]),
    .Z(net360));
 BUF_X4 buffer361 (.A(\icache.data_mem_data_li [388]),
    .Z(net361));
 BUF_X4 buffer362 (.A(\icache.data_mem_data_li [387]),
    .Z(net362));
 BUF_X4 buffer363 (.A(\icache.data_mem_data_li [386]),
    .Z(net363));
 BUF_X4 buffer364 (.A(\icache.data_mem_data_li [385]),
    .Z(net364));
 BUF_X4 buffer365 (.A(\icache.data_mem_data_li [384]),
    .Z(net365));
 BUF_X4 buffer366 (.A(\icache.data_mem_data_li [383]),
    .Z(net366));
 BUF_X4 buffer367 (.A(\icache.data_mem_data_li [382]),
    .Z(net367));
 BUF_X4 buffer368 (.A(\icache.data_mem_data_li [381]),
    .Z(net368));
 BUF_X4 buffer369 (.A(\icache.data_mem_data_li [380]),
    .Z(net369));
 BUF_X4 buffer37 (.A(_23782_),
    .Z(net37));
 BUF_X4 buffer370 (.A(\icache.data_mem_data_li [379]),
    .Z(net370));
 BUF_X4 buffer371 (.A(\icache.data_mem_data_li [378]),
    .Z(net371));
 BUF_X4 buffer372 (.A(\icache.data_mem_data_li [377]),
    .Z(net372));
 BUF_X4 buffer373 (.A(\icache.data_mem_data_li [376]),
    .Z(net373));
 BUF_X4 buffer374 (.A(\icache.data_mem_data_li [375]),
    .Z(net374));
 BUF_X4 buffer375 (.A(\icache.data_mem_data_li [374]),
    .Z(net375));
 BUF_X4 buffer376 (.A(\icache.data_mem_data_li [373]),
    .Z(net376));
 BUF_X4 buffer377 (.A(\icache.data_mem_data_li [372]),
    .Z(net377));
 BUF_X4 buffer378 (.A(\icache.data_mem_data_li [371]),
    .Z(net378));
 BUF_X4 buffer379 (.A(\icache.data_mem_data_li [370]),
    .Z(net379));
 BUF_X4 buffer38 (.A(_23497_),
    .Z(net38));
 BUF_X4 buffer380 (.A(\icache.data_mem_data_li [369]),
    .Z(net380));
 BUF_X4 buffer381 (.A(\icache.data_mem_data_li [368]),
    .Z(net381));
 BUF_X4 buffer382 (.A(\icache.data_mem_data_li [367]),
    .Z(net382));
 BUF_X4 buffer383 (.A(\icache.data_mem_data_li [366]),
    .Z(net383));
 BUF_X4 buffer384 (.A(\icache.data_mem_data_li [365]),
    .Z(net384));
 BUF_X4 buffer385 (.A(\icache.data_mem_data_li [364]),
    .Z(net385));
 BUF_X4 buffer386 (.A(\icache.data_mem_data_li [363]),
    .Z(net386));
 BUF_X4 buffer387 (.A(\icache.data_mem_data_li [362]),
    .Z(net387));
 BUF_X4 buffer388 (.A(\icache.data_mem_data_li [361]),
    .Z(net388));
 BUF_X4 buffer389 (.A(\icache.data_mem_data_li [360]),
    .Z(net389));
 BUF_X4 buffer39 (.A(_23486_),
    .Z(net39));
 BUF_X4 buffer390 (.A(\icache.data_mem_data_li [359]),
    .Z(net390));
 BUF_X4 buffer391 (.A(\icache.data_mem_data_li [358]),
    .Z(net391));
 BUF_X4 buffer392 (.A(\icache.data_mem_data_li [357]),
    .Z(net392));
 BUF_X4 buffer393 (.A(\icache.data_mem_data_li [356]),
    .Z(net393));
 BUF_X4 buffer394 (.A(\icache.data_mem_data_li [355]),
    .Z(net394));
 BUF_X4 buffer395 (.A(\icache.data_mem_data_li [354]),
    .Z(net395));
 BUF_X4 buffer396 (.A(\icache.data_mem_data_li [353]),
    .Z(net396));
 BUF_X4 buffer397 (.A(\icache.data_mem_data_li [352]),
    .Z(net397));
 BUF_X4 buffer398 (.A(\icache.data_mem_data_li [351]),
    .Z(net398));
 BUF_X4 buffer399 (.A(\icache.data_mem_data_li [350]),
    .Z(net399));
 BUF_X4 buffer4 (.A(_24038_),
    .Z(net4));
 BUF_X4 buffer40 (.A(_23220_),
    .Z(net40));
 BUF_X4 buffer400 (.A(\icache.data_mem_data_li [349]),
    .Z(net400));
 BUF_X4 buffer401 (.A(\icache.data_mem_data_li [348]),
    .Z(net401));
 BUF_X4 buffer402 (.A(\icache.data_mem_data_li [347]),
    .Z(net402));
 BUF_X4 buffer403 (.A(\icache.data_mem_data_li [346]),
    .Z(net403));
 BUF_X4 buffer404 (.A(\icache.data_mem_data_li [345]),
    .Z(net404));
 BUF_X4 buffer405 (.A(\icache.data_mem_data_li [344]),
    .Z(net405));
 BUF_X4 buffer406 (.A(\icache.data_mem_data_li [343]),
    .Z(net406));
 BUF_X4 buffer407 (.A(\icache.data_mem_data_li [342]),
    .Z(net407));
 BUF_X4 buffer408 (.A(\icache.data_mem_data_li [341]),
    .Z(net408));
 BUF_X4 buffer409 (.A(\icache.data_mem_data_li [340]),
    .Z(net409));
 BUF_X4 buffer41 (.A(_26262_),
    .Z(net41));
 BUF_X4 buffer410 (.A(\icache.data_mem_data_li [339]),
    .Z(net410));
 BUF_X4 buffer411 (.A(\icache.data_mem_data_li [338]),
    .Z(net411));
 BUF_X4 buffer412 (.A(\icache.data_mem_data_li [337]),
    .Z(net412));
 BUF_X4 buffer413 (.A(\icache.data_mem_data_li [336]),
    .Z(net413));
 BUF_X4 buffer414 (.A(\icache.data_mem_data_li [335]),
    .Z(net414));
 BUF_X4 buffer415 (.A(\icache.data_mem_data_li [334]),
    .Z(net415));
 BUF_X4 buffer416 (.A(\icache.data_mem_data_li [333]),
    .Z(net416));
 BUF_X4 buffer417 (.A(\icache.data_mem_data_li [332]),
    .Z(net417));
 BUF_X4 buffer418 (.A(\icache.data_mem_data_li [331]),
    .Z(net418));
 BUF_X4 buffer419 (.A(\icache.data_mem_data_li [330]),
    .Z(net419));
 BUF_X4 buffer42 (.A(_26253_),
    .Z(net42));
 BUF_X4 buffer420 (.A(\icache.data_mem_data_li [329]),
    .Z(net420));
 BUF_X4 buffer421 (.A(\icache.data_mem_data_li [328]),
    .Z(net421));
 BUF_X4 buffer422 (.A(\icache.data_mem_data_li [327]),
    .Z(net422));
 BUF_X4 buffer423 (.A(\icache.data_mem_data_li [326]),
    .Z(net423));
 BUF_X4 buffer424 (.A(\icache.data_mem_data_li [325]),
    .Z(net424));
 BUF_X4 buffer425 (.A(\icache.data_mem_data_li [324]),
    .Z(net425));
 BUF_X4 buffer426 (.A(\icache.data_mem_data_li [323]),
    .Z(net426));
 BUF_X4 buffer427 (.A(\icache.data_mem_data_li [322]),
    .Z(net427));
 BUF_X4 buffer428 (.A(\icache.data_mem_data_li [321]),
    .Z(net428));
 BUF_X4 buffer429 (.A(\icache.data_mem_data_li [320]),
    .Z(net429));
 BUF_X4 buffer43 (.A(_25501_),
    .Z(net43));
 BUF_X4 buffer430 (.A(\icache.data_mem_data_li [319]),
    .Z(net430));
 BUF_X4 buffer431 (.A(\icache.data_mem_data_li [318]),
    .Z(net431));
 BUF_X4 buffer432 (.A(\icache.data_mem_data_li [317]),
    .Z(net432));
 BUF_X4 buffer433 (.A(\icache.data_mem_data_li [316]),
    .Z(net433));
 BUF_X4 buffer434 (.A(\icache.data_mem_data_li [315]),
    .Z(net434));
 BUF_X4 buffer435 (.A(\icache.data_mem_data_li [314]),
    .Z(net435));
 BUF_X4 buffer436 (.A(\icache.data_mem_data_li [313]),
    .Z(net436));
 BUF_X4 buffer437 (.A(\icache.data_mem_data_li [312]),
    .Z(net437));
 BUF_X4 buffer438 (.A(\icache.data_mem_data_li [311]),
    .Z(net438));
 BUF_X4 buffer439 (.A(\icache.data_mem_data_li [310]),
    .Z(net439));
 BUF_X4 buffer44 (.A(_25095_),
    .Z(net44));
 BUF_X4 buffer440 (.A(\icache.data_mem_data_li [309]),
    .Z(net440));
 BUF_X4 buffer441 (.A(\icache.data_mem_data_li [308]),
    .Z(net441));
 BUF_X4 buffer442 (.A(\icache.data_mem_data_li [307]),
    .Z(net442));
 BUF_X4 buffer443 (.A(\icache.data_mem_data_li [306]),
    .Z(net443));
 BUF_X4 buffer444 (.A(\icache.data_mem_data_li [305]),
    .Z(net444));
 BUF_X4 buffer445 (.A(\icache.data_mem_data_li [304]),
    .Z(net445));
 BUF_X4 buffer446 (.A(\icache.data_mem_data_li [303]),
    .Z(net446));
 BUF_X4 buffer447 (.A(\icache.data_mem_data_li [302]),
    .Z(net447));
 BUF_X4 buffer448 (.A(\icache.data_mem_data_li [301]),
    .Z(net448));
 BUF_X4 buffer449 (.A(\icache.data_mem_data_li [300]),
    .Z(net449));
 BUF_X4 buffer45 (.A(_24954_),
    .Z(net45));
 BUF_X4 buffer450 (.A(\icache.data_mem_data_li [299]),
    .Z(net450));
 BUF_X4 buffer451 (.A(\icache.data_mem_data_li [298]),
    .Z(net451));
 BUF_X4 buffer452 (.A(\icache.data_mem_data_li [297]),
    .Z(net452));
 BUF_X4 buffer453 (.A(\icache.data_mem_data_li [296]),
    .Z(net453));
 BUF_X4 buffer454 (.A(\icache.data_mem_data_li [295]),
    .Z(net454));
 BUF_X4 buffer455 (.A(\icache.data_mem_data_li [294]),
    .Z(net455));
 BUF_X4 buffer456 (.A(\icache.data_mem_data_li [293]),
    .Z(net456));
 BUF_X4 buffer457 (.A(\icache.data_mem_data_li [292]),
    .Z(net457));
 BUF_X4 buffer458 (.A(\icache.data_mem_data_li [291]),
    .Z(net458));
 BUF_X4 buffer459 (.A(\icache.data_mem_data_li [290]),
    .Z(net459));
 BUF_X4 buffer46 (.A(_24950_),
    .Z(net46));
 BUF_X4 buffer460 (.A(\icache.data_mem_data_li [289]),
    .Z(net460));
 BUF_X4 buffer461 (.A(\icache.data_mem_data_li [288]),
    .Z(net461));
 BUF_X4 buffer462 (.A(\icache.data_mem_data_li [287]),
    .Z(net462));
 BUF_X4 buffer463 (.A(\icache.data_mem_data_li [286]),
    .Z(net463));
 BUF_X4 buffer464 (.A(\icache.data_mem_data_li [285]),
    .Z(net464));
 BUF_X4 buffer465 (.A(\icache.data_mem_data_li [284]),
    .Z(net465));
 BUF_X4 buffer466 (.A(\icache.data_mem_data_li [283]),
    .Z(net466));
 BUF_X4 buffer467 (.A(\icache.data_mem_data_li [282]),
    .Z(net467));
 BUF_X4 buffer468 (.A(\icache.data_mem_data_li [281]),
    .Z(net468));
 BUF_X4 buffer469 (.A(\icache.data_mem_data_li [280]),
    .Z(net469));
 BUF_X4 buffer47 (.A(_24784_),
    .Z(net47));
 BUF_X4 buffer470 (.A(\icache.data_mem_data_li [279]),
    .Z(net470));
 BUF_X4 buffer471 (.A(\icache.data_mem_data_li [278]),
    .Z(net471));
 BUF_X4 buffer472 (.A(\icache.data_mem_data_li [277]),
    .Z(net472));
 BUF_X4 buffer473 (.A(\icache.data_mem_data_li [276]),
    .Z(net473));
 BUF_X4 buffer474 (.A(\icache.data_mem_data_li [275]),
    .Z(net474));
 BUF_X4 buffer475 (.A(\icache.data_mem_data_li [274]),
    .Z(net475));
 BUF_X4 buffer476 (.A(\icache.data_mem_data_li [273]),
    .Z(net476));
 BUF_X4 buffer477 (.A(\icache.data_mem_data_li [272]),
    .Z(net477));
 BUF_X4 buffer478 (.A(\icache.data_mem_data_li [271]),
    .Z(net478));
 BUF_X4 buffer479 (.A(\icache.data_mem_data_li [270]),
    .Z(net479));
 BUF_X4 buffer48 (.A(_24577_),
    .Z(net48));
 BUF_X4 buffer480 (.A(\icache.data_mem_data_li [269]),
    .Z(net480));
 BUF_X4 buffer481 (.A(\icache.data_mem_data_li [268]),
    .Z(net481));
 BUF_X4 buffer482 (.A(\icache.data_mem_data_li [267]),
    .Z(net482));
 BUF_X4 buffer483 (.A(\icache.data_mem_data_li [266]),
    .Z(net483));
 BUF_X4 buffer484 (.A(\icache.data_mem_data_li [265]),
    .Z(net484));
 BUF_X4 buffer485 (.A(\icache.data_mem_data_li [264]),
    .Z(net485));
 BUF_X4 buffer486 (.A(\icache.data_mem_data_li [263]),
    .Z(net486));
 BUF_X4 buffer487 (.A(\icache.data_mem_data_li [262]),
    .Z(net487));
 BUF_X4 buffer488 (.A(\icache.data_mem_data_li [261]),
    .Z(net488));
 BUF_X4 buffer489 (.A(\icache.data_mem_data_li [260]),
    .Z(net489));
 BUF_X4 buffer49 (.A(_24532_),
    .Z(net49));
 BUF_X4 buffer490 (.A(\icache.data_mem_data_li [259]),
    .Z(net490));
 BUF_X4 buffer491 (.A(\icache.data_mem_data_li [258]),
    .Z(net491));
 BUF_X4 buffer492 (.A(\icache.data_mem_data_li [257]),
    .Z(net492));
 BUF_X4 buffer493 (.A(\icache.data_mem_data_li [256]),
    .Z(net493));
 BUF_X4 buffer494 (.A(\icache.data_mem_data_li [255]),
    .Z(net494));
 BUF_X4 buffer495 (.A(\icache.data_mem_data_li [254]),
    .Z(net495));
 BUF_X4 buffer496 (.A(\icache.data_mem_data_li [253]),
    .Z(net496));
 BUF_X4 buffer497 (.A(\icache.data_mem_data_li [252]),
    .Z(net497));
 BUF_X4 buffer498 (.A(\icache.data_mem_data_li [251]),
    .Z(net498));
 BUF_X4 buffer499 (.A(\icache.data_mem_data_li [250]),
    .Z(net499));
 BUF_X4 buffer5 (.A(_26279_),
    .Z(net5));
 BUF_X4 buffer50 (.A(_24292_),
    .Z(net50));
 BUF_X4 buffer500 (.A(\icache.data_mem_data_li [249]),
    .Z(net500));
 BUF_X4 buffer501 (.A(\icache.data_mem_data_li [248]),
    .Z(net501));
 BUF_X4 buffer502 (.A(\icache.data_mem_data_li [247]),
    .Z(net502));
 BUF_X4 buffer503 (.A(\icache.data_mem_data_li [246]),
    .Z(net503));
 BUF_X4 buffer504 (.A(\icache.data_mem_data_li [245]),
    .Z(net504));
 BUF_X4 buffer505 (.A(\icache.data_mem_data_li [244]),
    .Z(net505));
 BUF_X4 buffer506 (.A(\icache.data_mem_data_li [243]),
    .Z(net506));
 BUF_X4 buffer507 (.A(\icache.data_mem_data_li [242]),
    .Z(net507));
 BUF_X4 buffer508 (.A(\icache.data_mem_data_li [241]),
    .Z(net508));
 BUF_X4 buffer509 (.A(\icache.data_mem_data_li [240]),
    .Z(net509));
 BUF_X4 buffer51 (.A(_24075_),
    .Z(net51));
 BUF_X4 buffer510 (.A(\icache.data_mem_data_li [239]),
    .Z(net510));
 BUF_X4 buffer511 (.A(\icache.data_mem_data_li [238]),
    .Z(net511));
 BUF_X4 buffer512 (.A(\icache.data_mem_data_li [237]),
    .Z(net512));
 BUF_X4 buffer513 (.A(\icache.data_mem_data_li [236]),
    .Z(net513));
 BUF_X4 buffer514 (.A(\icache.data_mem_data_li [235]),
    .Z(net514));
 BUF_X4 buffer515 (.A(\icache.data_mem_data_li [234]),
    .Z(net515));
 BUF_X4 buffer516 (.A(\icache.data_mem_data_li [233]),
    .Z(net516));
 BUF_X4 buffer517 (.A(\icache.data_mem_data_li [232]),
    .Z(net517));
 BUF_X4 buffer518 (.A(\icache.data_mem_data_li [231]),
    .Z(net518));
 BUF_X4 buffer519 (.A(\icache.data_mem_data_li [230]),
    .Z(net519));
 BUF_X4 buffer52 (.A(_23989_),
    .Z(net52));
 BUF_X4 buffer520 (.A(\icache.data_mem_data_li [229]),
    .Z(net520));
 BUF_X4 buffer521 (.A(\icache.data_mem_data_li [228]),
    .Z(net521));
 BUF_X4 buffer522 (.A(\icache.data_mem_data_li [227]),
    .Z(net522));
 BUF_X4 buffer523 (.A(\icache.data_mem_data_li [226]),
    .Z(net523));
 BUF_X4 buffer524 (.A(\icache.data_mem_data_li [225]),
    .Z(net524));
 BUF_X4 buffer525 (.A(\icache.data_mem_data_li [224]),
    .Z(net525));
 BUF_X4 buffer526 (.A(\icache.data_mem_data_li [223]),
    .Z(net526));
 BUF_X4 buffer527 (.A(\icache.data_mem_data_li [222]),
    .Z(net527));
 BUF_X4 buffer528 (.A(\icache.data_mem_data_li [221]),
    .Z(net528));
 BUF_X4 buffer529 (.A(\icache.data_mem_data_li [220]),
    .Z(net529));
 BUF_X4 buffer53 (.A(_23650_),
    .Z(net53));
 BUF_X4 buffer530 (.A(\icache.data_mem_data_li [219]),
    .Z(net530));
 BUF_X4 buffer531 (.A(\icache.data_mem_data_li [218]),
    .Z(net531));
 BUF_X4 buffer532 (.A(\icache.data_mem_data_li [217]),
    .Z(net532));
 BUF_X4 buffer533 (.A(\icache.data_mem_data_li [216]),
    .Z(net533));
 BUF_X4 buffer534 (.A(\icache.data_mem_data_li [215]),
    .Z(net534));
 BUF_X4 buffer535 (.A(\icache.data_mem_data_li [214]),
    .Z(net535));
 BUF_X4 buffer536 (.A(\icache.data_mem_data_li [213]),
    .Z(net536));
 BUF_X4 buffer537 (.A(\icache.data_mem_data_li [212]),
    .Z(net537));
 BUF_X4 buffer538 (.A(\icache.data_mem_data_li [211]),
    .Z(net538));
 BUF_X4 buffer539 (.A(\icache.data_mem_data_li [210]),
    .Z(net539));
 BUF_X4 buffer54 (.A(_23462_),
    .Z(net54));
 BUF_X4 buffer540 (.A(\icache.data_mem_data_li [209]),
    .Z(net540));
 BUF_X4 buffer541 (.A(\icache.data_mem_data_li [208]),
    .Z(net541));
 BUF_X4 buffer542 (.A(\icache.data_mem_data_li [207]),
    .Z(net542));
 BUF_X4 buffer543 (.A(\icache.data_mem_data_li [206]),
    .Z(net543));
 BUF_X4 buffer544 (.A(\icache.data_mem_data_li [205]),
    .Z(net544));
 BUF_X4 buffer545 (.A(\icache.data_mem_data_li [204]),
    .Z(net545));
 BUF_X4 buffer546 (.A(\icache.data_mem_data_li [203]),
    .Z(net546));
 BUF_X4 buffer547 (.A(\icache.data_mem_data_li [202]),
    .Z(net547));
 BUF_X4 buffer548 (.A(\icache.data_mem_data_li [201]),
    .Z(net548));
 BUF_X4 buffer549 (.A(\icache.data_mem_data_li [200]),
    .Z(net549));
 BUF_X4 buffer55 (.A(_23287_),
    .Z(net55));
 BUF_X4 buffer550 (.A(\icache.data_mem_data_li [199]),
    .Z(net550));
 BUF_X4 buffer551 (.A(\icache.data_mem_data_li [198]),
    .Z(net551));
 BUF_X4 buffer552 (.A(\icache.data_mem_data_li [197]),
    .Z(net552));
 BUF_X4 buffer553 (.A(\icache.data_mem_data_li [196]),
    .Z(net553));
 BUF_X4 buffer554 (.A(\icache.data_mem_data_li [195]),
    .Z(net554));
 BUF_X4 buffer555 (.A(\icache.data_mem_data_li [194]),
    .Z(net555));
 BUF_X4 buffer556 (.A(\icache.data_mem_data_li [193]),
    .Z(net556));
 BUF_X4 buffer557 (.A(\icache.data_mem_data_li [192]),
    .Z(net557));
 BUF_X4 buffer558 (.A(\icache.data_mem_data_li [191]),
    .Z(net558));
 BUF_X4 buffer559 (.A(\icache.data_mem_data_li [190]),
    .Z(net559));
 BUF_X4 buffer56 (.A(_23105_),
    .Z(net56));
 BUF_X4 buffer560 (.A(\icache.data_mem_data_li [189]),
    .Z(net560));
 BUF_X4 buffer561 (.A(\icache.data_mem_data_li [188]),
    .Z(net561));
 BUF_X4 buffer562 (.A(\icache.data_mem_data_li [187]),
    .Z(net562));
 BUF_X4 buffer563 (.A(\icache.data_mem_data_li [186]),
    .Z(net563));
 BUF_X4 buffer564 (.A(\icache.data_mem_data_li [185]),
    .Z(net564));
 BUF_X4 buffer565 (.A(\icache.data_mem_data_li [184]),
    .Z(net565));
 BUF_X4 buffer566 (.A(\icache.data_mem_data_li [183]),
    .Z(net566));
 BUF_X4 buffer567 (.A(\icache.data_mem_data_li [182]),
    .Z(net567));
 BUF_X4 buffer568 (.A(\icache.data_mem_data_li [181]),
    .Z(net568));
 BUF_X4 buffer569 (.A(\icache.data_mem_data_li [180]),
    .Z(net569));
 BUF_X4 buffer57 (.A(_26190_),
    .Z(net57));
 BUF_X4 buffer570 (.A(\icache.data_mem_data_li [179]),
    .Z(net570));
 BUF_X4 buffer571 (.A(\icache.data_mem_data_li [178]),
    .Z(net571));
 BUF_X4 buffer572 (.A(\icache.data_mem_data_li [177]),
    .Z(net572));
 BUF_X4 buffer573 (.A(\icache.data_mem_data_li [176]),
    .Z(net573));
 BUF_X4 buffer574 (.A(\icache.data_mem_data_li [175]),
    .Z(net574));
 BUF_X4 buffer575 (.A(\icache.data_mem_data_li [174]),
    .Z(net575));
 BUF_X4 buffer576 (.A(\icache.data_mem_data_li [173]),
    .Z(net576));
 BUF_X4 buffer577 (.A(\icache.data_mem_data_li [172]),
    .Z(net577));
 BUF_X4 buffer578 (.A(\icache.data_mem_data_li [171]),
    .Z(net578));
 BUF_X4 buffer579 (.A(\icache.data_mem_data_li [170]),
    .Z(net579));
 BUF_X4 buffer58 (.A(_25377_),
    .Z(net58));
 BUF_X4 buffer580 (.A(\icache.data_mem_data_li [169]),
    .Z(net580));
 BUF_X4 buffer581 (.A(\icache.data_mem_data_li [168]),
    .Z(net581));
 BUF_X4 buffer582 (.A(\icache.data_mem_data_li [167]),
    .Z(net582));
 BUF_X4 buffer583 (.A(\icache.data_mem_data_li [166]),
    .Z(net583));
 BUF_X4 buffer584 (.A(\icache.data_mem_data_li [165]),
    .Z(net584));
 BUF_X4 buffer585 (.A(\icache.data_mem_data_li [164]),
    .Z(net585));
 BUF_X4 buffer586 (.A(\icache.data_mem_data_li [163]),
    .Z(net586));
 BUF_X4 buffer587 (.A(\icache.data_mem_data_li [162]),
    .Z(net587));
 BUF_X4 buffer588 (.A(\icache.data_mem_data_li [161]),
    .Z(net588));
 BUF_X4 buffer589 (.A(\icache.data_mem_data_li [160]),
    .Z(net589));
 BUF_X4 buffer59 (.A(_24249_),
    .Z(net59));
 BUF_X4 buffer590 (.A(\icache.data_mem_data_li [159]),
    .Z(net590));
 BUF_X4 buffer591 (.A(\icache.data_mem_data_li [158]),
    .Z(net591));
 BUF_X4 buffer592 (.A(\icache.data_mem_data_li [157]),
    .Z(net592));
 BUF_X4 buffer593 (.A(\icache.data_mem_data_li [156]),
    .Z(net593));
 BUF_X4 buffer594 (.A(\icache.data_mem_data_li [155]),
    .Z(net594));
 BUF_X4 buffer595 (.A(\icache.data_mem_data_li [154]),
    .Z(net595));
 BUF_X4 buffer596 (.A(\icache.data_mem_data_li [153]),
    .Z(net596));
 BUF_X4 buffer597 (.A(\icache.data_mem_data_li [152]),
    .Z(net597));
 BUF_X4 buffer598 (.A(\icache.data_mem_data_li [151]),
    .Z(net598));
 BUF_X4 buffer599 (.A(\icache.data_mem_data_li [150]),
    .Z(net599));
 BUF_X4 buffer6 (.A(_26251_),
    .Z(net6));
 BUF_X4 buffer60 (.A(_10872_),
    .Z(net60));
 BUF_X4 buffer600 (.A(\icache.data_mem_data_li [149]),
    .Z(net600));
 BUF_X4 buffer601 (.A(\icache.data_mem_data_li [148]),
    .Z(net601));
 BUF_X4 buffer602 (.A(\icache.data_mem_data_li [147]),
    .Z(net602));
 BUF_X4 buffer603 (.A(\icache.data_mem_data_li [146]),
    .Z(net603));
 BUF_X4 buffer604 (.A(\icache.data_mem_data_li [145]),
    .Z(net604));
 BUF_X4 buffer605 (.A(\icache.data_mem_data_li [144]),
    .Z(net605));
 BUF_X4 buffer606 (.A(\icache.data_mem_data_li [143]),
    .Z(net606));
 BUF_X4 buffer607 (.A(\icache.data_mem_data_li [142]),
    .Z(net607));
 BUF_X4 buffer608 (.A(\icache.data_mem_data_li [141]),
    .Z(net608));
 BUF_X4 buffer609 (.A(\icache.data_mem_data_li [140]),
    .Z(net609));
 BUF_X4 buffer61 (.A(net60),
    .Z(net61));
 BUF_X4 buffer610 (.A(\icache.data_mem_data_li [139]),
    .Z(net610));
 BUF_X4 buffer611 (.A(\icache.data_mem_data_li [138]),
    .Z(net611));
 BUF_X4 buffer612 (.A(\icache.data_mem_data_li [137]),
    .Z(net612));
 BUF_X4 buffer613 (.A(\icache.data_mem_data_li [136]),
    .Z(net613));
 BUF_X4 buffer614 (.A(\icache.data_mem_data_li [135]),
    .Z(net614));
 BUF_X4 buffer615 (.A(\icache.data_mem_data_li [134]),
    .Z(net615));
 BUF_X4 buffer616 (.A(\icache.data_mem_data_li [133]),
    .Z(net616));
 BUF_X4 buffer617 (.A(\icache.data_mem_data_li [132]),
    .Z(net617));
 BUF_X4 buffer618 (.A(\icache.data_mem_data_li [131]),
    .Z(net618));
 BUF_X4 buffer619 (.A(\icache.data_mem_data_li [130]),
    .Z(net619));
 BUF_X4 buffer62 (.A(net60),
    .Z(net62));
 BUF_X4 buffer620 (.A(\icache.data_mem_data_li [129]),
    .Z(net620));
 BUF_X4 buffer621 (.A(\icache.data_mem_data_li [128]),
    .Z(net621));
 BUF_X4 buffer622 (.A(\icache.data_mem_data_li [127]),
    .Z(net622));
 BUF_X4 buffer623 (.A(\icache.data_mem_data_li [126]),
    .Z(net623));
 BUF_X4 buffer624 (.A(\icache.data_mem_data_li [125]),
    .Z(net624));
 BUF_X4 buffer625 (.A(\icache.data_mem_data_li [124]),
    .Z(net625));
 BUF_X4 buffer626 (.A(\icache.data_mem_data_li [123]),
    .Z(net626));
 BUF_X4 buffer627 (.A(\icache.data_mem_data_li [122]),
    .Z(net627));
 BUF_X4 buffer628 (.A(\icache.data_mem_data_li [121]),
    .Z(net628));
 BUF_X4 buffer629 (.A(\icache.data_mem_data_li [120]),
    .Z(net629));
 BUF_X4 buffer63 (.A(_10862_),
    .Z(net63));
 BUF_X4 buffer630 (.A(\icache.data_mem_data_li [119]),
    .Z(net630));
 BUF_X4 buffer631 (.A(\icache.data_mem_data_li [118]),
    .Z(net631));
 BUF_X4 buffer632 (.A(\icache.data_mem_data_li [117]),
    .Z(net632));
 BUF_X4 buffer633 (.A(\icache.data_mem_data_li [116]),
    .Z(net633));
 BUF_X4 buffer634 (.A(\icache.data_mem_data_li [115]),
    .Z(net634));
 BUF_X4 buffer635 (.A(\icache.data_mem_data_li [114]),
    .Z(net635));
 BUF_X4 buffer636 (.A(\icache.data_mem_data_li [113]),
    .Z(net636));
 BUF_X4 buffer637 (.A(\icache.data_mem_data_li [112]),
    .Z(net637));
 BUF_X4 buffer638 (.A(\icache.data_mem_data_li [111]),
    .Z(net638));
 BUF_X4 buffer639 (.A(\icache.data_mem_data_li [110]),
    .Z(net639));
 BUF_X4 buffer64 (.A(net63),
    .Z(net64));
 BUF_X4 buffer640 (.A(\icache.data_mem_data_li [109]),
    .Z(net640));
 BUF_X4 buffer641 (.A(\icache.data_mem_data_li [108]),
    .Z(net641));
 BUF_X4 buffer642 (.A(\icache.data_mem_data_li [107]),
    .Z(net642));
 BUF_X4 buffer643 (.A(\icache.data_mem_data_li [106]),
    .Z(net643));
 BUF_X4 buffer644 (.A(\icache.data_mem_data_li [105]),
    .Z(net644));
 BUF_X4 buffer645 (.A(\icache.data_mem_data_li [104]),
    .Z(net645));
 BUF_X4 buffer646 (.A(\icache.data_mem_data_li [103]),
    .Z(net646));
 BUF_X4 buffer647 (.A(\icache.data_mem_data_li [102]),
    .Z(net647));
 BUF_X4 buffer648 (.A(\icache.data_mem_data_li [101]),
    .Z(net648));
 BUF_X4 buffer649 (.A(\icache.data_mem_data_li [100]),
    .Z(net649));
 BUF_X4 buffer65 (.A(net63),
    .Z(net65));
 BUF_X4 buffer650 (.A(\icache.data_mem_data_li [99]),
    .Z(net650));
 BUF_X4 buffer651 (.A(\icache.data_mem_data_li [98]),
    .Z(net651));
 BUF_X4 buffer652 (.A(\icache.data_mem_data_li [97]),
    .Z(net652));
 BUF_X4 buffer653 (.A(\icache.data_mem_data_li [96]),
    .Z(net653));
 BUF_X4 buffer654 (.A(\icache.data_mem_data_li [95]),
    .Z(net654));
 BUF_X4 buffer655 (.A(\icache.data_mem_data_li [94]),
    .Z(net655));
 BUF_X4 buffer656 (.A(\icache.data_mem_data_li [93]),
    .Z(net656));
 BUF_X4 buffer657 (.A(\icache.data_mem_data_li [92]),
    .Z(net657));
 BUF_X4 buffer658 (.A(\icache.data_mem_data_li [91]),
    .Z(net658));
 BUF_X4 buffer659 (.A(\icache.data_mem_data_li [90]),
    .Z(net659));
 BUF_X4 buffer66 (.A(_10862_),
    .Z(net66));
 BUF_X4 buffer660 (.A(\icache.data_mem_data_li [89]),
    .Z(net660));
 BUF_X4 buffer661 (.A(\icache.data_mem_data_li [88]),
    .Z(net661));
 BUF_X4 buffer662 (.A(\icache.data_mem_data_li [87]),
    .Z(net662));
 BUF_X4 buffer663 (.A(\icache.data_mem_data_li [86]),
    .Z(net663));
 BUF_X4 buffer664 (.A(\icache.data_mem_data_li [85]),
    .Z(net664));
 BUF_X4 buffer665 (.A(\icache.data_mem_data_li [84]),
    .Z(net665));
 BUF_X4 buffer666 (.A(\icache.data_mem_data_li [83]),
    .Z(net666));
 BUF_X4 buffer667 (.A(\icache.data_mem_data_li [82]),
    .Z(net667));
 BUF_X4 buffer668 (.A(\icache.data_mem_data_li [81]),
    .Z(net668));
 BUF_X4 buffer669 (.A(\icache.data_mem_data_li [80]),
    .Z(net669));
 BUF_X4 buffer67 (.A(net66),
    .Z(net67));
 BUF_X4 buffer670 (.A(\icache.data_mem_data_li [79]),
    .Z(net670));
 BUF_X4 buffer671 (.A(\icache.data_mem_data_li [78]),
    .Z(net671));
 BUF_X4 buffer672 (.A(\icache.data_mem_data_li [77]),
    .Z(net672));
 BUF_X4 buffer673 (.A(\icache.data_mem_data_li [76]),
    .Z(net673));
 BUF_X4 buffer674 (.A(\icache.data_mem_data_li [75]),
    .Z(net674));
 BUF_X4 buffer675 (.A(\icache.data_mem_data_li [74]),
    .Z(net675));
 BUF_X4 buffer676 (.A(\icache.data_mem_data_li [73]),
    .Z(net676));
 BUF_X4 buffer677 (.A(\icache.data_mem_data_li [72]),
    .Z(net677));
 BUF_X4 buffer678 (.A(\icache.data_mem_data_li [71]),
    .Z(net678));
 BUF_X4 buffer679 (.A(\icache.data_mem_data_li [70]),
    .Z(net679));
 BUF_X4 buffer68 (.A(net66),
    .Z(net68));
 BUF_X4 buffer680 (.A(\icache.data_mem_data_li [69]),
    .Z(net680));
 BUF_X4 buffer681 (.A(\icache.data_mem_data_li [68]),
    .Z(net681));
 BUF_X4 buffer682 (.A(\icache.data_mem_data_li [67]),
    .Z(net682));
 BUF_X4 buffer683 (.A(\icache.data_mem_data_li [66]),
    .Z(net683));
 BUF_X4 buffer684 (.A(\icache.data_mem_data_li [65]),
    .Z(net684));
 BUF_X4 buffer685 (.A(\icache.data_mem_data_li [64]),
    .Z(net685));
 BUF_X4 buffer686 (.A(\icache.data_mem_data_li [63]),
    .Z(net686));
 BUF_X4 buffer687 (.A(\icache.data_mem_data_li [62]),
    .Z(net687));
 BUF_X4 buffer688 (.A(\icache.data_mem_data_li [61]),
    .Z(net688));
 BUF_X4 buffer689 (.A(\icache.data_mem_data_li [60]),
    .Z(net689));
 BUF_X4 buffer69 (.A(_10837_),
    .Z(net69));
 BUF_X4 buffer690 (.A(\icache.data_mem_data_li [59]),
    .Z(net690));
 BUF_X4 buffer691 (.A(\icache.data_mem_data_li [58]),
    .Z(net691));
 BUF_X4 buffer692 (.A(\icache.data_mem_data_li [57]),
    .Z(net692));
 BUF_X4 buffer693 (.A(\icache.data_mem_data_li [56]),
    .Z(net693));
 BUF_X4 buffer694 (.A(\icache.data_mem_data_li [55]),
    .Z(net694));
 BUF_X4 buffer695 (.A(\icache.data_mem_data_li [54]),
    .Z(net695));
 BUF_X4 buffer696 (.A(\icache.data_mem_data_li [53]),
    .Z(net696));
 BUF_X4 buffer697 (.A(\icache.data_mem_data_li [52]),
    .Z(net697));
 BUF_X4 buffer698 (.A(\icache.data_mem_data_li [51]),
    .Z(net698));
 BUF_X4 buffer699 (.A(\icache.data_mem_data_li [50]),
    .Z(net699));
 BUF_X4 buffer7 (.A(_25020_),
    .Z(net7));
 BUF_X4 buffer70 (.A(net69),
    .Z(net70));
 BUF_X4 buffer700 (.A(\icache.data_mem_data_li [49]),
    .Z(net700));
 BUF_X4 buffer701 (.A(\icache.data_mem_data_li [48]),
    .Z(net701));
 BUF_X4 buffer702 (.A(\icache.data_mem_data_li [47]),
    .Z(net702));
 BUF_X4 buffer703 (.A(\icache.data_mem_data_li [46]),
    .Z(net703));
 BUF_X4 buffer704 (.A(\icache.data_mem_data_li [45]),
    .Z(net704));
 BUF_X4 buffer705 (.A(\icache.data_mem_data_li [44]),
    .Z(net705));
 BUF_X4 buffer706 (.A(\icache.data_mem_data_li [43]),
    .Z(net706));
 BUF_X4 buffer707 (.A(\icache.data_mem_data_li [42]),
    .Z(net707));
 BUF_X4 buffer708 (.A(\icache.data_mem_data_li [41]),
    .Z(net708));
 BUF_X4 buffer709 (.A(\icache.data_mem_data_li [40]),
    .Z(net709));
 BUF_X4 buffer71 (.A(net69),
    .Z(net71));
 BUF_X4 buffer710 (.A(\icache.data_mem_data_li [39]),
    .Z(net710));
 BUF_X4 buffer711 (.A(\icache.data_mem_data_li [38]),
    .Z(net711));
 BUF_X4 buffer712 (.A(\icache.data_mem_data_li [37]),
    .Z(net712));
 BUF_X4 buffer713 (.A(\icache.data_mem_data_li [36]),
    .Z(net713));
 BUF_X4 buffer714 (.A(\icache.data_mem_data_li [35]),
    .Z(net714));
 BUF_X4 buffer715 (.A(\icache.data_mem_data_li [34]),
    .Z(net715));
 BUF_X4 buffer716 (.A(\icache.data_mem_data_li [33]),
    .Z(net716));
 BUF_X4 buffer717 (.A(\icache.data_mem_data_li [32]),
    .Z(net717));
 BUF_X4 buffer718 (.A(\icache.data_mem_data_li [31]),
    .Z(net718));
 BUF_X4 buffer719 (.A(\icache.data_mem_data_li [30]),
    .Z(net719));
 BUF_X4 buffer72 (.A(net69),
    .Z(net72));
 BUF_X4 buffer720 (.A(\icache.data_mem_data_li [29]),
    .Z(net720));
 BUF_X4 buffer721 (.A(\icache.data_mem_data_li [28]),
    .Z(net721));
 BUF_X4 buffer722 (.A(\icache.data_mem_data_li [27]),
    .Z(net722));
 BUF_X4 buffer723 (.A(\icache.data_mem_data_li [26]),
    .Z(net723));
 BUF_X4 buffer724 (.A(\icache.data_mem_data_li [25]),
    .Z(net724));
 BUF_X4 buffer725 (.A(\icache.data_mem_data_li [24]),
    .Z(net725));
 BUF_X4 buffer726 (.A(\icache.data_mem_data_li [23]),
    .Z(net726));
 BUF_X4 buffer727 (.A(\icache.data_mem_data_li [22]),
    .Z(net727));
 BUF_X4 buffer728 (.A(\icache.data_mem_data_li [21]),
    .Z(net728));
 BUF_X4 buffer729 (.A(\icache.data_mem_data_li [20]),
    .Z(net729));
 BUF_X4 buffer73 (.A(net69),
    .Z(net73));
 BUF_X4 buffer730 (.A(\icache.data_mem_data_li [19]),
    .Z(net730));
 BUF_X4 buffer731 (.A(\icache.data_mem_data_li [18]),
    .Z(net731));
 BUF_X4 buffer732 (.A(\icache.data_mem_data_li [17]),
    .Z(net732));
 BUF_X4 buffer733 (.A(\icache.data_mem_data_li [16]),
    .Z(net733));
 BUF_X4 buffer734 (.A(\icache.data_mem_data_li [15]),
    .Z(net734));
 BUF_X4 buffer735 (.A(\icache.data_mem_data_li [14]),
    .Z(net735));
 BUF_X4 buffer736 (.A(\icache.data_mem_data_li [13]),
    .Z(net736));
 BUF_X4 buffer737 (.A(\icache.data_mem_data_li [12]),
    .Z(net737));
 BUF_X4 buffer738 (.A(\icache.data_mem_data_li [11]),
    .Z(net738));
 BUF_X4 buffer739 (.A(\icache.data_mem_data_li [10]),
    .Z(net739));
 BUF_X4 buffer74 (.A(net69),
    .Z(net74));
 BUF_X4 buffer740 (.A(\icache.data_mem_data_li [9]),
    .Z(net740));
 BUF_X4 buffer741 (.A(\icache.data_mem_data_li [8]),
    .Z(net741));
 BUF_X4 buffer742 (.A(\icache.data_mem_data_li [7]),
    .Z(net742));
 BUF_X4 buffer743 (.A(\icache.data_mem_data_li [6]),
    .Z(net743));
 BUF_X4 buffer744 (.A(\icache.data_mem_data_li [5]),
    .Z(net744));
 BUF_X4 buffer745 (.A(\icache.data_mem_data_li [4]),
    .Z(net745));
 BUF_X4 buffer746 (.A(\icache.data_mem_data_li [3]),
    .Z(net746));
 BUF_X4 buffer747 (.A(\icache.data_mem_data_li [2]),
    .Z(net747));
 BUF_X4 buffer748 (.A(\icache.data_mem_data_li [1]),
    .Z(net748));
 BUF_X4 buffer749 (.A(\icache.data_mem_data_li [0]),
    .Z(net749));
 BUF_X4 buffer75 (.A(net74),
    .Z(net75));
 BUF_X4 buffer750 (.A(\icache.tag_mem.w_mask_i [143]),
    .Z(net750));
 BUF_X4 buffer751 (.A(\icache.tag_mem.w_mask_i [143]),
    .Z(net751));
 BUF_X4 buffer752 (.A(\icache.tag_mem.w_mask_i [116]),
    .Z(net752));
 BUF_X4 buffer753 (.A(net752),
    .Z(net753));
 BUF_X4 buffer754 (.A(net752),
    .Z(net754));
 BUF_X4 buffer755 (.A(net752),
    .Z(net755));
 BUF_X4 buffer756 (.A(net752),
    .Z(net756));
 BUF_X4 buffer757 (.A(net752),
    .Z(net757));
 BUF_X4 buffer758 (.A(net752),
    .Z(net758));
 BUF_X4 buffer759 (.A(net752),
    .Z(net759));
 BUF_X4 buffer76 (.A(net74),
    .Z(net76));
 BUF_X4 buffer760 (.A(net752),
    .Z(net760));
 BUF_X4 buffer761 (.A(net752),
    .Z(net761));
 BUF_X4 buffer762 (.A(net752),
    .Z(net762));
 BUF_X4 buffer763 (.A(net752),
    .Z(net763));
 BUF_X4 buffer764 (.A(net752),
    .Z(net764));
 BUF_X4 buffer765 (.A(net752),
    .Z(net765));
 BUF_X4 buffer766 (.A(net752),
    .Z(net766));
 BUF_X4 buffer767 (.A(net752),
    .Z(net767));
 BUF_X4 buffer768 (.A(net752),
    .Z(net768));
 BUF_X4 buffer769 (.A(net752),
    .Z(net769));
 BUF_X4 buffer77 (.A(_10823_),
    .Z(net77));
 BUF_X4 buffer770 (.A(net752),
    .Z(net770));
 BUF_X4 buffer771 (.A(net752),
    .Z(net771));
 BUF_X4 buffer772 (.A(net752),
    .Z(net772));
 BUF_X4 buffer773 (.A(net752),
    .Z(net773));
 BUF_X4 buffer774 (.A(net752),
    .Z(net774));
 BUF_X4 buffer775 (.A(net752),
    .Z(net775));
 BUF_X4 buffer776 (.A(net752),
    .Z(net776));
 BUF_X4 buffer777 (.A(net752),
    .Z(net777));
 BUF_X4 buffer778 (.A(net752),
    .Z(net778));
 BUF_X4 buffer779 (.A(net752),
    .Z(net779));
 BUF_X4 buffer78 (.A(net77),
    .Z(net78));
 BUF_X4 buffer780 (.A(\icache.tag_mem.w_mask_i [114]),
    .Z(net780));
 BUF_X4 buffer781 (.A(\icache.tag_mem.w_mask_i [114]),
    .Z(net781));
 BUF_X4 buffer782 (.A(\icache.tag_mem.w_mask_i [100]),
    .Z(net782));
 BUF_X4 buffer783 (.A(net782),
    .Z(net783));
 BUF_X4 buffer784 (.A(net782),
    .Z(net784));
 BUF_X4 buffer785 (.A(net782),
    .Z(net785));
 BUF_X4 buffer786 (.A(net782),
    .Z(net786));
 BUF_X4 buffer787 (.A(net782),
    .Z(net787));
 BUF_X4 buffer788 (.A(net782),
    .Z(net788));
 BUF_X4 buffer789 (.A(net782),
    .Z(net789));
 BUF_X4 buffer79 (.A(net77),
    .Z(net79));
 BUF_X4 buffer790 (.A(net782),
    .Z(net790));
 BUF_X4 buffer791 (.A(net782),
    .Z(net791));
 BUF_X4 buffer792 (.A(net782),
    .Z(net792));
 BUF_X4 buffer793 (.A(net782),
    .Z(net793));
 BUF_X4 buffer794 (.A(net782),
    .Z(net794));
 BUF_X4 buffer795 (.A(net782),
    .Z(net795));
 BUF_X4 buffer796 (.A(net782),
    .Z(net796));
 BUF_X4 buffer797 (.A(net782),
    .Z(net797));
 BUF_X4 buffer798 (.A(net782),
    .Z(net798));
 BUF_X4 buffer799 (.A(net782),
    .Z(net799));
 BUF_X4 buffer8 (.A(_24964_),
    .Z(net8));
 BUF_X4 buffer80 (.A(net79),
    .Z(net80));
 BUF_X4 buffer800 (.A(net782),
    .Z(net800));
 BUF_X4 buffer801 (.A(net782),
    .Z(net801));
 BUF_X4 buffer802 (.A(net782),
    .Z(net802));
 BUF_X4 buffer803 (.A(net782),
    .Z(net803));
 BUF_X4 buffer804 (.A(net782),
    .Z(net804));
 BUF_X4 buffer805 (.A(net782),
    .Z(net805));
 BUF_X4 buffer806 (.A(net782),
    .Z(net806));
 BUF_X4 buffer807 (.A(net782),
    .Z(net807));
 BUF_X4 buffer808 (.A(net782),
    .Z(net808));
 BUF_X4 buffer809 (.A(net782),
    .Z(net809));
 BUF_X4 buffer81 (.A(net77),
    .Z(net81));
 BUF_X4 buffer810 (.A(\icache.tag_mem.w_mask_i [85]),
    .Z(net810));
 BUF_X4 buffer811 (.A(\icache.tag_mem.w_mask_i [85]),
    .Z(net811));
 BUF_X4 buffer812 (.A(\icache.tag_mem.w_mask_i [58]),
    .Z(net812));
 BUF_X4 buffer813 (.A(net812),
    .Z(net813));
 BUF_X4 buffer814 (.A(net812),
    .Z(net814));
 BUF_X4 buffer815 (.A(net812),
    .Z(net815));
 BUF_X4 buffer816 (.A(net812),
    .Z(net816));
 BUF_X4 buffer817 (.A(net812),
    .Z(net817));
 BUF_X4 buffer818 (.A(net812),
    .Z(net818));
 BUF_X4 buffer819 (.A(net812),
    .Z(net819));
 BUF_X4 buffer82 (.A(net81),
    .Z(net82));
 BUF_X4 buffer820 (.A(net812),
    .Z(net820));
 BUF_X4 buffer821 (.A(net812),
    .Z(net821));
 BUF_X4 buffer822 (.A(net812),
    .Z(net822));
 BUF_X4 buffer823 (.A(net812),
    .Z(net823));
 BUF_X4 buffer824 (.A(net812),
    .Z(net824));
 BUF_X4 buffer825 (.A(net812),
    .Z(net825));
 BUF_X4 buffer826 (.A(net812),
    .Z(net826));
 BUF_X4 buffer827 (.A(net812),
    .Z(net827));
 BUF_X4 buffer828 (.A(net812),
    .Z(net828));
 BUF_X4 buffer829 (.A(net812),
    .Z(net829));
 BUF_X4 buffer83 (.A(_10810_),
    .Z(net83));
 BUF_X4 buffer830 (.A(net812),
    .Z(net830));
 BUF_X4 buffer831 (.A(net812),
    .Z(net831));
 BUF_X4 buffer832 (.A(net812),
    .Z(net832));
 BUF_X4 buffer833 (.A(net812),
    .Z(net833));
 BUF_X4 buffer834 (.A(net812),
    .Z(net834));
 BUF_X4 buffer835 (.A(net812),
    .Z(net835));
 BUF_X4 buffer836 (.A(net812),
    .Z(net836));
 BUF_X4 buffer837 (.A(net812),
    .Z(net837));
 BUF_X4 buffer838 (.A(net812),
    .Z(net838));
 BUF_X4 buffer839 (.A(net812),
    .Z(net839));
 BUF_X4 buffer84 (.A(_10810_),
    .Z(net84));
 BUF_X4 buffer840 (.A(\icache.tag_mem.w_mask_i [56]),
    .Z(net840));
 BUF_X4 buffer841 (.A(\icache.tag_mem.w_mask_i [56]),
    .Z(net841));
 BUF_X4 buffer842 (.A(\icache.tag_mem.w_mask_i [29]),
    .Z(net842));
 BUF_X4 buffer843 (.A(net842),
    .Z(net843));
 BUF_X4 buffer844 (.A(net842),
    .Z(net844));
 BUF_X4 buffer845 (.A(net842),
    .Z(net845));
 BUF_X4 buffer846 (.A(net842),
    .Z(net846));
 BUF_X4 buffer847 (.A(net842),
    .Z(net847));
 BUF_X4 buffer848 (.A(net842),
    .Z(net848));
 BUF_X4 buffer849 (.A(net842),
    .Z(net849));
 BUF_X4 buffer85 (.A(_10810_),
    .Z(net85));
 BUF_X4 buffer850 (.A(net842),
    .Z(net850));
 BUF_X4 buffer851 (.A(net842),
    .Z(net851));
 BUF_X4 buffer852 (.A(net842),
    .Z(net852));
 BUF_X4 buffer853 (.A(net842),
    .Z(net853));
 BUF_X4 buffer854 (.A(net842),
    .Z(net854));
 BUF_X4 buffer855 (.A(net842),
    .Z(net855));
 BUF_X4 buffer856 (.A(net842),
    .Z(net856));
 BUF_X4 buffer857 (.A(net842),
    .Z(net857));
 BUF_X4 buffer858 (.A(net842),
    .Z(net858));
 BUF_X4 buffer859 (.A(net842),
    .Z(net859));
 BUF_X4 buffer86 (.A(_10810_),
    .Z(net86));
 BUF_X4 buffer860 (.A(net842),
    .Z(net860));
 BUF_X4 buffer861 (.A(net842),
    .Z(net861));
 BUF_X4 buffer862 (.A(net842),
    .Z(net862));
 BUF_X4 buffer863 (.A(net842),
    .Z(net863));
 BUF_X4 buffer864 (.A(net842),
    .Z(net864));
 BUF_X4 buffer865 (.A(net842),
    .Z(net865));
 BUF_X4 buffer866 (.A(net842),
    .Z(net866));
 BUF_X4 buffer867 (.A(net842),
    .Z(net867));
 BUF_X4 buffer868 (.A(net842),
    .Z(net868));
 BUF_X4 buffer869 (.A(net842),
    .Z(net869));
 BUF_X4 buffer87 (.A(_10810_),
    .Z(net87));
 BUF_X4 buffer870 (.A(\icache.tag_mem.w_mask_i [0]),
    .Z(net870));
 BUF_X4 buffer871 (.A(net870),
    .Z(net871));
 BUF_X4 buffer872 (.A(net870),
    .Z(net872));
 BUF_X4 buffer873 (.A(net870),
    .Z(net873));
 BUF_X4 buffer874 (.A(net870),
    .Z(net874));
 BUF_X4 buffer875 (.A(net870),
    .Z(net875));
 BUF_X4 buffer876 (.A(net870),
    .Z(net876));
 BUF_X4 buffer877 (.A(net870),
    .Z(net877));
 BUF_X4 buffer878 (.A(net870),
    .Z(net878));
 BUF_X4 buffer879 (.A(net870),
    .Z(net879));
 BUF_X4 buffer88 (.A(_10796_),
    .Z(net88));
 BUF_X4 buffer880 (.A(net870),
    .Z(net880));
 BUF_X4 buffer881 (.A(net870),
    .Z(net881));
 BUF_X4 buffer882 (.A(net870),
    .Z(net882));
 BUF_X4 buffer883 (.A(net870),
    .Z(net883));
 BUF_X4 buffer884 (.A(net870),
    .Z(net884));
 BUF_X4 buffer885 (.A(net870),
    .Z(net885));
 BUF_X4 buffer886 (.A(net870),
    .Z(net886));
 BUF_X4 buffer887 (.A(net870),
    .Z(net887));
 BUF_X4 buffer888 (.A(net870),
    .Z(net888));
 BUF_X4 buffer889 (.A(net870),
    .Z(net889));
 BUF_X4 buffer89 (.A(_10796_),
    .Z(net89));
 BUF_X4 buffer890 (.A(net870),
    .Z(net890));
 BUF_X4 buffer891 (.A(net870),
    .Z(net891));
 BUF_X4 buffer892 (.A(net870),
    .Z(net892));
 BUF_X4 buffer893 (.A(net870),
    .Z(net893));
 BUF_X4 buffer894 (.A(net870),
    .Z(net894));
 BUF_X4 buffer895 (.A(net870),
    .Z(net895));
 BUF_X4 buffer896 (.A(net870),
    .Z(net896));
 BUF_X4 buffer897 (.A(net870),
    .Z(net897));
 BUF_X4 buffer898 (.A(\icache.tag_mem.w_mask_i [230]),
    .Z(net898));
 BUF_X4 buffer899 (.A(\icache.tag_mem.w_mask_i [230]),
    .Z(net899));
 BUF_X4 buffer9 (.A(_24796_),
    .Z(net9));
 BUF_X4 buffer90 (.A(net89),
    .Z(net90));
 BUF_X4 buffer900 (.A(\icache.tag_mem.w_mask_i [203]),
    .Z(net900));
 BUF_X4 buffer901 (.A(net900),
    .Z(net901));
 BUF_X4 buffer902 (.A(net900),
    .Z(net902));
 BUF_X4 buffer903 (.A(net900),
    .Z(net903));
 BUF_X4 buffer904 (.A(net900),
    .Z(net904));
 BUF_X4 buffer905 (.A(net900),
    .Z(net905));
 BUF_X4 buffer906 (.A(net900),
    .Z(net906));
 BUF_X4 buffer907 (.A(net900),
    .Z(net907));
 BUF_X4 buffer908 (.A(net900),
    .Z(net908));
 BUF_X4 buffer909 (.A(net900),
    .Z(net909));
 BUF_X4 buffer91 (.A(_10796_),
    .Z(net91));
 BUF_X4 buffer910 (.A(net900),
    .Z(net910));
 BUF_X4 buffer911 (.A(net900),
    .Z(net911));
 BUF_X4 buffer912 (.A(net900),
    .Z(net912));
 BUF_X4 buffer913 (.A(net900),
    .Z(net913));
 BUF_X4 buffer914 (.A(net900),
    .Z(net914));
 BUF_X4 buffer915 (.A(net900),
    .Z(net915));
 BUF_X4 buffer916 (.A(net900),
    .Z(net916));
 BUF_X4 buffer917 (.A(net900),
    .Z(net917));
 BUF_X4 buffer918 (.A(net900),
    .Z(net918));
 BUF_X4 buffer919 (.A(net900),
    .Z(net919));
 BUF_X4 buffer92 (.A(net91),
    .Z(net92));
 BUF_X4 buffer920 (.A(net900),
    .Z(net920));
 BUF_X4 buffer921 (.A(net900),
    .Z(net921));
 BUF_X4 buffer922 (.A(net900),
    .Z(net922));
 BUF_X4 buffer923 (.A(net900),
    .Z(net923));
 BUF_X4 buffer924 (.A(net900),
    .Z(net924));
 BUF_X4 buffer925 (.A(net900),
    .Z(net925));
 BUF_X4 buffer926 (.A(net900),
    .Z(net926));
 BUF_X4 buffer927 (.A(net900),
    .Z(net927));
 BUF_X4 buffer928 (.A(\icache.tag_mem.w_mask_i [172]),
    .Z(net928));
 BUF_X4 buffer929 (.A(\icache.tag_mem.w_mask_i [172]),
    .Z(net929));
 BUF_X4 buffer93 (.A(net91),
    .Z(net93));
 BUF_X4 buffer930 (.A(\icache.tag_mem.w_mask_i [145]),
    .Z(net930));
 BUF_X4 buffer931 (.A(net930),
    .Z(net931));
 BUF_X4 buffer932 (.A(net930),
    .Z(net932));
 BUF_X4 buffer933 (.A(net930),
    .Z(net933));
 BUF_X4 buffer934 (.A(net930),
    .Z(net934));
 BUF_X4 buffer935 (.A(net930),
    .Z(net935));
 BUF_X4 buffer936 (.A(net930),
    .Z(net936));
 BUF_X4 buffer937 (.A(net930),
    .Z(net937));
 BUF_X4 buffer938 (.A(net930),
    .Z(net938));
 BUF_X4 buffer939 (.A(net930),
    .Z(net939));
 BUF_X4 buffer94 (.A(_11074_),
    .Z(net94));
 BUF_X4 buffer940 (.A(net930),
    .Z(net940));
 BUF_X4 buffer941 (.A(net930),
    .Z(net941));
 BUF_X4 buffer942 (.A(net930),
    .Z(net942));
 BUF_X4 buffer943 (.A(net930),
    .Z(net943));
 BUF_X4 buffer944 (.A(net930),
    .Z(net944));
 BUF_X4 buffer945 (.A(net930),
    .Z(net945));
 BUF_X4 buffer946 (.A(net930),
    .Z(net946));
 BUF_X4 buffer947 (.A(net930),
    .Z(net947));
 BUF_X4 buffer948 (.A(net930),
    .Z(net948));
 BUF_X4 buffer949 (.A(net930),
    .Z(net949));
 BUF_X4 buffer95 (.A(net94),
    .Z(net95));
 BUF_X4 buffer950 (.A(net930),
    .Z(net950));
 BUF_X4 buffer951 (.A(net930),
    .Z(net951));
 BUF_X4 buffer952 (.A(net930),
    .Z(net952));
 BUF_X4 buffer953 (.A(net930),
    .Z(net953));
 BUF_X4 buffer954 (.A(net930),
    .Z(net954));
 BUF_X4 buffer955 (.A(net930),
    .Z(net955));
 BUF_X4 buffer956 (.A(net930),
    .Z(net956));
 BUF_X4 buffer957 (.A(net930),
    .Z(net957));
 BUF_X4 buffer958 (.A(_07997_),
    .Z(net958));
 BUF_X4 buffer959 (.A(\icache.tag_mem.w_mask_i [201]),
    .Z(net959));
 BUF_X4 buffer96 (.A(net95),
    .Z(net96));
 BUF_X4 buffer960 (.A(\icache.tag_mem.w_mask_i [201]),
    .Z(net960));
 BUF_X4 buffer961 (.A(\icache.tag_mem.w_mask_i [174]),
    .Z(net961));
 BUF_X4 buffer962 (.A(net961),
    .Z(net962));
 BUF_X4 buffer963 (.A(net961),
    .Z(net963));
 BUF_X4 buffer964 (.A(net961),
    .Z(net964));
 BUF_X4 buffer965 (.A(net961),
    .Z(net965));
 BUF_X4 buffer966 (.A(net961),
    .Z(net966));
 BUF_X4 buffer967 (.A(net961),
    .Z(net967));
 BUF_X4 buffer968 (.A(net961),
    .Z(net968));
 BUF_X4 buffer969 (.A(net961),
    .Z(net969));
 BUF_X4 buffer97 (.A(_11030_),
    .Z(net97));
 BUF_X4 buffer970 (.A(net961),
    .Z(net970));
 BUF_X4 buffer971 (.A(net961),
    .Z(net971));
 BUF_X4 buffer972 (.A(net961),
    .Z(net972));
 BUF_X4 buffer973 (.A(net961),
    .Z(net973));
 BUF_X4 buffer974 (.A(net961),
    .Z(net974));
 BUF_X4 buffer975 (.A(net961),
    .Z(net975));
 BUF_X4 buffer976 (.A(net961),
    .Z(net976));
 BUF_X4 buffer977 (.A(net961),
    .Z(net977));
 BUF_X4 buffer978 (.A(net961),
    .Z(net978));
 BUF_X4 buffer979 (.A(net961),
    .Z(net979));
 BUF_X4 buffer98 (.A(net97),
    .Z(net98));
 BUF_X4 buffer980 (.A(net961),
    .Z(net980));
 BUF_X4 buffer981 (.A(net961),
    .Z(net981));
 BUF_X4 buffer982 (.A(net961),
    .Z(net982));
 BUF_X4 buffer983 (.A(net961),
    .Z(net983));
 BUF_X4 buffer984 (.A(net961),
    .Z(net984));
 BUF_X4 buffer985 (.A(net961),
    .Z(net985));
 BUF_X4 buffer986 (.A(net961),
    .Z(net986));
 BUF_X4 buffer987 (.A(net961),
    .Z(net987));
 BUF_X4 buffer988 (.A(net961),
    .Z(net988));
 BUF_X4 buffer989 (.A(\icache.tag_mem.w_mask_i [27]),
    .Z(net989));
 BUF_X4 buffer99 (.A(net97),
    .Z(net99));
 BUF_X4 buffer990 (.A(net989),
    .Z(net990));
 BUF_X4 buffer991 (.A(net990),
    .Z(net991));
 BUF_X4 buffer992 (.A(net990),
    .Z(net992));
 BUF_X4 buffer993 (.A(\icache.stat_mem.w_i ),
    .Z(net993));
 BUF_X4 buffer994 (.A(\icache.stat_mem.data_i [3]),
    .Z(net994));
 BUF_X4 buffer995 (.A(\icache.stat_mem.data_i [1]),
    .Z(net995));
 BUF_X4 buffer996 (.A(\icache.stat_mem.w_mask_i [3]),
    .Z(net996));
 BUF_X4 buffer997 (.A(\icache.stat_mem.w_mask_i [1]),
    .Z(net997));
 BUF_X4 buffer998 (.A(\icache.stat_mem.w_mask_i [6]),
    .Z(net998));
 BUF_X4 buffer999 (.A(\icache.stat_mem.w_mask_i [2]),
    .Z(net999));
 nangate45_64x512_1P_BM \icache.data_mems_0__data_mem.macro_mem  (.we_in(net214),
    .clk(clk_i),
    .ce_in(net226),
    .addr_in({net125,
    net134,
    net143,
    net152,
    net189,
    net198,
    net161,
    net166,
    net115}),
    .rd_out({\icache.data_mems_0__data_mem.data_o [63],
    \icache.data_mems_0__data_mem.data_o [62],
    \icache.data_mems_0__data_mem.data_o [61],
    \icache.data_mems_0__data_mem.data_o [60],
    \icache.data_mems_0__data_mem.data_o [59],
    \icache.data_mems_0__data_mem.data_o [58],
    \icache.data_mems_0__data_mem.data_o [57],
    \icache.data_mems_0__data_mem.data_o [56],
    \icache.data_mems_0__data_mem.data_o [55],
    \icache.data_mems_0__data_mem.data_o [54],
    \icache.data_mems_0__data_mem.data_o [53],
    \icache.data_mems_0__data_mem.data_o [52],
    \icache.data_mems_0__data_mem.data_o [51],
    \icache.data_mems_0__data_mem.data_o [50],
    \icache.data_mems_0__data_mem.data_o [49],
    \icache.data_mems_0__data_mem.data_o [48],
    \icache.data_mems_0__data_mem.data_o [47],
    \icache.data_mems_0__data_mem.data_o [46],
    \icache.data_mems_0__data_mem.data_o [45],
    \icache.data_mems_0__data_mem.data_o [44],
    \icache.data_mems_0__data_mem.data_o [43],
    \icache.data_mems_0__data_mem.data_o [42],
    \icache.data_mems_0__data_mem.data_o [41],
    \icache.data_mems_0__data_mem.data_o [40],
    \icache.data_mems_0__data_mem.data_o [39],
    \icache.data_mems_0__data_mem.data_o [38],
    \icache.data_mems_0__data_mem.data_o [37],
    \icache.data_mems_0__data_mem.data_o [36],
    \icache.data_mems_0__data_mem.data_o [35],
    \icache.data_mems_0__data_mem.data_o [34],
    \icache.data_mems_0__data_mem.data_o [33],
    \icache.data_mems_0__data_mem.data_o [32],
    \icache.data_mems_0__data_mem.data_o [31],
    \icache.data_mems_0__data_mem.data_o [30],
    \icache.data_mems_0__data_mem.data_o [29],
    \icache.data_mems_0__data_mem.data_o [28],
    \icache.data_mems_0__data_mem.data_o [27],
    \icache.data_mems_0__data_mem.data_o [26],
    \icache.data_mems_0__data_mem.data_o [25],
    \icache.data_mems_0__data_mem.data_o [24],
    \icache.data_mems_0__data_mem.data_o [23],
    \icache.data_mems_0__data_mem.data_o [22],
    \icache.data_mems_0__data_mem.data_o [21],
    \icache.data_mems_0__data_mem.data_o [20],
    \icache.data_mems_0__data_mem.data_o [19],
    \icache.data_mems_0__data_mem.data_o [18],
    \icache.data_mems_0__data_mem.data_o [17],
    \icache.data_mems_0__data_mem.data_o [16],
    \icache.data_mems_0__data_mem.data_o [15],
    \icache.data_mems_0__data_mem.data_o [14],
    \icache.data_mems_0__data_mem.data_o [13],
    \icache.data_mems_0__data_mem.data_o [12],
    \icache.data_mems_0__data_mem.data_o [11],
    \icache.data_mems_0__data_mem.data_o [10],
    \icache.data_mems_0__data_mem.data_o [9],
    \icache.data_mems_0__data_mem.data_o [8],
    \icache.data_mems_0__data_mem.data_o [7],
    \icache.data_mems_0__data_mem.data_o [6],
    \icache.data_mems_0__data_mem.data_o [5],
    \icache.data_mems_0__data_mem.data_o [4],
    \icache.data_mems_0__data_mem.data_o [3],
    \icache.data_mems_0__data_mem.data_o [2],
    \icache.data_mems_0__data_mem.data_o [1],
    \icache.data_mems_0__data_mem.data_o [0]}),
    .w_mask_in({_NC1,
    _NC2,
    _NC3,
    _NC4,
    _NC5,
    _NC6,
    _NC7,
    _NC8,
    _NC9,
    _NC10,
    _NC11,
    _NC12,
    _NC13,
    _NC14,
    _NC15,
    _NC16,
    _NC17,
    _NC18,
    _NC19,
    _NC20,
    _NC21,
    _NC22,
    _NC23,
    _NC24,
    _NC25,
    _NC26,
    _NC27,
    _NC28,
    _NC29,
    _NC30,
    _NC31,
    _NC32,
    _NC33,
    _NC34,
    _NC35,
    _NC36,
    _NC37,
    _NC38,
    _NC39,
    _NC40,
    _NC41,
    _NC42,
    _NC43,
    _NC44,
    _NC45,
    _NC46,
    _NC47,
    _NC48,
    _NC49,
    _NC50,
    _NC51,
    _NC52,
    _NC53,
    _NC54,
    _NC55,
    _NC56,
    _NC57,
    _NC58,
    _NC59,
    _NC60,
    _NC61,
    _NC62,
    _NC63,
    _NC64}),
    .wd_in({net686,
    net687,
    net688,
    net689,
    net690,
    net691,
    net692,
    net693,
    net694,
    net695,
    net696,
    net697,
    net698,
    net699,
    net700,
    net701,
    net702,
    net703,
    net704,
    net705,
    net706,
    net707,
    net708,
    net709,
    net710,
    net711,
    net712,
    net713,
    net714,
    net715,
    net716,
    net717,
    net718,
    net719,
    net720,
    net721,
    net722,
    net723,
    net724,
    net725,
    net726,
    net727,
    net728,
    net729,
    net730,
    net731,
    net732,
    net733,
    net734,
    net735,
    net736,
    net737,
    net738,
    net739,
    net740,
    net741,
    net742,
    net743,
    net744,
    net745,
    net746,
    net747,
    net748,
    net749}));
 nangate45_64x512_1P_BM \icache.data_mems_1__data_mem.macro_mem  (.we_in(net215),
    .clk(clk_i),
    .ce_in(net227),
    .addr_in({net126,
    net135,
    net144,
    net153,
    net190,
    net199,
    net162,
    net167,
    net120}),
    .rd_out({\icache.data_mems_1__data_mem.data_o [63],
    \icache.data_mems_1__data_mem.data_o [62],
    \icache.data_mems_1__data_mem.data_o [61],
    \icache.data_mems_1__data_mem.data_o [60],
    \icache.data_mems_1__data_mem.data_o [59],
    \icache.data_mems_1__data_mem.data_o [58],
    \icache.data_mems_1__data_mem.data_o [57],
    \icache.data_mems_1__data_mem.data_o [56],
    \icache.data_mems_1__data_mem.data_o [55],
    \icache.data_mems_1__data_mem.data_o [54],
    \icache.data_mems_1__data_mem.data_o [53],
    \icache.data_mems_1__data_mem.data_o [52],
    \icache.data_mems_1__data_mem.data_o [51],
    \icache.data_mems_1__data_mem.data_o [50],
    \icache.data_mems_1__data_mem.data_o [49],
    \icache.data_mems_1__data_mem.data_o [48],
    \icache.data_mems_1__data_mem.data_o [47],
    \icache.data_mems_1__data_mem.data_o [46],
    \icache.data_mems_1__data_mem.data_o [45],
    \icache.data_mems_1__data_mem.data_o [44],
    \icache.data_mems_1__data_mem.data_o [43],
    \icache.data_mems_1__data_mem.data_o [42],
    \icache.data_mems_1__data_mem.data_o [41],
    \icache.data_mems_1__data_mem.data_o [40],
    \icache.data_mems_1__data_mem.data_o [39],
    \icache.data_mems_1__data_mem.data_o [38],
    \icache.data_mems_1__data_mem.data_o [37],
    \icache.data_mems_1__data_mem.data_o [36],
    \icache.data_mems_1__data_mem.data_o [35],
    \icache.data_mems_1__data_mem.data_o [34],
    \icache.data_mems_1__data_mem.data_o [33],
    \icache.data_mems_1__data_mem.data_o [32],
    \icache.data_mems_1__data_mem.data_o [31],
    \icache.data_mems_1__data_mem.data_o [30],
    \icache.data_mems_1__data_mem.data_o [29],
    \icache.data_mems_1__data_mem.data_o [28],
    \icache.data_mems_1__data_mem.data_o [27],
    \icache.data_mems_1__data_mem.data_o [26],
    \icache.data_mems_1__data_mem.data_o [25],
    \icache.data_mems_1__data_mem.data_o [24],
    \icache.data_mems_1__data_mem.data_o [23],
    \icache.data_mems_1__data_mem.data_o [22],
    \icache.data_mems_1__data_mem.data_o [21],
    \icache.data_mems_1__data_mem.data_o [20],
    \icache.data_mems_1__data_mem.data_o [19],
    \icache.data_mems_1__data_mem.data_o [18],
    \icache.data_mems_1__data_mem.data_o [17],
    \icache.data_mems_1__data_mem.data_o [16],
    \icache.data_mems_1__data_mem.data_o [15],
    \icache.data_mems_1__data_mem.data_o [14],
    \icache.data_mems_1__data_mem.data_o [13],
    \icache.data_mems_1__data_mem.data_o [12],
    \icache.data_mems_1__data_mem.data_o [11],
    \icache.data_mems_1__data_mem.data_o [10],
    \icache.data_mems_1__data_mem.data_o [9],
    \icache.data_mems_1__data_mem.data_o [8],
    \icache.data_mems_1__data_mem.data_o [7],
    \icache.data_mems_1__data_mem.data_o [6],
    \icache.data_mems_1__data_mem.data_o [5],
    \icache.data_mems_1__data_mem.data_o [4],
    \icache.data_mems_1__data_mem.data_o [3],
    \icache.data_mems_1__data_mem.data_o [2],
    \icache.data_mems_1__data_mem.data_o [1],
    \icache.data_mems_1__data_mem.data_o [0]}),
    .w_mask_in({_NC65,
    _NC66,
    _NC67,
    _NC68,
    _NC69,
    _NC70,
    _NC71,
    _NC72,
    _NC73,
    _NC74,
    _NC75,
    _NC76,
    _NC77,
    _NC78,
    _NC79,
    _NC80,
    _NC81,
    _NC82,
    _NC83,
    _NC84,
    _NC85,
    _NC86,
    _NC87,
    _NC88,
    _NC89,
    _NC90,
    _NC91,
    _NC92,
    _NC93,
    _NC94,
    _NC95,
    _NC96,
    _NC97,
    _NC98,
    _NC99,
    _NC100,
    _NC101,
    _NC102,
    _NC103,
    _NC104,
    _NC105,
    _NC106,
    _NC107,
    _NC108,
    _NC109,
    _NC110,
    _NC111,
    _NC112,
    _NC113,
    _NC114,
    _NC115,
    _NC116,
    _NC117,
    _NC118,
    _NC119,
    _NC120,
    _NC121,
    _NC122,
    _NC123,
    _NC124,
    _NC125,
    _NC126,
    _NC127,
    _NC128}),
    .wd_in({net622,
    net623,
    net624,
    net625,
    net626,
    net627,
    net628,
    net629,
    net630,
    net631,
    net632,
    net633,
    net634,
    net635,
    net636,
    net637,
    net638,
    net639,
    net640,
    net641,
    net642,
    net643,
    net644,
    net645,
    net646,
    net647,
    net648,
    net649,
    net650,
    net651,
    net652,
    net653,
    net654,
    net655,
    net656,
    net657,
    net658,
    net659,
    net660,
    net661,
    net662,
    net663,
    net664,
    net665,
    net666,
    net667,
    net668,
    net669,
    net670,
    net671,
    net672,
    net673,
    net674,
    net675,
    net676,
    net677,
    net678,
    net679,
    net680,
    net681,
    net682,
    net683,
    net684,
    net685}));
 nangate45_64x512_1P_BM \icache.data_mems_2__data_mem.macro_mem  (.we_in(net216),
    .clk(clk_i),
    .ce_in(net228),
    .addr_in({net127,
    net136,
    net145,
    net154,
    net191,
    net200,
    net164,
    net171,
    net116}),
    .rd_out({\icache.data_mems_2__data_mem.data_o [63],
    \icache.data_mems_2__data_mem.data_o [62],
    \icache.data_mems_2__data_mem.data_o [61],
    \icache.data_mems_2__data_mem.data_o [60],
    \icache.data_mems_2__data_mem.data_o [59],
    \icache.data_mems_2__data_mem.data_o [58],
    \icache.data_mems_2__data_mem.data_o [57],
    \icache.data_mems_2__data_mem.data_o [56],
    \icache.data_mems_2__data_mem.data_o [55],
    \icache.data_mems_2__data_mem.data_o [54],
    \icache.data_mems_2__data_mem.data_o [53],
    \icache.data_mems_2__data_mem.data_o [52],
    \icache.data_mems_2__data_mem.data_o [51],
    \icache.data_mems_2__data_mem.data_o [50],
    \icache.data_mems_2__data_mem.data_o [49],
    \icache.data_mems_2__data_mem.data_o [48],
    \icache.data_mems_2__data_mem.data_o [47],
    \icache.data_mems_2__data_mem.data_o [46],
    \icache.data_mems_2__data_mem.data_o [45],
    \icache.data_mems_2__data_mem.data_o [44],
    \icache.data_mems_2__data_mem.data_o [43],
    \icache.data_mems_2__data_mem.data_o [42],
    \icache.data_mems_2__data_mem.data_o [41],
    \icache.data_mems_2__data_mem.data_o [40],
    \icache.data_mems_2__data_mem.data_o [39],
    \icache.data_mems_2__data_mem.data_o [38],
    \icache.data_mems_2__data_mem.data_o [37],
    \icache.data_mems_2__data_mem.data_o [36],
    \icache.data_mems_2__data_mem.data_o [35],
    \icache.data_mems_2__data_mem.data_o [34],
    \icache.data_mems_2__data_mem.data_o [33],
    \icache.data_mems_2__data_mem.data_o [32],
    \icache.data_mems_2__data_mem.data_o [31],
    \icache.data_mems_2__data_mem.data_o [30],
    \icache.data_mems_2__data_mem.data_o [29],
    \icache.data_mems_2__data_mem.data_o [28],
    \icache.data_mems_2__data_mem.data_o [27],
    \icache.data_mems_2__data_mem.data_o [26],
    \icache.data_mems_2__data_mem.data_o [25],
    \icache.data_mems_2__data_mem.data_o [24],
    \icache.data_mems_2__data_mem.data_o [23],
    \icache.data_mems_2__data_mem.data_o [22],
    \icache.data_mems_2__data_mem.data_o [21],
    \icache.data_mems_2__data_mem.data_o [20],
    \icache.data_mems_2__data_mem.data_o [19],
    \icache.data_mems_2__data_mem.data_o [18],
    \icache.data_mems_2__data_mem.data_o [17],
    \icache.data_mems_2__data_mem.data_o [16],
    \icache.data_mems_2__data_mem.data_o [15],
    \icache.data_mems_2__data_mem.data_o [14],
    \icache.data_mems_2__data_mem.data_o [13],
    \icache.data_mems_2__data_mem.data_o [12],
    \icache.data_mems_2__data_mem.data_o [11],
    \icache.data_mems_2__data_mem.data_o [10],
    \icache.data_mems_2__data_mem.data_o [9],
    \icache.data_mems_2__data_mem.data_o [8],
    \icache.data_mems_2__data_mem.data_o [7],
    \icache.data_mems_2__data_mem.data_o [6],
    \icache.data_mems_2__data_mem.data_o [5],
    \icache.data_mems_2__data_mem.data_o [4],
    \icache.data_mems_2__data_mem.data_o [3],
    \icache.data_mems_2__data_mem.data_o [2],
    \icache.data_mems_2__data_mem.data_o [1],
    \icache.data_mems_2__data_mem.data_o [0]}),
    .w_mask_in({_NC129,
    _NC130,
    _NC131,
    _NC132,
    _NC133,
    _NC134,
    _NC135,
    _NC136,
    _NC137,
    _NC138,
    _NC139,
    _NC140,
    _NC141,
    _NC142,
    _NC143,
    _NC144,
    _NC145,
    _NC146,
    _NC147,
    _NC148,
    _NC149,
    _NC150,
    _NC151,
    _NC152,
    _NC153,
    _NC154,
    _NC155,
    _NC156,
    _NC157,
    _NC158,
    _NC159,
    _NC160,
    _NC161,
    _NC162,
    _NC163,
    _NC164,
    _NC165,
    _NC166,
    _NC167,
    _NC168,
    _NC169,
    _NC170,
    _NC171,
    _NC172,
    _NC173,
    _NC174,
    _NC175,
    _NC176,
    _NC177,
    _NC178,
    _NC179,
    _NC180,
    _NC181,
    _NC182,
    _NC183,
    _NC184,
    _NC185,
    _NC186,
    _NC187,
    _NC188,
    _NC189,
    _NC190,
    _NC191,
    _NC192}),
    .wd_in({net558,
    net559,
    net560,
    net561,
    net562,
    net563,
    net564,
    net565,
    net566,
    net567,
    net568,
    net569,
    net570,
    net571,
    net572,
    net573,
    net574,
    net575,
    net576,
    net577,
    net578,
    net579,
    net580,
    net581,
    net582,
    net583,
    net584,
    net585,
    net586,
    net587,
    net588,
    net589,
    net590,
    net591,
    net592,
    net593,
    net594,
    net595,
    net596,
    net597,
    net598,
    net599,
    net600,
    net601,
    net602,
    net603,
    net604,
    net605,
    net606,
    net607,
    net608,
    net609,
    net610,
    net611,
    net612,
    net613,
    net614,
    net615,
    net616,
    net617,
    net618,
    net619,
    net620,
    net621}));
 nangate45_64x512_1P_BM \icache.data_mems_3__data_mem.macro_mem  (.we_in(net217),
    .clk(clk_i),
    .ce_in(net229),
    .addr_in({net128,
    net137,
    net146,
    net155,
    net192,
    net201,
    net163,
    net172,
    net121}),
    .rd_out({\icache.data_mems_3__data_mem.data_o [63],
    \icache.data_mems_3__data_mem.data_o [62],
    \icache.data_mems_3__data_mem.data_o [61],
    \icache.data_mems_3__data_mem.data_o [60],
    \icache.data_mems_3__data_mem.data_o [59],
    \icache.data_mems_3__data_mem.data_o [58],
    \icache.data_mems_3__data_mem.data_o [57],
    \icache.data_mems_3__data_mem.data_o [56],
    \icache.data_mems_3__data_mem.data_o [55],
    \icache.data_mems_3__data_mem.data_o [54],
    \icache.data_mems_3__data_mem.data_o [53],
    \icache.data_mems_3__data_mem.data_o [52],
    \icache.data_mems_3__data_mem.data_o [51],
    \icache.data_mems_3__data_mem.data_o [50],
    \icache.data_mems_3__data_mem.data_o [49],
    \icache.data_mems_3__data_mem.data_o [48],
    \icache.data_mems_3__data_mem.data_o [47],
    \icache.data_mems_3__data_mem.data_o [46],
    \icache.data_mems_3__data_mem.data_o [45],
    \icache.data_mems_3__data_mem.data_o [44],
    \icache.data_mems_3__data_mem.data_o [43],
    \icache.data_mems_3__data_mem.data_o [42],
    \icache.data_mems_3__data_mem.data_o [41],
    \icache.data_mems_3__data_mem.data_o [40],
    \icache.data_mems_3__data_mem.data_o [39],
    \icache.data_mems_3__data_mem.data_o [38],
    \icache.data_mems_3__data_mem.data_o [37],
    \icache.data_mems_3__data_mem.data_o [36],
    \icache.data_mems_3__data_mem.data_o [35],
    \icache.data_mems_3__data_mem.data_o [34],
    \icache.data_mems_3__data_mem.data_o [33],
    \icache.data_mems_3__data_mem.data_o [32],
    \icache.data_mems_3__data_mem.data_o [31],
    \icache.data_mems_3__data_mem.data_o [30],
    \icache.data_mems_3__data_mem.data_o [29],
    \icache.data_mems_3__data_mem.data_o [28],
    \icache.data_mems_3__data_mem.data_o [27],
    \icache.data_mems_3__data_mem.data_o [26],
    \icache.data_mems_3__data_mem.data_o [25],
    \icache.data_mems_3__data_mem.data_o [24],
    \icache.data_mems_3__data_mem.data_o [23],
    \icache.data_mems_3__data_mem.data_o [22],
    \icache.data_mems_3__data_mem.data_o [21],
    \icache.data_mems_3__data_mem.data_o [20],
    \icache.data_mems_3__data_mem.data_o [19],
    \icache.data_mems_3__data_mem.data_o [18],
    \icache.data_mems_3__data_mem.data_o [17],
    \icache.data_mems_3__data_mem.data_o [16],
    \icache.data_mems_3__data_mem.data_o [15],
    \icache.data_mems_3__data_mem.data_o [14],
    \icache.data_mems_3__data_mem.data_o [13],
    \icache.data_mems_3__data_mem.data_o [12],
    \icache.data_mems_3__data_mem.data_o [11],
    \icache.data_mems_3__data_mem.data_o [10],
    \icache.data_mems_3__data_mem.data_o [9],
    \icache.data_mems_3__data_mem.data_o [8],
    \icache.data_mems_3__data_mem.data_o [7],
    \icache.data_mems_3__data_mem.data_o [6],
    \icache.data_mems_3__data_mem.data_o [5],
    \icache.data_mems_3__data_mem.data_o [4],
    \icache.data_mems_3__data_mem.data_o [3],
    \icache.data_mems_3__data_mem.data_o [2],
    \icache.data_mems_3__data_mem.data_o [1],
    \icache.data_mems_3__data_mem.data_o [0]}),
    .w_mask_in({_NC193,
    _NC194,
    _NC195,
    _NC196,
    _NC197,
    _NC198,
    _NC199,
    _NC200,
    _NC201,
    _NC202,
    _NC203,
    _NC204,
    _NC205,
    _NC206,
    _NC207,
    _NC208,
    _NC209,
    _NC210,
    _NC211,
    _NC212,
    _NC213,
    _NC214,
    _NC215,
    _NC216,
    _NC217,
    _NC218,
    _NC219,
    _NC220,
    _NC221,
    _NC222,
    _NC223,
    _NC224,
    _NC225,
    _NC226,
    _NC227,
    _NC228,
    _NC229,
    _NC230,
    _NC231,
    _NC232,
    _NC233,
    _NC234,
    _NC235,
    _NC236,
    _NC237,
    _NC238,
    _NC239,
    _NC240,
    _NC241,
    _NC242,
    _NC243,
    _NC244,
    _NC245,
    _NC246,
    _NC247,
    _NC248,
    _NC249,
    _NC250,
    _NC251,
    _NC252,
    _NC253,
    _NC254,
    _NC255,
    _NC256}),
    .wd_in({net494,
    net495,
    net496,
    net497,
    net498,
    net499,
    net500,
    net501,
    net502,
    net503,
    net504,
    net505,
    net506,
    net507,
    net508,
    net509,
    net510,
    net511,
    net512,
    net513,
    net514,
    net515,
    net516,
    net517,
    net518,
    net519,
    net520,
    net521,
    net522,
    net523,
    net524,
    net525,
    net526,
    net527,
    net528,
    net529,
    net530,
    net531,
    net532,
    net533,
    net534,
    net535,
    net536,
    net537,
    net538,
    net539,
    net540,
    net541,
    net542,
    net543,
    net544,
    net545,
    net546,
    net547,
    net548,
    net549,
    net550,
    net551,
    net552,
    net553,
    net554,
    net555,
    net556,
    net557}));
 nangate45_64x512_1P_BM \icache.data_mems_4__data_mem.macro_mem  (.we_in(net218),
    .clk(clk_i),
    .ce_in(net230),
    .addr_in({net129,
    net138,
    net147,
    net156,
    net193,
    net202,
    net176,
    net169,
    net118}),
    .rd_out({\icache.data_mems_4__data_mem.data_o [63],
    \icache.data_mems_4__data_mem.data_o [62],
    \icache.data_mems_4__data_mem.data_o [61],
    \icache.data_mems_4__data_mem.data_o [60],
    \icache.data_mems_4__data_mem.data_o [59],
    \icache.data_mems_4__data_mem.data_o [58],
    \icache.data_mems_4__data_mem.data_o [57],
    \icache.data_mems_4__data_mem.data_o [56],
    \icache.data_mems_4__data_mem.data_o [55],
    \icache.data_mems_4__data_mem.data_o [54],
    \icache.data_mems_4__data_mem.data_o [53],
    \icache.data_mems_4__data_mem.data_o [52],
    \icache.data_mems_4__data_mem.data_o [51],
    \icache.data_mems_4__data_mem.data_o [50],
    \icache.data_mems_4__data_mem.data_o [49],
    \icache.data_mems_4__data_mem.data_o [48],
    \icache.data_mems_4__data_mem.data_o [47],
    \icache.data_mems_4__data_mem.data_o [46],
    \icache.data_mems_4__data_mem.data_o [45],
    \icache.data_mems_4__data_mem.data_o [44],
    \icache.data_mems_4__data_mem.data_o [43],
    \icache.data_mems_4__data_mem.data_o [42],
    \icache.data_mems_4__data_mem.data_o [41],
    \icache.data_mems_4__data_mem.data_o [40],
    \icache.data_mems_4__data_mem.data_o [39],
    \icache.data_mems_4__data_mem.data_o [38],
    \icache.data_mems_4__data_mem.data_o [37],
    \icache.data_mems_4__data_mem.data_o [36],
    \icache.data_mems_4__data_mem.data_o [35],
    \icache.data_mems_4__data_mem.data_o [34],
    \icache.data_mems_4__data_mem.data_o [33],
    \icache.data_mems_4__data_mem.data_o [32],
    \icache.data_mems_4__data_mem.data_o [31],
    \icache.data_mems_4__data_mem.data_o [30],
    \icache.data_mems_4__data_mem.data_o [29],
    \icache.data_mems_4__data_mem.data_o [28],
    \icache.data_mems_4__data_mem.data_o [27],
    \icache.data_mems_4__data_mem.data_o [26],
    \icache.data_mems_4__data_mem.data_o [25],
    \icache.data_mems_4__data_mem.data_o [24],
    \icache.data_mems_4__data_mem.data_o [23],
    \icache.data_mems_4__data_mem.data_o [22],
    \icache.data_mems_4__data_mem.data_o [21],
    \icache.data_mems_4__data_mem.data_o [20],
    \icache.data_mems_4__data_mem.data_o [19],
    \icache.data_mems_4__data_mem.data_o [18],
    \icache.data_mems_4__data_mem.data_o [17],
    \icache.data_mems_4__data_mem.data_o [16],
    \icache.data_mems_4__data_mem.data_o [15],
    \icache.data_mems_4__data_mem.data_o [14],
    \icache.data_mems_4__data_mem.data_o [13],
    \icache.data_mems_4__data_mem.data_o [12],
    \icache.data_mems_4__data_mem.data_o [11],
    \icache.data_mems_4__data_mem.data_o [10],
    \icache.data_mems_4__data_mem.data_o [9],
    \icache.data_mems_4__data_mem.data_o [8],
    \icache.data_mems_4__data_mem.data_o [7],
    \icache.data_mems_4__data_mem.data_o [6],
    \icache.data_mems_4__data_mem.data_o [5],
    \icache.data_mems_4__data_mem.data_o [4],
    \icache.data_mems_4__data_mem.data_o [3],
    \icache.data_mems_4__data_mem.data_o [2],
    \icache.data_mems_4__data_mem.data_o [1],
    \icache.data_mems_4__data_mem.data_o [0]}),
    .w_mask_in({_NC257,
    _NC258,
    _NC259,
    _NC260,
    _NC261,
    _NC262,
    _NC263,
    _NC264,
    _NC265,
    _NC266,
    _NC267,
    _NC268,
    _NC269,
    _NC270,
    _NC271,
    _NC272,
    _NC273,
    _NC274,
    _NC275,
    _NC276,
    _NC277,
    _NC278,
    _NC279,
    _NC280,
    _NC281,
    _NC282,
    _NC283,
    _NC284,
    _NC285,
    _NC286,
    _NC287,
    _NC288,
    _NC289,
    _NC290,
    _NC291,
    _NC292,
    _NC293,
    _NC294,
    _NC295,
    _NC296,
    _NC297,
    _NC298,
    _NC299,
    _NC300,
    _NC301,
    _NC302,
    _NC303,
    _NC304,
    _NC305,
    _NC306,
    _NC307,
    _NC308,
    _NC309,
    _NC310,
    _NC311,
    _NC312,
    _NC313,
    _NC314,
    _NC315,
    _NC316,
    _NC317,
    _NC318,
    _NC319,
    _NC320}),
    .wd_in({net430,
    net431,
    net432,
    net433,
    net434,
    net435,
    net436,
    net437,
    net438,
    net439,
    net440,
    net441,
    net442,
    net443,
    net444,
    net445,
    net446,
    net447,
    net448,
    net449,
    net450,
    net451,
    net452,
    net453,
    net454,
    net455,
    net456,
    net457,
    net458,
    net459,
    net460,
    net461,
    net462,
    net463,
    net464,
    net465,
    net466,
    net467,
    net468,
    net469,
    net470,
    net471,
    net472,
    net473,
    net474,
    net475,
    net476,
    net477,
    net478,
    net479,
    net480,
    net481,
    net482,
    net483,
    net484,
    net485,
    net486,
    net487,
    net488,
    net489,
    net490,
    net491,
    net492,
    net493}));
 nangate45_64x512_1P_BM \icache.data_mems_5__data_mem.macro_mem  (.we_in(net219),
    .clk(clk_i),
    .ce_in(net231),
    .addr_in({net130,
    net139,
    net148,
    net157,
    net194,
    net203,
    net177,
    net168,
    net123}),
    .rd_out({\icache.data_mems_5__data_mem.data_o [63],
    \icache.data_mems_5__data_mem.data_o [62],
    \icache.data_mems_5__data_mem.data_o [61],
    \icache.data_mems_5__data_mem.data_o [60],
    \icache.data_mems_5__data_mem.data_o [59],
    \icache.data_mems_5__data_mem.data_o [58],
    \icache.data_mems_5__data_mem.data_o [57],
    \icache.data_mems_5__data_mem.data_o [56],
    \icache.data_mems_5__data_mem.data_o [55],
    \icache.data_mems_5__data_mem.data_o [54],
    \icache.data_mems_5__data_mem.data_o [53],
    \icache.data_mems_5__data_mem.data_o [52],
    \icache.data_mems_5__data_mem.data_o [51],
    \icache.data_mems_5__data_mem.data_o [50],
    \icache.data_mems_5__data_mem.data_o [49],
    \icache.data_mems_5__data_mem.data_o [48],
    \icache.data_mems_5__data_mem.data_o [47],
    \icache.data_mems_5__data_mem.data_o [46],
    \icache.data_mems_5__data_mem.data_o [45],
    \icache.data_mems_5__data_mem.data_o [44],
    \icache.data_mems_5__data_mem.data_o [43],
    \icache.data_mems_5__data_mem.data_o [42],
    \icache.data_mems_5__data_mem.data_o [41],
    \icache.data_mems_5__data_mem.data_o [40],
    \icache.data_mems_5__data_mem.data_o [39],
    \icache.data_mems_5__data_mem.data_o [38],
    \icache.data_mems_5__data_mem.data_o [37],
    \icache.data_mems_5__data_mem.data_o [36],
    \icache.data_mems_5__data_mem.data_o [35],
    \icache.data_mems_5__data_mem.data_o [34],
    \icache.data_mems_5__data_mem.data_o [33],
    \icache.data_mems_5__data_mem.data_o [32],
    \icache.data_mems_5__data_mem.data_o [31],
    \icache.data_mems_5__data_mem.data_o [30],
    \icache.data_mems_5__data_mem.data_o [29],
    \icache.data_mems_5__data_mem.data_o [28],
    \icache.data_mems_5__data_mem.data_o [27],
    \icache.data_mems_5__data_mem.data_o [26],
    \icache.data_mems_5__data_mem.data_o [25],
    \icache.data_mems_5__data_mem.data_o [24],
    \icache.data_mems_5__data_mem.data_o [23],
    \icache.data_mems_5__data_mem.data_o [22],
    \icache.data_mems_5__data_mem.data_o [21],
    \icache.data_mems_5__data_mem.data_o [20],
    \icache.data_mems_5__data_mem.data_o [19],
    \icache.data_mems_5__data_mem.data_o [18],
    \icache.data_mems_5__data_mem.data_o [17],
    \icache.data_mems_5__data_mem.data_o [16],
    \icache.data_mems_5__data_mem.data_o [15],
    \icache.data_mems_5__data_mem.data_o [14],
    \icache.data_mems_5__data_mem.data_o [13],
    \icache.data_mems_5__data_mem.data_o [12],
    \icache.data_mems_5__data_mem.data_o [11],
    \icache.data_mems_5__data_mem.data_o [10],
    \icache.data_mems_5__data_mem.data_o [9],
    \icache.data_mems_5__data_mem.data_o [8],
    \icache.data_mems_5__data_mem.data_o [7],
    \icache.data_mems_5__data_mem.data_o [6],
    \icache.data_mems_5__data_mem.data_o [5],
    \icache.data_mems_5__data_mem.data_o [4],
    \icache.data_mems_5__data_mem.data_o [3],
    \icache.data_mems_5__data_mem.data_o [2],
    \icache.data_mems_5__data_mem.data_o [1],
    \icache.data_mems_5__data_mem.data_o [0]}),
    .w_mask_in({_NC321,
    _NC322,
    _NC323,
    _NC324,
    _NC325,
    _NC326,
    _NC327,
    _NC328,
    _NC329,
    _NC330,
    _NC331,
    _NC332,
    _NC333,
    _NC334,
    _NC335,
    _NC336,
    _NC337,
    _NC338,
    _NC339,
    _NC340,
    _NC341,
    _NC342,
    _NC343,
    _NC344,
    _NC345,
    _NC346,
    _NC347,
    _NC348,
    _NC349,
    _NC350,
    _NC351,
    _NC352,
    _NC353,
    _NC354,
    _NC355,
    _NC356,
    _NC357,
    _NC358,
    _NC359,
    _NC360,
    _NC361,
    _NC362,
    _NC363,
    _NC364,
    _NC365,
    _NC366,
    _NC367,
    _NC368,
    _NC369,
    _NC370,
    _NC371,
    _NC372,
    _NC373,
    _NC374,
    _NC375,
    _NC376,
    _NC377,
    _NC378,
    _NC379,
    _NC380,
    _NC381,
    _NC382,
    _NC383,
    _NC384}),
    .wd_in({net366,
    net367,
    net368,
    net369,
    net370,
    net371,
    net372,
    net373,
    net374,
    net375,
    net376,
    net377,
    net378,
    net379,
    net380,
    net381,
    net382,
    net383,
    net384,
    net385,
    net386,
    net387,
    net388,
    net389,
    net390,
    net391,
    net392,
    net393,
    net394,
    net395,
    net396,
    net397,
    net398,
    net399,
    net400,
    net401,
    net402,
    net403,
    net404,
    net405,
    net406,
    net407,
    net408,
    net409,
    net410,
    net411,
    net412,
    net413,
    net414,
    net415,
    net416,
    net417,
    net418,
    net419,
    net420,
    net421,
    net422,
    net423,
    net424,
    net425,
    net426,
    net427,
    net428,
    net429}));
 nangate45_64x512_1P_BM \icache.data_mems_6__data_mem.macro_mem  (.we_in(net221),
    .clk(clk_i),
    .ce_in(net233),
    .addr_in({net132,
    net141,
    net150,
    net159,
    net196,
    net205,
    net179,
    net174,
    net117}),
    .rd_out({\icache.data_mems_6__data_mem.data_o [63],
    \icache.data_mems_6__data_mem.data_o [62],
    \icache.data_mems_6__data_mem.data_o [61],
    \icache.data_mems_6__data_mem.data_o [60],
    \icache.data_mems_6__data_mem.data_o [59],
    \icache.data_mems_6__data_mem.data_o [58],
    \icache.data_mems_6__data_mem.data_o [57],
    \icache.data_mems_6__data_mem.data_o [56],
    \icache.data_mems_6__data_mem.data_o [55],
    \icache.data_mems_6__data_mem.data_o [54],
    \icache.data_mems_6__data_mem.data_o [53],
    \icache.data_mems_6__data_mem.data_o [52],
    \icache.data_mems_6__data_mem.data_o [51],
    \icache.data_mems_6__data_mem.data_o [50],
    \icache.data_mems_6__data_mem.data_o [49],
    \icache.data_mems_6__data_mem.data_o [48],
    \icache.data_mems_6__data_mem.data_o [47],
    \icache.data_mems_6__data_mem.data_o [46],
    \icache.data_mems_6__data_mem.data_o [45],
    \icache.data_mems_6__data_mem.data_o [44],
    \icache.data_mems_6__data_mem.data_o [43],
    \icache.data_mems_6__data_mem.data_o [42],
    \icache.data_mems_6__data_mem.data_o [41],
    \icache.data_mems_6__data_mem.data_o [40],
    \icache.data_mems_6__data_mem.data_o [39],
    \icache.data_mems_6__data_mem.data_o [38],
    \icache.data_mems_6__data_mem.data_o [37],
    \icache.data_mems_6__data_mem.data_o [36],
    \icache.data_mems_6__data_mem.data_o [35],
    \icache.data_mems_6__data_mem.data_o [34],
    \icache.data_mems_6__data_mem.data_o [33],
    \icache.data_mems_6__data_mem.data_o [32],
    \icache.data_mems_6__data_mem.data_o [31],
    \icache.data_mems_6__data_mem.data_o [30],
    \icache.data_mems_6__data_mem.data_o [29],
    \icache.data_mems_6__data_mem.data_o [28],
    \icache.data_mems_6__data_mem.data_o [27],
    \icache.data_mems_6__data_mem.data_o [26],
    \icache.data_mems_6__data_mem.data_o [25],
    \icache.data_mems_6__data_mem.data_o [24],
    \icache.data_mems_6__data_mem.data_o [23],
    \icache.data_mems_6__data_mem.data_o [22],
    \icache.data_mems_6__data_mem.data_o [21],
    \icache.data_mems_6__data_mem.data_o [20],
    \icache.data_mems_6__data_mem.data_o [19],
    \icache.data_mems_6__data_mem.data_o [18],
    \icache.data_mems_6__data_mem.data_o [17],
    \icache.data_mems_6__data_mem.data_o [16],
    \icache.data_mems_6__data_mem.data_o [15],
    \icache.data_mems_6__data_mem.data_o [14],
    \icache.data_mems_6__data_mem.data_o [13],
    \icache.data_mems_6__data_mem.data_o [12],
    \icache.data_mems_6__data_mem.data_o [11],
    \icache.data_mems_6__data_mem.data_o [10],
    \icache.data_mems_6__data_mem.data_o [9],
    \icache.data_mems_6__data_mem.data_o [8],
    \icache.data_mems_6__data_mem.data_o [7],
    \icache.data_mems_6__data_mem.data_o [6],
    \icache.data_mems_6__data_mem.data_o [5],
    \icache.data_mems_6__data_mem.data_o [4],
    \icache.data_mems_6__data_mem.data_o [3],
    \icache.data_mems_6__data_mem.data_o [2],
    \icache.data_mems_6__data_mem.data_o [1],
    \icache.data_mems_6__data_mem.data_o [0]}),
    .w_mask_in({_NC385,
    _NC386,
    _NC387,
    _NC388,
    _NC389,
    _NC390,
    _NC391,
    _NC392,
    _NC393,
    _NC394,
    _NC395,
    _NC396,
    _NC397,
    _NC398,
    _NC399,
    _NC400,
    _NC401,
    _NC402,
    _NC403,
    _NC404,
    _NC405,
    _NC406,
    _NC407,
    _NC408,
    _NC409,
    _NC410,
    _NC411,
    _NC412,
    _NC413,
    _NC414,
    _NC415,
    _NC416,
    _NC417,
    _NC418,
    _NC419,
    _NC420,
    _NC421,
    _NC422,
    _NC423,
    _NC424,
    _NC425,
    _NC426,
    _NC427,
    _NC428,
    _NC429,
    _NC430,
    _NC431,
    _NC432,
    _NC433,
    _NC434,
    _NC435,
    _NC436,
    _NC437,
    _NC438,
    _NC439,
    _NC440,
    _NC441,
    _NC442,
    _NC443,
    _NC444,
    _NC445,
    _NC446,
    _NC447,
    _NC448}),
    .wd_in({net302,
    net303,
    net304,
    net305,
    net306,
    net307,
    net308,
    net309,
    net310,
    net311,
    net312,
    net313,
    net314,
    net315,
    net316,
    net317,
    net318,
    net319,
    net320,
    net321,
    net322,
    net323,
    net324,
    net325,
    net326,
    net327,
    net328,
    net329,
    net330,
    net331,
    net332,
    net333,
    net334,
    net335,
    net336,
    net337,
    net338,
    net339,
    net340,
    net341,
    net342,
    net343,
    net344,
    net345,
    net346,
    net347,
    net348,
    net349,
    net350,
    net351,
    net352,
    net353,
    net354,
    net355,
    net356,
    net357,
    net358,
    net359,
    net360,
    net361,
    net362,
    net363,
    net364,
    net365}));
 nangate45_64x512_1P_BM \icache.data_mems_7__data_mem.macro_mem  (.we_in(net220),
    .clk(clk_i),
    .ce_in(net232),
    .addr_in({net131,
    net140,
    net149,
    net158,
    net195,
    net204,
    net178,
    net173,
    net122}),
    .rd_out({\icache.data_mems_7__data_mem.data_o [63],
    \icache.data_mems_7__data_mem.data_o [62],
    \icache.data_mems_7__data_mem.data_o [61],
    \icache.data_mems_7__data_mem.data_o [60],
    \icache.data_mems_7__data_mem.data_o [59],
    \icache.data_mems_7__data_mem.data_o [58],
    \icache.data_mems_7__data_mem.data_o [57],
    \icache.data_mems_7__data_mem.data_o [56],
    \icache.data_mems_7__data_mem.data_o [55],
    \icache.data_mems_7__data_mem.data_o [54],
    \icache.data_mems_7__data_mem.data_o [53],
    \icache.data_mems_7__data_mem.data_o [52],
    \icache.data_mems_7__data_mem.data_o [51],
    \icache.data_mems_7__data_mem.data_o [50],
    \icache.data_mems_7__data_mem.data_o [49],
    \icache.data_mems_7__data_mem.data_o [48],
    \icache.data_mems_7__data_mem.data_o [47],
    \icache.data_mems_7__data_mem.data_o [46],
    \icache.data_mems_7__data_mem.data_o [45],
    \icache.data_mems_7__data_mem.data_o [44],
    \icache.data_mems_7__data_mem.data_o [43],
    \icache.data_mems_7__data_mem.data_o [42],
    \icache.data_mems_7__data_mem.data_o [41],
    \icache.data_mems_7__data_mem.data_o [40],
    \icache.data_mems_7__data_mem.data_o [39],
    \icache.data_mems_7__data_mem.data_o [38],
    \icache.data_mems_7__data_mem.data_o [37],
    \icache.data_mems_7__data_mem.data_o [36],
    \icache.data_mems_7__data_mem.data_o [35],
    \icache.data_mems_7__data_mem.data_o [34],
    \icache.data_mems_7__data_mem.data_o [33],
    \icache.data_mems_7__data_mem.data_o [32],
    \icache.data_mems_7__data_mem.data_o [31],
    \icache.data_mems_7__data_mem.data_o [30],
    \icache.data_mems_7__data_mem.data_o [29],
    \icache.data_mems_7__data_mem.data_o [28],
    \icache.data_mems_7__data_mem.data_o [27],
    \icache.data_mems_7__data_mem.data_o [26],
    \icache.data_mems_7__data_mem.data_o [25],
    \icache.data_mems_7__data_mem.data_o [24],
    \icache.data_mems_7__data_mem.data_o [23],
    \icache.data_mems_7__data_mem.data_o [22],
    \icache.data_mems_7__data_mem.data_o [21],
    \icache.data_mems_7__data_mem.data_o [20],
    \icache.data_mems_7__data_mem.data_o [19],
    \icache.data_mems_7__data_mem.data_o [18],
    \icache.data_mems_7__data_mem.data_o [17],
    \icache.data_mems_7__data_mem.data_o [16],
    \icache.data_mems_7__data_mem.data_o [15],
    \icache.data_mems_7__data_mem.data_o [14],
    \icache.data_mems_7__data_mem.data_o [13],
    \icache.data_mems_7__data_mem.data_o [12],
    \icache.data_mems_7__data_mem.data_o [11],
    \icache.data_mems_7__data_mem.data_o [10],
    \icache.data_mems_7__data_mem.data_o [9],
    \icache.data_mems_7__data_mem.data_o [8],
    \icache.data_mems_7__data_mem.data_o [7],
    \icache.data_mems_7__data_mem.data_o [6],
    \icache.data_mems_7__data_mem.data_o [5],
    \icache.data_mems_7__data_mem.data_o [4],
    \icache.data_mems_7__data_mem.data_o [3],
    \icache.data_mems_7__data_mem.data_o [2],
    \icache.data_mems_7__data_mem.data_o [1],
    \icache.data_mems_7__data_mem.data_o [0]}),
    .w_mask_in({_NC449,
    _NC450,
    _NC451,
    _NC452,
    _NC453,
    _NC454,
    _NC455,
    _NC456,
    _NC457,
    _NC458,
    _NC459,
    _NC460,
    _NC461,
    _NC462,
    _NC463,
    _NC464,
    _NC465,
    _NC466,
    _NC467,
    _NC468,
    _NC469,
    _NC470,
    _NC471,
    _NC472,
    _NC473,
    _NC474,
    _NC475,
    _NC476,
    _NC477,
    _NC478,
    _NC479,
    _NC480,
    _NC481,
    _NC482,
    _NC483,
    _NC484,
    _NC485,
    _NC486,
    _NC487,
    _NC488,
    _NC489,
    _NC490,
    _NC491,
    _NC492,
    _NC493,
    _NC494,
    _NC495,
    _NC496,
    _NC497,
    _NC498,
    _NC499,
    _NC500,
    _NC501,
    _NC502,
    _NC503,
    _NC504,
    _NC505,
    _NC506,
    _NC507,
    _NC508,
    _NC509,
    _NC510,
    _NC511,
    _NC512}),
    .wd_in({net238,
    net239,
    net240,
    net241,
    net242,
    net243,
    net244,
    net245,
    net246,
    net247,
    net248,
    net249,
    net250,
    net251,
    net252,
    net253,
    net254,
    net255,
    net256,
    net257,
    net258,
    net259,
    net260,
    net261,
    net262,
    net263,
    net264,
    net265,
    net266,
    net267,
    net268,
    net269,
    net270,
    net271,
    net272,
    net273,
    net274,
    net275,
    net276,
    net277,
    net278,
    net279,
    net280,
    net281,
    net282,
    net283,
    net284,
    net285,
    net286,
    net287,
    net288,
    net289,
    net290,
    net291,
    net292,
    net293,
    net294,
    net295,
    net296,
    net297,
    net298,
    net299,
    net300,
    net301}));
 nangate45_8x64_1P_bit \icache.stat_mem.macro_mem  (.we_in(net993),
    .clk(clk_i),
    .ce_in(net1003),
    .addr_in({net1085,
    net1086,
    net1087,
    net1088,
    net1089,
    net1090}),
    .rd_out({_32505_,
    \icache.lru_encoder.lru_i [6],
    \icache.lru_encoder.lru_i [5],
    \icache.lru_encoder.lru_i [4],
    \icache.lru_encoder.lru_i [3],
    \icache.lru_encoder.lru_i [2],
    \icache.lru_encoder.lru_i [1],
    \icache.lru_encode [2]}),
    .w_mask_in({_NC513,
    net998,
    net1002,
    \icache.stat_mem.w_mask_i [4],
    net996,
    net999,
    net997,
    _NC514}),
    .wd_in({_NC515,
    net1000,
    \icache.stat_mem.data_i [5],
    net1004,
    net994,
    \icache.stat_mem.data_i [2],
    net995,
    \icache.stat_mem.data_i [0]}));
 nangate45_120x64_1P_bit \icache.tag_mem.macro_mem0  (.we_in(net237),
    .clk(clk_i),
    .ce_in(net224),
    .addr_in({net181,
    net183,
    net185,
    net187,
    net207,
    net209}),
    .rd_out({_32513_,
    _32512_,
    _32511_,
    _32510_,
    \icache.tag_mem.data_o [115],
    \icache.tag_mem.data_o [114],
    \icache.tag_mem.data_o [113],
    \icache.tag_mem.data_o [112],
    \icache.tag_mem.data_o [111],
    \icache.tag_mem.data_o [110],
    \icache.tag_mem.data_o [109],
    \icache.tag_mem.data_o [108],
    \icache.tag_mem.data_o [107],
    \icache.tag_mem.data_o [106],
    \icache.tag_mem.data_o [105],
    \icache.tag_mem.data_o [104],
    \icache.tag_mem.data_o [103],
    \icache.tag_mem.data_o [102],
    \icache.tag_mem.data_o [101],
    \icache.tag_mem.data_o [100],
    \icache.tag_mem.data_o [99],
    \icache.tag_mem.data_o [98],
    \icache.tag_mem.data_o [97],
    \icache.tag_mem.data_o [96],
    \icache.tag_mem.data_o [95],
    \icache.tag_mem.data_o [94],
    \icache.tag_mem.data_o [93],
    \icache.tag_mem.data_o [92],
    \icache.tag_mem.data_o [91],
    \icache.tag_mem.data_o [90],
    \icache.tag_mem.data_o [89],
    \icache.tag_mem.data_o [88],
    \icache.tag_mem.data_o [87],
    \icache.tag_mem.data_o [86],
    \icache.tag_mem.data_o [85],
    \icache.tag_mem.data_o [84],
    \icache.tag_mem.data_o [83],
    \icache.tag_mem.data_o [82],
    \icache.tag_mem.data_o [81],
    \icache.tag_mem.data_o [80],
    \icache.tag_mem.data_o [79],
    \icache.tag_mem.data_o [78],
    \icache.tag_mem.data_o [77],
    \icache.tag_mem.data_o [76],
    \icache.tag_mem.data_o [75],
    \icache.tag_mem.data_o [74],
    \icache.tag_mem.data_o [73],
    \icache.tag_mem.data_o [72],
    \icache.tag_mem.data_o [71],
    \icache.tag_mem.data_o [70],
    \icache.tag_mem.data_o [69],
    \icache.tag_mem.data_o [68],
    \icache.tag_mem.data_o [67],
    \icache.tag_mem.data_o [66],
    \icache.tag_mem.data_o [65],
    \icache.tag_mem.data_o [64],
    \icache.tag_mem.data_o [63],
    \icache.tag_mem.data_o [62],
    \icache.tag_mem.data_o [61],
    \icache.tag_mem.data_o [60],
    \icache.tag_mem.data_o [59],
    \icache.tag_mem.data_o [58],
    \icache.tag_mem.data_o [57],
    \icache.tag_mem.data_o [56],
    \icache.tag_mem.data_o [55],
    \icache.tag_mem.data_o [54],
    \icache.tag_mem.data_o [53],
    \icache.tag_mem.data_o [52],
    \icache.tag_mem.data_o [51],
    \icache.tag_mem.data_o [50],
    \icache.tag_mem.data_o [49],
    \icache.tag_mem.data_o [48],
    \icache.tag_mem.data_o [47],
    \icache.tag_mem.data_o [46],
    \icache.tag_mem.data_o [45],
    \icache.tag_mem.data_o [44],
    \icache.tag_mem.data_o [43],
    \icache.tag_mem.data_o [42],
    \icache.tag_mem.data_o [41],
    \icache.tag_mem.data_o [40],
    \icache.tag_mem.data_o [39],
    \icache.tag_mem.data_o [38],
    \icache.tag_mem.data_o [37],
    \icache.tag_mem.data_o [36],
    \icache.tag_mem.data_o [35],
    \icache.tag_mem.data_o [34],
    \icache.tag_mem.data_o [33],
    \icache.tag_mem.data_o [32],
    \icache.tag_mem.data_o [31],
    \icache.tag_mem.data_o [30],
    \icache.tag_mem.data_o [29],
    \icache.tag_mem.data_o [28],
    \icache.tag_mem.data_o [27],
    \icache.tag_mem.data_o [26],
    \icache.tag_mem.data_o [25],
    \icache.tag_mem.data_o [24],
    \icache.tag_mem.data_o [23],
    \icache.tag_mem.data_o [22],
    \icache.tag_mem.data_o [21],
    \icache.tag_mem.data_o [20],
    \icache.tag_mem.data_o [19],
    \icache.tag_mem.data_o [18],
    \icache.tag_mem.data_o [17],
    \icache.tag_mem.data_o [16],
    \icache.tag_mem.data_o [15],
    \icache.tag_mem.data_o [14],
    \icache.tag_mem.data_o [13],
    \icache.tag_mem.data_o [12],
    \icache.tag_mem.data_o [11],
    \icache.tag_mem.data_o [10],
    \icache.tag_mem.data_o [9],
    \icache.tag_mem.data_o [8],
    \icache.tag_mem.data_o [7],
    \icache.tag_mem.data_o [6],
    \icache.tag_mem.data_o [5],
    \icache.tag_mem.data_o [4],
    \icache.tag_mem.data_o [3],
    \icache.tag_mem.data_o [2],
    \icache.tag_mem.data_o [1],
    \icache.tag_mem.data_o [0]}),
    .w_mask_in({_NC516,
    _NC517,
    _NC518,
    _NC519,
    net780,
    net781,
    net796,
    net795,
    net794,
    net793,
    net792,
    net791,
    net790,
    net789,
    net788,
    net787,
    net786,
    net785,
    net784,
    net783,
    net808,
    net809,
    net807,
    net806,
    net805,
    net804,
    net803,
    net802,
    net801,
    net800,
    net799,
    net798,
    net797,
    net810,
    net811,
    net838,
    net839,
    net837,
    net836,
    net835,
    net834,
    net833,
    net832,
    net831,
    net830,
    net829,
    net828,
    net827,
    net826,
    net825,
    net824,
    net823,
    net822,
    net821,
    net820,
    net819,
    net818,
    net817,
    net816,
    net815,
    net814,
    net813,
    net840,
    net841,
    net868,
    net869,
    net867,
    net866,
    net865,
    net864,
    net863,
    net862,
    net861,
    net860,
    net859,
    net858,
    net857,
    net856,
    net855,
    net854,
    net853,
    net852,
    net851,
    net850,
    net849,
    net848,
    net847,
    net846,
    net845,
    net844,
    net843,
    net991,
    net992,
    net889,
    net888,
    net887,
    net886,
    net885,
    net884,
    net883,
    net881,
    net880,
    net879,
    net878,
    net877,
    net876,
    net875,
    net874,
    net873,
    net872,
    net896,
    net897,
    net895,
    net894,
    net893,
    net892,
    net891,
    net890,
    net882,
    net871}),
    .wd_in({_NC520,
    _NC521,
    _NC522,
    _NC523,
    net1091,
    net1099,
    net1217,
    net1226,
    net1107,
    net1235,
    net1244,
    net1253,
    net1116,
    net1125,
    net1133,
    net1142,
    net1005,
    net1013,
    net1151,
    net1160,
    net1024,
    net1032,
    net1172,
    net1039,
    net1048,
    net1181,
    net1190,
    net1056,
    net1064,
    net1072,
    net1199,
    net1080,
    net1208,
    net1094,
    net1102,
    net1220,
    net1229,
    net1110,
    net1238,
    net1247,
    net1256,
    net1119,
    net1128,
    net1136,
    net1145,
    net1008,
    net1016,
    net1154,
    net1163,
    net1023,
    net1031,
    net1171,
    net1038,
    net1046,
    net1179,
    net1188,
    net1055,
    net1063,
    net1071,
    net1198,
    net1079,
    net1207,
    net1093,
    net1101,
    net1219,
    net1228,
    net1109,
    net1237,
    net1246,
    net1255,
    net1118,
    net1127,
    net1135,
    net1144,
    net1007,
    net1015,
    net1153,
    net1162,
    net1022,
    net1030,
    net1170,
    net1037,
    net1045,
    net1178,
    net1187,
    net1053,
    net1061,
    net1069,
    net1197,
    net1078,
    net1206,
    net1092,
    net1100,
    net1218,
    net1227,
    net1108,
    net1236,
    net1245,
    net1254,
    net1117,
    net1126,
    net1134,
    net1143,
    net1006,
    net1014,
    net1152,
    net1161,
    net1021,
    net1029,
    net1169,
    net1040,
    net1047,
    net1180,
    net1189,
    net1054,
    net1062,
    net1070,
    net1196,
    net1077,
    net1205}));
 nangate45_120x64_1P_bit \icache.tag_mem.macro_mem1  (.we_in(net236),
    .clk(clk_i),
    .ce_in(net223),
    .addr_in({net180,
    net182,
    net184,
    net186,
    net206,
    net208}),
    .rd_out({_32509_,
    _32508_,
    _32507_,
    _32506_,
    \icache.tag_mem.data_o [231],
    \icache.tag_mem.data_o [230],
    \icache.tag_mem.data_o [229],
    \icache.tag_mem.data_o [228],
    \icache.tag_mem.data_o [227],
    \icache.tag_mem.data_o [226],
    \icache.tag_mem.data_o [225],
    \icache.tag_mem.data_o [224],
    \icache.tag_mem.data_o [223],
    \icache.tag_mem.data_o [222],
    \icache.tag_mem.data_o [221],
    \icache.tag_mem.data_o [220],
    \icache.tag_mem.data_o [219],
    \icache.tag_mem.data_o [218],
    \icache.tag_mem.data_o [217],
    \icache.tag_mem.data_o [216],
    \icache.tag_mem.data_o [215],
    \icache.tag_mem.data_o [214],
    \icache.tag_mem.data_o [213],
    \icache.tag_mem.data_o [212],
    \icache.tag_mem.data_o [211],
    \icache.tag_mem.data_o [210],
    \icache.tag_mem.data_o [209],
    \icache.tag_mem.data_o [208],
    \icache.tag_mem.data_o [207],
    \icache.tag_mem.data_o [206],
    \icache.tag_mem.data_o [205],
    \icache.tag_mem.data_o [204],
    \icache.tag_mem.data_o [203],
    \icache.tag_mem.data_o [202],
    \icache.tag_mem.data_o [201],
    \icache.tag_mem.data_o [200],
    \icache.tag_mem.data_o [199],
    \icache.tag_mem.data_o [198],
    \icache.tag_mem.data_o [197],
    \icache.tag_mem.data_o [196],
    \icache.tag_mem.data_o [195],
    \icache.tag_mem.data_o [194],
    \icache.tag_mem.data_o [193],
    \icache.tag_mem.data_o [192],
    \icache.tag_mem.data_o [191],
    \icache.tag_mem.data_o [190],
    \icache.tag_mem.data_o [189],
    \icache.tag_mem.data_o [188],
    \icache.tag_mem.data_o [187],
    \icache.tag_mem.data_o [186],
    \icache.tag_mem.data_o [185],
    \icache.tag_mem.data_o [184],
    \icache.tag_mem.data_o [183],
    \icache.tag_mem.data_o [182],
    \icache.tag_mem.data_o [181],
    \icache.tag_mem.data_o [180],
    \icache.tag_mem.data_o [179],
    \icache.tag_mem.data_o [178],
    \icache.tag_mem.data_o [177],
    \icache.tag_mem.data_o [176],
    \icache.tag_mem.data_o [175],
    \icache.tag_mem.data_o [174],
    \icache.tag_mem.data_o [173],
    \icache.tag_mem.data_o [172],
    \icache.tag_mem.data_o [171],
    \icache.tag_mem.data_o [170],
    \icache.tag_mem.data_o [169],
    \icache.tag_mem.data_o [168],
    \icache.tag_mem.data_o [167],
    \icache.tag_mem.data_o [166],
    \icache.tag_mem.data_o [165],
    \icache.tag_mem.data_o [164],
    \icache.tag_mem.data_o [163],
    \icache.tag_mem.data_o [162],
    \icache.tag_mem.data_o [161],
    \icache.tag_mem.data_o [160],
    \icache.tag_mem.data_o [159],
    \icache.tag_mem.data_o [158],
    \icache.tag_mem.data_o [157],
    \icache.tag_mem.data_o [156],
    \icache.tag_mem.data_o [155],
    \icache.tag_mem.data_o [154],
    \icache.tag_mem.data_o [153],
    \icache.tag_mem.data_o [152],
    \icache.tag_mem.data_o [151],
    \icache.tag_mem.data_o [150],
    \icache.tag_mem.data_o [149],
    \icache.tag_mem.data_o [148],
    \icache.tag_mem.data_o [147],
    \icache.tag_mem.data_o [146],
    \icache.tag_mem.data_o [145],
    \icache.tag_mem.data_o [144],
    \icache.tag_mem.data_o [143],
    \icache.tag_mem.data_o [142],
    \icache.tag_mem.data_o [141],
    \icache.tag_mem.data_o [140],
    \icache.tag_mem.data_o [139],
    \icache.tag_mem.data_o [138],
    \icache.tag_mem.data_o [137],
    \icache.tag_mem.data_o [136],
    \icache.tag_mem.data_o [135],
    \icache.tag_mem.data_o [134],
    \icache.tag_mem.data_o [133],
    \icache.tag_mem.data_o [132],
    \icache.tag_mem.data_o [131],
    \icache.tag_mem.data_o [130],
    \icache.tag_mem.data_o [129],
    \icache.tag_mem.data_o [128],
    \icache.tag_mem.data_o [127],
    \icache.tag_mem.data_o [126],
    \icache.tag_mem.data_o [125],
    \icache.tag_mem.data_o [124],
    \icache.tag_mem.data_o [123],
    \icache.tag_mem.data_o [122],
    \icache.tag_mem.data_o [121],
    \icache.tag_mem.data_o [120],
    \icache.tag_mem.data_o [119],
    \icache.tag_mem.data_o [118],
    \icache.tag_mem.data_o [117],
    \icache.tag_mem.data_o [116]}),
    .w_mask_in({_NC524,
    _NC525,
    _NC526,
    _NC527,
    net898,
    net899,
    net914,
    net913,
    net912,
    net911,
    net910,
    net909,
    net908,
    net907,
    net906,
    net905,
    net904,
    net903,
    net902,
    net901,
    net926,
    net927,
    net925,
    net924,
    net923,
    net922,
    net921,
    net920,
    net919,
    net918,
    net917,
    net916,
    net915,
    net959,
    net960,
    net987,
    net988,
    net986,
    net985,
    net984,
    net983,
    net982,
    net981,
    net980,
    net979,
    net978,
    net977,
    net976,
    net975,
    net974,
    net973,
    net972,
    net971,
    net970,
    net969,
    net968,
    net967,
    net966,
    net965,
    net964,
    net963,
    net962,
    net928,
    net929,
    net956,
    net957,
    net955,
    net954,
    net953,
    net952,
    net951,
    net950,
    net949,
    net948,
    net947,
    net946,
    net945,
    net944,
    net943,
    net942,
    net941,
    net940,
    net939,
    net938,
    net937,
    net936,
    net935,
    net934,
    net933,
    net932,
    net931,
    net750,
    net751,
    net771,
    net770,
    net769,
    net768,
    net767,
    net766,
    net765,
    net763,
    net762,
    net761,
    net760,
    net759,
    net758,
    net757,
    net756,
    net755,
    net754,
    net778,
    net779,
    net777,
    net776,
    net775,
    net774,
    net773,
    net772,
    net764,
    net753}),
    .wd_in({_NC528,
    _NC529,
    _NC530,
    _NC531,
    net1095,
    net1103,
    net1221,
    net1230,
    net1111,
    net1239,
    net1248,
    net1257,
    net1120,
    net1129,
    net1137,
    net1146,
    net1009,
    net1017,
    net1155,
    net1164,
    net1027,
    net1035,
    net1175,
    net1044,
    net1051,
    net1184,
    net1193,
    net1059,
    net1067,
    net1075,
    net1202,
    net1083,
    net1211,
    net1097,
    net1105,
    net1223,
    net1232,
    net1113,
    net1241,
    net1250,
    net1259,
    net1122,
    net1131,
    net1139,
    net1148,
    net1011,
    net1019,
    net1157,
    net1166,
    net1028,
    net1036,
    net1176,
    net1042,
    net1050,
    net1183,
    net1192,
    net1060,
    net1068,
    net1076,
    net1203,
    net1084,
    net1212,
    net1098,
    net1106,
    net1224,
    net1233,
    net1114,
    net1242,
    net1251,
    net1260,
    net1123,
    net1132,
    net1140,
    net1149,
    net1012,
    net1020,
    net1158,
    net1167,
    net1026,
    net1034,
    net1174,
    net1041,
    net1049,
    net1182,
    net1191,
    net1057,
    net1065,
    net1073,
    net1201,
    net1082,
    net1210,
    net1096,
    net1104,
    net1222,
    net1231,
    net1112,
    net1240,
    net1249,
    net1258,
    net1121,
    net1130,
    net1138,
    net1147,
    net1010,
    net1018,
    net1156,
    net1165,
    net1025,
    net1033,
    net1173,
    net1043,
    net1052,
    net1185,
    net1194,
    net1058,
    net1066,
    net1074,
    net1200,
    net1081,
    net1209}));
endmodule
