module nangate45_120x64_1P_bit
(
   rd_out,
   addr_in,
   we_in,
   wd_in,
   w_mask_in,
   clk,
   ce_in
);
   parameter                BITS = 120;
   parameter                WORD_DEPTH = 64;
   parameter                ADDR_WIDTH = 6;
   parameter                corrupt_mem_on_X_p = 1;

   output reg [BITS-1:0]    rd_out;
   input  [ADDR_WIDTH-1:0]  addr_in;
   input                    we_in;
   input  [BITS-1:0]        wd_in;
   input  [BITS-1:0]        w_mask_in;
   input                    clk;
   input                    ce_in;

endmodule

module nangate45_64x512_1P_BM
(
   rd_out,
   addr_in,
   we_in,
   wd_in,
   w_mask_in,
   clk,
   ce_in
);
   parameter                BITS = 64;
   parameter                WORD_DEPTH = 512;
   parameter                ADDR_WIDTH = 9;
   parameter                corrupt_mem_on_X_p = 1;

   output reg [BITS-1:0]    rd_out;
   input  [ADDR_WIDTH-1:0]  addr_in;
   input                    we_in;
   input  [BITS-1:0]        wd_in;
   input  [BITS-1:0]        w_mask_in;
   input                    clk;
   input                    ce_in;

endmodule

module nangate45_8x64_1P_bit
(
   rd_out,
   addr_in,
   we_in,
   wd_in,
   w_mask_in,
   clk,
   ce_in
);
   parameter                BITS = 8;
   parameter                WORD_DEPTH = 64;
   parameter                ADDR_WIDTH = 6;
   parameter                corrupt_mem_on_X_p = 1;

   output reg [BITS-1:0]    rd_out;
   input  [ADDR_WIDTH-1:0]  addr_in;
   input                    we_in;
   input  [BITS-1:0]        wd_in;
   input  [BITS-1:0]        w_mask_in;
   input                    clk;
   input                    ce_in;

endmodule

module bsg_dff_reset_en_width_p27
(
  clk_i,
  reset_i,
  en_i,
  data_i,
  data_o
);

  input [26:0] data_i;
  output [26:0] data_o;
  input clk_i;
  input reset_i;
  input en_i;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32;
  reg [26:0] data_o;
  assign N3 = (N0)? 1'b1 : 
              (N32)? 1'b1 : 
              (N2)? 1'b0 : 1'b0;
  assign N0 = reset_i;
  assign { N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4 } = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                               (N32)? data_i : 1'b0;
  assign N1 = en_i | reset_i;
  assign N2 = ~N1;
  assign N31 = ~reset_i;
  assign N32 = en_i & N31;

  always @(posedge clk_i) begin
    if(N3) begin
      { data_o[26:0] } <= { N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4 };
    end 
  end


endmodule



module bsg_mem_1r1w_synth_width_p49_els_p64_read_write_same_addr_p0_harden_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [5:0] w_addr_i;
  input [48:0] w_data_i;
  input [5:0] r_addr_i;
  output [48:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [48:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294;
  reg [3135:0] mem;
  assign r_data_o[48] = (N76)? mem[48] : 
                        (N78)? mem[97] : 
                        (N80)? mem[146] : 
                        (N82)? mem[195] : 
                        (N84)? mem[244] : 
                        (N86)? mem[293] : 
                        (N88)? mem[342] : 
                        (N90)? mem[391] : 
                        (N92)? mem[440] : 
                        (N94)? mem[489] : 
                        (N96)? mem[538] : 
                        (N98)? mem[587] : 
                        (N100)? mem[636] : 
                        (N102)? mem[685] : 
                        (N104)? mem[734] : 
                        (N106)? mem[783] : 
                        (N108)? mem[832] : 
                        (N110)? mem[881] : 
                        (N112)? mem[930] : 
                        (N114)? mem[979] : 
                        (N116)? mem[1028] : 
                        (N118)? mem[1077] : 
                        (N120)? mem[1126] : 
                        (N122)? mem[1175] : 
                        (N124)? mem[1224] : 
                        (N126)? mem[1273] : 
                        (N128)? mem[1322] : 
                        (N130)? mem[1371] : 
                        (N132)? mem[1420] : 
                        (N134)? mem[1469] : 
                        (N136)? mem[1518] : 
                        (N138)? mem[1567] : 
                        (N77)? mem[1616] : 
                        (N79)? mem[1665] : 
                        (N81)? mem[1714] : 
                        (N83)? mem[1763] : 
                        (N85)? mem[1812] : 
                        (N87)? mem[1861] : 
                        (N89)? mem[1910] : 
                        (N91)? mem[1959] : 
                        (N93)? mem[2008] : 
                        (N95)? mem[2057] : 
                        (N97)? mem[2106] : 
                        (N99)? mem[2155] : 
                        (N101)? mem[2204] : 
                        (N103)? mem[2253] : 
                        (N105)? mem[2302] : 
                        (N107)? mem[2351] : 
                        (N109)? mem[2400] : 
                        (N111)? mem[2449] : 
                        (N113)? mem[2498] : 
                        (N115)? mem[2547] : 
                        (N117)? mem[2596] : 
                        (N119)? mem[2645] : 
                        (N121)? mem[2694] : 
                        (N123)? mem[2743] : 
                        (N125)? mem[2792] : 
                        (N127)? mem[2841] : 
                        (N129)? mem[2890] : 
                        (N131)? mem[2939] : 
                        (N133)? mem[2988] : 
                        (N135)? mem[3037] : 
                        (N137)? mem[3086] : 
                        (N139)? mem[3135] : 1'b0;
  assign r_data_o[47] = (N76)? mem[47] : 
                        (N78)? mem[96] : 
                        (N80)? mem[145] : 
                        (N82)? mem[194] : 
                        (N84)? mem[243] : 
                        (N86)? mem[292] : 
                        (N88)? mem[341] : 
                        (N90)? mem[390] : 
                        (N92)? mem[439] : 
                        (N94)? mem[488] : 
                        (N96)? mem[537] : 
                        (N98)? mem[586] : 
                        (N100)? mem[635] : 
                        (N102)? mem[684] : 
                        (N104)? mem[733] : 
                        (N106)? mem[782] : 
                        (N108)? mem[831] : 
                        (N110)? mem[880] : 
                        (N112)? mem[929] : 
                        (N114)? mem[978] : 
                        (N116)? mem[1027] : 
                        (N118)? mem[1076] : 
                        (N120)? mem[1125] : 
                        (N122)? mem[1174] : 
                        (N124)? mem[1223] : 
                        (N126)? mem[1272] : 
                        (N128)? mem[1321] : 
                        (N130)? mem[1370] : 
                        (N132)? mem[1419] : 
                        (N134)? mem[1468] : 
                        (N136)? mem[1517] : 
                        (N138)? mem[1566] : 
                        (N77)? mem[1615] : 
                        (N79)? mem[1664] : 
                        (N81)? mem[1713] : 
                        (N83)? mem[1762] : 
                        (N85)? mem[1811] : 
                        (N87)? mem[1860] : 
                        (N89)? mem[1909] : 
                        (N91)? mem[1958] : 
                        (N93)? mem[2007] : 
                        (N95)? mem[2056] : 
                        (N97)? mem[2105] : 
                        (N99)? mem[2154] : 
                        (N101)? mem[2203] : 
                        (N103)? mem[2252] : 
                        (N105)? mem[2301] : 
                        (N107)? mem[2350] : 
                        (N109)? mem[2399] : 
                        (N111)? mem[2448] : 
                        (N113)? mem[2497] : 
                        (N115)? mem[2546] : 
                        (N117)? mem[2595] : 
                        (N119)? mem[2644] : 
                        (N121)? mem[2693] : 
                        (N123)? mem[2742] : 
                        (N125)? mem[2791] : 
                        (N127)? mem[2840] : 
                        (N129)? mem[2889] : 
                        (N131)? mem[2938] : 
                        (N133)? mem[2987] : 
                        (N135)? mem[3036] : 
                        (N137)? mem[3085] : 
                        (N139)? mem[3134] : 1'b0;
  assign r_data_o[46] = (N76)? mem[46] : 
                        (N78)? mem[95] : 
                        (N80)? mem[144] : 
                        (N82)? mem[193] : 
                        (N84)? mem[242] : 
                        (N86)? mem[291] : 
                        (N88)? mem[340] : 
                        (N90)? mem[389] : 
                        (N92)? mem[438] : 
                        (N94)? mem[487] : 
                        (N96)? mem[536] : 
                        (N98)? mem[585] : 
                        (N100)? mem[634] : 
                        (N102)? mem[683] : 
                        (N104)? mem[732] : 
                        (N106)? mem[781] : 
                        (N108)? mem[830] : 
                        (N110)? mem[879] : 
                        (N112)? mem[928] : 
                        (N114)? mem[977] : 
                        (N116)? mem[1026] : 
                        (N118)? mem[1075] : 
                        (N120)? mem[1124] : 
                        (N122)? mem[1173] : 
                        (N124)? mem[1222] : 
                        (N126)? mem[1271] : 
                        (N128)? mem[1320] : 
                        (N130)? mem[1369] : 
                        (N132)? mem[1418] : 
                        (N134)? mem[1467] : 
                        (N136)? mem[1516] : 
                        (N138)? mem[1565] : 
                        (N77)? mem[1614] : 
                        (N79)? mem[1663] : 
                        (N81)? mem[1712] : 
                        (N83)? mem[1761] : 
                        (N85)? mem[1810] : 
                        (N87)? mem[1859] : 
                        (N89)? mem[1908] : 
                        (N91)? mem[1957] : 
                        (N93)? mem[2006] : 
                        (N95)? mem[2055] : 
                        (N97)? mem[2104] : 
                        (N99)? mem[2153] : 
                        (N101)? mem[2202] : 
                        (N103)? mem[2251] : 
                        (N105)? mem[2300] : 
                        (N107)? mem[2349] : 
                        (N109)? mem[2398] : 
                        (N111)? mem[2447] : 
                        (N113)? mem[2496] : 
                        (N115)? mem[2545] : 
                        (N117)? mem[2594] : 
                        (N119)? mem[2643] : 
                        (N121)? mem[2692] : 
                        (N123)? mem[2741] : 
                        (N125)? mem[2790] : 
                        (N127)? mem[2839] : 
                        (N129)? mem[2888] : 
                        (N131)? mem[2937] : 
                        (N133)? mem[2986] : 
                        (N135)? mem[3035] : 
                        (N137)? mem[3084] : 
                        (N139)? mem[3133] : 1'b0;
  assign r_data_o[45] = (N76)? mem[45] : 
                        (N78)? mem[94] : 
                        (N80)? mem[143] : 
                        (N82)? mem[192] : 
                        (N84)? mem[241] : 
                        (N86)? mem[290] : 
                        (N88)? mem[339] : 
                        (N90)? mem[388] : 
                        (N92)? mem[437] : 
                        (N94)? mem[486] : 
                        (N96)? mem[535] : 
                        (N98)? mem[584] : 
                        (N100)? mem[633] : 
                        (N102)? mem[682] : 
                        (N104)? mem[731] : 
                        (N106)? mem[780] : 
                        (N108)? mem[829] : 
                        (N110)? mem[878] : 
                        (N112)? mem[927] : 
                        (N114)? mem[976] : 
                        (N116)? mem[1025] : 
                        (N118)? mem[1074] : 
                        (N120)? mem[1123] : 
                        (N122)? mem[1172] : 
                        (N124)? mem[1221] : 
                        (N126)? mem[1270] : 
                        (N128)? mem[1319] : 
                        (N130)? mem[1368] : 
                        (N132)? mem[1417] : 
                        (N134)? mem[1466] : 
                        (N136)? mem[1515] : 
                        (N138)? mem[1564] : 
                        (N77)? mem[1613] : 
                        (N79)? mem[1662] : 
                        (N81)? mem[1711] : 
                        (N83)? mem[1760] : 
                        (N85)? mem[1809] : 
                        (N87)? mem[1858] : 
                        (N89)? mem[1907] : 
                        (N91)? mem[1956] : 
                        (N93)? mem[2005] : 
                        (N95)? mem[2054] : 
                        (N97)? mem[2103] : 
                        (N99)? mem[2152] : 
                        (N101)? mem[2201] : 
                        (N103)? mem[2250] : 
                        (N105)? mem[2299] : 
                        (N107)? mem[2348] : 
                        (N109)? mem[2397] : 
                        (N111)? mem[2446] : 
                        (N113)? mem[2495] : 
                        (N115)? mem[2544] : 
                        (N117)? mem[2593] : 
                        (N119)? mem[2642] : 
                        (N121)? mem[2691] : 
                        (N123)? mem[2740] : 
                        (N125)? mem[2789] : 
                        (N127)? mem[2838] : 
                        (N129)? mem[2887] : 
                        (N131)? mem[2936] : 
                        (N133)? mem[2985] : 
                        (N135)? mem[3034] : 
                        (N137)? mem[3083] : 
                        (N139)? mem[3132] : 1'b0;
  assign r_data_o[44] = (N76)? mem[44] : 
                        (N78)? mem[93] : 
                        (N80)? mem[142] : 
                        (N82)? mem[191] : 
                        (N84)? mem[240] : 
                        (N86)? mem[289] : 
                        (N88)? mem[338] : 
                        (N90)? mem[387] : 
                        (N92)? mem[436] : 
                        (N94)? mem[485] : 
                        (N96)? mem[534] : 
                        (N98)? mem[583] : 
                        (N100)? mem[632] : 
                        (N102)? mem[681] : 
                        (N104)? mem[730] : 
                        (N106)? mem[779] : 
                        (N108)? mem[828] : 
                        (N110)? mem[877] : 
                        (N112)? mem[926] : 
                        (N114)? mem[975] : 
                        (N116)? mem[1024] : 
                        (N118)? mem[1073] : 
                        (N120)? mem[1122] : 
                        (N122)? mem[1171] : 
                        (N124)? mem[1220] : 
                        (N126)? mem[1269] : 
                        (N128)? mem[1318] : 
                        (N130)? mem[1367] : 
                        (N132)? mem[1416] : 
                        (N134)? mem[1465] : 
                        (N136)? mem[1514] : 
                        (N138)? mem[1563] : 
                        (N77)? mem[1612] : 
                        (N79)? mem[1661] : 
                        (N81)? mem[1710] : 
                        (N83)? mem[1759] : 
                        (N85)? mem[1808] : 
                        (N87)? mem[1857] : 
                        (N89)? mem[1906] : 
                        (N91)? mem[1955] : 
                        (N93)? mem[2004] : 
                        (N95)? mem[2053] : 
                        (N97)? mem[2102] : 
                        (N99)? mem[2151] : 
                        (N101)? mem[2200] : 
                        (N103)? mem[2249] : 
                        (N105)? mem[2298] : 
                        (N107)? mem[2347] : 
                        (N109)? mem[2396] : 
                        (N111)? mem[2445] : 
                        (N113)? mem[2494] : 
                        (N115)? mem[2543] : 
                        (N117)? mem[2592] : 
                        (N119)? mem[2641] : 
                        (N121)? mem[2690] : 
                        (N123)? mem[2739] : 
                        (N125)? mem[2788] : 
                        (N127)? mem[2837] : 
                        (N129)? mem[2886] : 
                        (N131)? mem[2935] : 
                        (N133)? mem[2984] : 
                        (N135)? mem[3033] : 
                        (N137)? mem[3082] : 
                        (N139)? mem[3131] : 1'b0;
  assign r_data_o[43] = (N76)? mem[43] : 
                        (N78)? mem[92] : 
                        (N80)? mem[141] : 
                        (N82)? mem[190] : 
                        (N84)? mem[239] : 
                        (N86)? mem[288] : 
                        (N88)? mem[337] : 
                        (N90)? mem[386] : 
                        (N92)? mem[435] : 
                        (N94)? mem[484] : 
                        (N96)? mem[533] : 
                        (N98)? mem[582] : 
                        (N100)? mem[631] : 
                        (N102)? mem[680] : 
                        (N104)? mem[729] : 
                        (N106)? mem[778] : 
                        (N108)? mem[827] : 
                        (N110)? mem[876] : 
                        (N112)? mem[925] : 
                        (N114)? mem[974] : 
                        (N116)? mem[1023] : 
                        (N118)? mem[1072] : 
                        (N120)? mem[1121] : 
                        (N122)? mem[1170] : 
                        (N124)? mem[1219] : 
                        (N126)? mem[1268] : 
                        (N128)? mem[1317] : 
                        (N130)? mem[1366] : 
                        (N132)? mem[1415] : 
                        (N134)? mem[1464] : 
                        (N136)? mem[1513] : 
                        (N138)? mem[1562] : 
                        (N77)? mem[1611] : 
                        (N79)? mem[1660] : 
                        (N81)? mem[1709] : 
                        (N83)? mem[1758] : 
                        (N85)? mem[1807] : 
                        (N87)? mem[1856] : 
                        (N89)? mem[1905] : 
                        (N91)? mem[1954] : 
                        (N93)? mem[2003] : 
                        (N95)? mem[2052] : 
                        (N97)? mem[2101] : 
                        (N99)? mem[2150] : 
                        (N101)? mem[2199] : 
                        (N103)? mem[2248] : 
                        (N105)? mem[2297] : 
                        (N107)? mem[2346] : 
                        (N109)? mem[2395] : 
                        (N111)? mem[2444] : 
                        (N113)? mem[2493] : 
                        (N115)? mem[2542] : 
                        (N117)? mem[2591] : 
                        (N119)? mem[2640] : 
                        (N121)? mem[2689] : 
                        (N123)? mem[2738] : 
                        (N125)? mem[2787] : 
                        (N127)? mem[2836] : 
                        (N129)? mem[2885] : 
                        (N131)? mem[2934] : 
                        (N133)? mem[2983] : 
                        (N135)? mem[3032] : 
                        (N137)? mem[3081] : 
                        (N139)? mem[3130] : 1'b0;
  assign r_data_o[42] = (N76)? mem[42] : 
                        (N78)? mem[91] : 
                        (N80)? mem[140] : 
                        (N82)? mem[189] : 
                        (N84)? mem[238] : 
                        (N86)? mem[287] : 
                        (N88)? mem[336] : 
                        (N90)? mem[385] : 
                        (N92)? mem[434] : 
                        (N94)? mem[483] : 
                        (N96)? mem[532] : 
                        (N98)? mem[581] : 
                        (N100)? mem[630] : 
                        (N102)? mem[679] : 
                        (N104)? mem[728] : 
                        (N106)? mem[777] : 
                        (N108)? mem[826] : 
                        (N110)? mem[875] : 
                        (N112)? mem[924] : 
                        (N114)? mem[973] : 
                        (N116)? mem[1022] : 
                        (N118)? mem[1071] : 
                        (N120)? mem[1120] : 
                        (N122)? mem[1169] : 
                        (N124)? mem[1218] : 
                        (N126)? mem[1267] : 
                        (N128)? mem[1316] : 
                        (N130)? mem[1365] : 
                        (N132)? mem[1414] : 
                        (N134)? mem[1463] : 
                        (N136)? mem[1512] : 
                        (N138)? mem[1561] : 
                        (N77)? mem[1610] : 
                        (N79)? mem[1659] : 
                        (N81)? mem[1708] : 
                        (N83)? mem[1757] : 
                        (N85)? mem[1806] : 
                        (N87)? mem[1855] : 
                        (N89)? mem[1904] : 
                        (N91)? mem[1953] : 
                        (N93)? mem[2002] : 
                        (N95)? mem[2051] : 
                        (N97)? mem[2100] : 
                        (N99)? mem[2149] : 
                        (N101)? mem[2198] : 
                        (N103)? mem[2247] : 
                        (N105)? mem[2296] : 
                        (N107)? mem[2345] : 
                        (N109)? mem[2394] : 
                        (N111)? mem[2443] : 
                        (N113)? mem[2492] : 
                        (N115)? mem[2541] : 
                        (N117)? mem[2590] : 
                        (N119)? mem[2639] : 
                        (N121)? mem[2688] : 
                        (N123)? mem[2737] : 
                        (N125)? mem[2786] : 
                        (N127)? mem[2835] : 
                        (N129)? mem[2884] : 
                        (N131)? mem[2933] : 
                        (N133)? mem[2982] : 
                        (N135)? mem[3031] : 
                        (N137)? mem[3080] : 
                        (N139)? mem[3129] : 1'b0;
  assign r_data_o[41] = (N76)? mem[41] : 
                        (N78)? mem[90] : 
                        (N80)? mem[139] : 
                        (N82)? mem[188] : 
                        (N84)? mem[237] : 
                        (N86)? mem[286] : 
                        (N88)? mem[335] : 
                        (N90)? mem[384] : 
                        (N92)? mem[433] : 
                        (N94)? mem[482] : 
                        (N96)? mem[531] : 
                        (N98)? mem[580] : 
                        (N100)? mem[629] : 
                        (N102)? mem[678] : 
                        (N104)? mem[727] : 
                        (N106)? mem[776] : 
                        (N108)? mem[825] : 
                        (N110)? mem[874] : 
                        (N112)? mem[923] : 
                        (N114)? mem[972] : 
                        (N116)? mem[1021] : 
                        (N118)? mem[1070] : 
                        (N120)? mem[1119] : 
                        (N122)? mem[1168] : 
                        (N124)? mem[1217] : 
                        (N126)? mem[1266] : 
                        (N128)? mem[1315] : 
                        (N130)? mem[1364] : 
                        (N132)? mem[1413] : 
                        (N134)? mem[1462] : 
                        (N136)? mem[1511] : 
                        (N138)? mem[1560] : 
                        (N77)? mem[1609] : 
                        (N79)? mem[1658] : 
                        (N81)? mem[1707] : 
                        (N83)? mem[1756] : 
                        (N85)? mem[1805] : 
                        (N87)? mem[1854] : 
                        (N89)? mem[1903] : 
                        (N91)? mem[1952] : 
                        (N93)? mem[2001] : 
                        (N95)? mem[2050] : 
                        (N97)? mem[2099] : 
                        (N99)? mem[2148] : 
                        (N101)? mem[2197] : 
                        (N103)? mem[2246] : 
                        (N105)? mem[2295] : 
                        (N107)? mem[2344] : 
                        (N109)? mem[2393] : 
                        (N111)? mem[2442] : 
                        (N113)? mem[2491] : 
                        (N115)? mem[2540] : 
                        (N117)? mem[2589] : 
                        (N119)? mem[2638] : 
                        (N121)? mem[2687] : 
                        (N123)? mem[2736] : 
                        (N125)? mem[2785] : 
                        (N127)? mem[2834] : 
                        (N129)? mem[2883] : 
                        (N131)? mem[2932] : 
                        (N133)? mem[2981] : 
                        (N135)? mem[3030] : 
                        (N137)? mem[3079] : 
                        (N139)? mem[3128] : 1'b0;
  assign r_data_o[40] = (N76)? mem[40] : 
                        (N78)? mem[89] : 
                        (N80)? mem[138] : 
                        (N82)? mem[187] : 
                        (N84)? mem[236] : 
                        (N86)? mem[285] : 
                        (N88)? mem[334] : 
                        (N90)? mem[383] : 
                        (N92)? mem[432] : 
                        (N94)? mem[481] : 
                        (N96)? mem[530] : 
                        (N98)? mem[579] : 
                        (N100)? mem[628] : 
                        (N102)? mem[677] : 
                        (N104)? mem[726] : 
                        (N106)? mem[775] : 
                        (N108)? mem[824] : 
                        (N110)? mem[873] : 
                        (N112)? mem[922] : 
                        (N114)? mem[971] : 
                        (N116)? mem[1020] : 
                        (N118)? mem[1069] : 
                        (N120)? mem[1118] : 
                        (N122)? mem[1167] : 
                        (N124)? mem[1216] : 
                        (N126)? mem[1265] : 
                        (N128)? mem[1314] : 
                        (N130)? mem[1363] : 
                        (N132)? mem[1412] : 
                        (N134)? mem[1461] : 
                        (N136)? mem[1510] : 
                        (N138)? mem[1559] : 
                        (N77)? mem[1608] : 
                        (N79)? mem[1657] : 
                        (N81)? mem[1706] : 
                        (N83)? mem[1755] : 
                        (N85)? mem[1804] : 
                        (N87)? mem[1853] : 
                        (N89)? mem[1902] : 
                        (N91)? mem[1951] : 
                        (N93)? mem[2000] : 
                        (N95)? mem[2049] : 
                        (N97)? mem[2098] : 
                        (N99)? mem[2147] : 
                        (N101)? mem[2196] : 
                        (N103)? mem[2245] : 
                        (N105)? mem[2294] : 
                        (N107)? mem[2343] : 
                        (N109)? mem[2392] : 
                        (N111)? mem[2441] : 
                        (N113)? mem[2490] : 
                        (N115)? mem[2539] : 
                        (N117)? mem[2588] : 
                        (N119)? mem[2637] : 
                        (N121)? mem[2686] : 
                        (N123)? mem[2735] : 
                        (N125)? mem[2784] : 
                        (N127)? mem[2833] : 
                        (N129)? mem[2882] : 
                        (N131)? mem[2931] : 
                        (N133)? mem[2980] : 
                        (N135)? mem[3029] : 
                        (N137)? mem[3078] : 
                        (N139)? mem[3127] : 1'b0;
  assign r_data_o[39] = (N76)? mem[39] : 
                        (N78)? mem[88] : 
                        (N80)? mem[137] : 
                        (N82)? mem[186] : 
                        (N84)? mem[235] : 
                        (N86)? mem[284] : 
                        (N88)? mem[333] : 
                        (N90)? mem[382] : 
                        (N92)? mem[431] : 
                        (N94)? mem[480] : 
                        (N96)? mem[529] : 
                        (N98)? mem[578] : 
                        (N100)? mem[627] : 
                        (N102)? mem[676] : 
                        (N104)? mem[725] : 
                        (N106)? mem[774] : 
                        (N108)? mem[823] : 
                        (N110)? mem[872] : 
                        (N112)? mem[921] : 
                        (N114)? mem[970] : 
                        (N116)? mem[1019] : 
                        (N118)? mem[1068] : 
                        (N120)? mem[1117] : 
                        (N122)? mem[1166] : 
                        (N124)? mem[1215] : 
                        (N126)? mem[1264] : 
                        (N128)? mem[1313] : 
                        (N130)? mem[1362] : 
                        (N132)? mem[1411] : 
                        (N134)? mem[1460] : 
                        (N136)? mem[1509] : 
                        (N138)? mem[1558] : 
                        (N77)? mem[1607] : 
                        (N79)? mem[1656] : 
                        (N81)? mem[1705] : 
                        (N83)? mem[1754] : 
                        (N85)? mem[1803] : 
                        (N87)? mem[1852] : 
                        (N89)? mem[1901] : 
                        (N91)? mem[1950] : 
                        (N93)? mem[1999] : 
                        (N95)? mem[2048] : 
                        (N97)? mem[2097] : 
                        (N99)? mem[2146] : 
                        (N101)? mem[2195] : 
                        (N103)? mem[2244] : 
                        (N105)? mem[2293] : 
                        (N107)? mem[2342] : 
                        (N109)? mem[2391] : 
                        (N111)? mem[2440] : 
                        (N113)? mem[2489] : 
                        (N115)? mem[2538] : 
                        (N117)? mem[2587] : 
                        (N119)? mem[2636] : 
                        (N121)? mem[2685] : 
                        (N123)? mem[2734] : 
                        (N125)? mem[2783] : 
                        (N127)? mem[2832] : 
                        (N129)? mem[2881] : 
                        (N131)? mem[2930] : 
                        (N133)? mem[2979] : 
                        (N135)? mem[3028] : 
                        (N137)? mem[3077] : 
                        (N139)? mem[3126] : 1'b0;
  assign r_data_o[38] = (N76)? mem[38] : 
                        (N78)? mem[87] : 
                        (N80)? mem[136] : 
                        (N82)? mem[185] : 
                        (N84)? mem[234] : 
                        (N86)? mem[283] : 
                        (N88)? mem[332] : 
                        (N90)? mem[381] : 
                        (N92)? mem[430] : 
                        (N94)? mem[479] : 
                        (N96)? mem[528] : 
                        (N98)? mem[577] : 
                        (N100)? mem[626] : 
                        (N102)? mem[675] : 
                        (N104)? mem[724] : 
                        (N106)? mem[773] : 
                        (N108)? mem[822] : 
                        (N110)? mem[871] : 
                        (N112)? mem[920] : 
                        (N114)? mem[969] : 
                        (N116)? mem[1018] : 
                        (N118)? mem[1067] : 
                        (N120)? mem[1116] : 
                        (N122)? mem[1165] : 
                        (N124)? mem[1214] : 
                        (N126)? mem[1263] : 
                        (N128)? mem[1312] : 
                        (N130)? mem[1361] : 
                        (N132)? mem[1410] : 
                        (N134)? mem[1459] : 
                        (N136)? mem[1508] : 
                        (N138)? mem[1557] : 
                        (N77)? mem[1606] : 
                        (N79)? mem[1655] : 
                        (N81)? mem[1704] : 
                        (N83)? mem[1753] : 
                        (N85)? mem[1802] : 
                        (N87)? mem[1851] : 
                        (N89)? mem[1900] : 
                        (N91)? mem[1949] : 
                        (N93)? mem[1998] : 
                        (N95)? mem[2047] : 
                        (N97)? mem[2096] : 
                        (N99)? mem[2145] : 
                        (N101)? mem[2194] : 
                        (N103)? mem[2243] : 
                        (N105)? mem[2292] : 
                        (N107)? mem[2341] : 
                        (N109)? mem[2390] : 
                        (N111)? mem[2439] : 
                        (N113)? mem[2488] : 
                        (N115)? mem[2537] : 
                        (N117)? mem[2586] : 
                        (N119)? mem[2635] : 
                        (N121)? mem[2684] : 
                        (N123)? mem[2733] : 
                        (N125)? mem[2782] : 
                        (N127)? mem[2831] : 
                        (N129)? mem[2880] : 
                        (N131)? mem[2929] : 
                        (N133)? mem[2978] : 
                        (N135)? mem[3027] : 
                        (N137)? mem[3076] : 
                        (N139)? mem[3125] : 1'b0;
  assign r_data_o[37] = (N76)? mem[37] : 
                        (N78)? mem[86] : 
                        (N80)? mem[135] : 
                        (N82)? mem[184] : 
                        (N84)? mem[233] : 
                        (N86)? mem[282] : 
                        (N88)? mem[331] : 
                        (N90)? mem[380] : 
                        (N92)? mem[429] : 
                        (N94)? mem[478] : 
                        (N96)? mem[527] : 
                        (N98)? mem[576] : 
                        (N100)? mem[625] : 
                        (N102)? mem[674] : 
                        (N104)? mem[723] : 
                        (N106)? mem[772] : 
                        (N108)? mem[821] : 
                        (N110)? mem[870] : 
                        (N112)? mem[919] : 
                        (N114)? mem[968] : 
                        (N116)? mem[1017] : 
                        (N118)? mem[1066] : 
                        (N120)? mem[1115] : 
                        (N122)? mem[1164] : 
                        (N124)? mem[1213] : 
                        (N126)? mem[1262] : 
                        (N128)? mem[1311] : 
                        (N130)? mem[1360] : 
                        (N132)? mem[1409] : 
                        (N134)? mem[1458] : 
                        (N136)? mem[1507] : 
                        (N138)? mem[1556] : 
                        (N77)? mem[1605] : 
                        (N79)? mem[1654] : 
                        (N81)? mem[1703] : 
                        (N83)? mem[1752] : 
                        (N85)? mem[1801] : 
                        (N87)? mem[1850] : 
                        (N89)? mem[1899] : 
                        (N91)? mem[1948] : 
                        (N93)? mem[1997] : 
                        (N95)? mem[2046] : 
                        (N97)? mem[2095] : 
                        (N99)? mem[2144] : 
                        (N101)? mem[2193] : 
                        (N103)? mem[2242] : 
                        (N105)? mem[2291] : 
                        (N107)? mem[2340] : 
                        (N109)? mem[2389] : 
                        (N111)? mem[2438] : 
                        (N113)? mem[2487] : 
                        (N115)? mem[2536] : 
                        (N117)? mem[2585] : 
                        (N119)? mem[2634] : 
                        (N121)? mem[2683] : 
                        (N123)? mem[2732] : 
                        (N125)? mem[2781] : 
                        (N127)? mem[2830] : 
                        (N129)? mem[2879] : 
                        (N131)? mem[2928] : 
                        (N133)? mem[2977] : 
                        (N135)? mem[3026] : 
                        (N137)? mem[3075] : 
                        (N139)? mem[3124] : 1'b0;
  assign r_data_o[36] = (N76)? mem[36] : 
                        (N78)? mem[85] : 
                        (N80)? mem[134] : 
                        (N82)? mem[183] : 
                        (N84)? mem[232] : 
                        (N86)? mem[281] : 
                        (N88)? mem[330] : 
                        (N90)? mem[379] : 
                        (N92)? mem[428] : 
                        (N94)? mem[477] : 
                        (N96)? mem[526] : 
                        (N98)? mem[575] : 
                        (N100)? mem[624] : 
                        (N102)? mem[673] : 
                        (N104)? mem[722] : 
                        (N106)? mem[771] : 
                        (N108)? mem[820] : 
                        (N110)? mem[869] : 
                        (N112)? mem[918] : 
                        (N114)? mem[967] : 
                        (N116)? mem[1016] : 
                        (N118)? mem[1065] : 
                        (N120)? mem[1114] : 
                        (N122)? mem[1163] : 
                        (N124)? mem[1212] : 
                        (N126)? mem[1261] : 
                        (N128)? mem[1310] : 
                        (N130)? mem[1359] : 
                        (N132)? mem[1408] : 
                        (N134)? mem[1457] : 
                        (N136)? mem[1506] : 
                        (N138)? mem[1555] : 
                        (N77)? mem[1604] : 
                        (N79)? mem[1653] : 
                        (N81)? mem[1702] : 
                        (N83)? mem[1751] : 
                        (N85)? mem[1800] : 
                        (N87)? mem[1849] : 
                        (N89)? mem[1898] : 
                        (N91)? mem[1947] : 
                        (N93)? mem[1996] : 
                        (N95)? mem[2045] : 
                        (N97)? mem[2094] : 
                        (N99)? mem[2143] : 
                        (N101)? mem[2192] : 
                        (N103)? mem[2241] : 
                        (N105)? mem[2290] : 
                        (N107)? mem[2339] : 
                        (N109)? mem[2388] : 
                        (N111)? mem[2437] : 
                        (N113)? mem[2486] : 
                        (N115)? mem[2535] : 
                        (N117)? mem[2584] : 
                        (N119)? mem[2633] : 
                        (N121)? mem[2682] : 
                        (N123)? mem[2731] : 
                        (N125)? mem[2780] : 
                        (N127)? mem[2829] : 
                        (N129)? mem[2878] : 
                        (N131)? mem[2927] : 
                        (N133)? mem[2976] : 
                        (N135)? mem[3025] : 
                        (N137)? mem[3074] : 
                        (N139)? mem[3123] : 1'b0;
  assign r_data_o[35] = (N76)? mem[35] : 
                        (N78)? mem[84] : 
                        (N80)? mem[133] : 
                        (N82)? mem[182] : 
                        (N84)? mem[231] : 
                        (N86)? mem[280] : 
                        (N88)? mem[329] : 
                        (N90)? mem[378] : 
                        (N92)? mem[427] : 
                        (N94)? mem[476] : 
                        (N96)? mem[525] : 
                        (N98)? mem[574] : 
                        (N100)? mem[623] : 
                        (N102)? mem[672] : 
                        (N104)? mem[721] : 
                        (N106)? mem[770] : 
                        (N108)? mem[819] : 
                        (N110)? mem[868] : 
                        (N112)? mem[917] : 
                        (N114)? mem[966] : 
                        (N116)? mem[1015] : 
                        (N118)? mem[1064] : 
                        (N120)? mem[1113] : 
                        (N122)? mem[1162] : 
                        (N124)? mem[1211] : 
                        (N126)? mem[1260] : 
                        (N128)? mem[1309] : 
                        (N130)? mem[1358] : 
                        (N132)? mem[1407] : 
                        (N134)? mem[1456] : 
                        (N136)? mem[1505] : 
                        (N138)? mem[1554] : 
                        (N77)? mem[1603] : 
                        (N79)? mem[1652] : 
                        (N81)? mem[1701] : 
                        (N83)? mem[1750] : 
                        (N85)? mem[1799] : 
                        (N87)? mem[1848] : 
                        (N89)? mem[1897] : 
                        (N91)? mem[1946] : 
                        (N93)? mem[1995] : 
                        (N95)? mem[2044] : 
                        (N97)? mem[2093] : 
                        (N99)? mem[2142] : 
                        (N101)? mem[2191] : 
                        (N103)? mem[2240] : 
                        (N105)? mem[2289] : 
                        (N107)? mem[2338] : 
                        (N109)? mem[2387] : 
                        (N111)? mem[2436] : 
                        (N113)? mem[2485] : 
                        (N115)? mem[2534] : 
                        (N117)? mem[2583] : 
                        (N119)? mem[2632] : 
                        (N121)? mem[2681] : 
                        (N123)? mem[2730] : 
                        (N125)? mem[2779] : 
                        (N127)? mem[2828] : 
                        (N129)? mem[2877] : 
                        (N131)? mem[2926] : 
                        (N133)? mem[2975] : 
                        (N135)? mem[3024] : 
                        (N137)? mem[3073] : 
                        (N139)? mem[3122] : 1'b0;
  assign r_data_o[34] = (N76)? mem[34] : 
                        (N78)? mem[83] : 
                        (N80)? mem[132] : 
                        (N82)? mem[181] : 
                        (N84)? mem[230] : 
                        (N86)? mem[279] : 
                        (N88)? mem[328] : 
                        (N90)? mem[377] : 
                        (N92)? mem[426] : 
                        (N94)? mem[475] : 
                        (N96)? mem[524] : 
                        (N98)? mem[573] : 
                        (N100)? mem[622] : 
                        (N102)? mem[671] : 
                        (N104)? mem[720] : 
                        (N106)? mem[769] : 
                        (N108)? mem[818] : 
                        (N110)? mem[867] : 
                        (N112)? mem[916] : 
                        (N114)? mem[965] : 
                        (N116)? mem[1014] : 
                        (N118)? mem[1063] : 
                        (N120)? mem[1112] : 
                        (N122)? mem[1161] : 
                        (N124)? mem[1210] : 
                        (N126)? mem[1259] : 
                        (N128)? mem[1308] : 
                        (N130)? mem[1357] : 
                        (N132)? mem[1406] : 
                        (N134)? mem[1455] : 
                        (N136)? mem[1504] : 
                        (N138)? mem[1553] : 
                        (N77)? mem[1602] : 
                        (N79)? mem[1651] : 
                        (N81)? mem[1700] : 
                        (N83)? mem[1749] : 
                        (N85)? mem[1798] : 
                        (N87)? mem[1847] : 
                        (N89)? mem[1896] : 
                        (N91)? mem[1945] : 
                        (N93)? mem[1994] : 
                        (N95)? mem[2043] : 
                        (N97)? mem[2092] : 
                        (N99)? mem[2141] : 
                        (N101)? mem[2190] : 
                        (N103)? mem[2239] : 
                        (N105)? mem[2288] : 
                        (N107)? mem[2337] : 
                        (N109)? mem[2386] : 
                        (N111)? mem[2435] : 
                        (N113)? mem[2484] : 
                        (N115)? mem[2533] : 
                        (N117)? mem[2582] : 
                        (N119)? mem[2631] : 
                        (N121)? mem[2680] : 
                        (N123)? mem[2729] : 
                        (N125)? mem[2778] : 
                        (N127)? mem[2827] : 
                        (N129)? mem[2876] : 
                        (N131)? mem[2925] : 
                        (N133)? mem[2974] : 
                        (N135)? mem[3023] : 
                        (N137)? mem[3072] : 
                        (N139)? mem[3121] : 1'b0;
  assign r_data_o[33] = (N76)? mem[33] : 
                        (N78)? mem[82] : 
                        (N80)? mem[131] : 
                        (N82)? mem[180] : 
                        (N84)? mem[229] : 
                        (N86)? mem[278] : 
                        (N88)? mem[327] : 
                        (N90)? mem[376] : 
                        (N92)? mem[425] : 
                        (N94)? mem[474] : 
                        (N96)? mem[523] : 
                        (N98)? mem[572] : 
                        (N100)? mem[621] : 
                        (N102)? mem[670] : 
                        (N104)? mem[719] : 
                        (N106)? mem[768] : 
                        (N108)? mem[817] : 
                        (N110)? mem[866] : 
                        (N112)? mem[915] : 
                        (N114)? mem[964] : 
                        (N116)? mem[1013] : 
                        (N118)? mem[1062] : 
                        (N120)? mem[1111] : 
                        (N122)? mem[1160] : 
                        (N124)? mem[1209] : 
                        (N126)? mem[1258] : 
                        (N128)? mem[1307] : 
                        (N130)? mem[1356] : 
                        (N132)? mem[1405] : 
                        (N134)? mem[1454] : 
                        (N136)? mem[1503] : 
                        (N138)? mem[1552] : 
                        (N77)? mem[1601] : 
                        (N79)? mem[1650] : 
                        (N81)? mem[1699] : 
                        (N83)? mem[1748] : 
                        (N85)? mem[1797] : 
                        (N87)? mem[1846] : 
                        (N89)? mem[1895] : 
                        (N91)? mem[1944] : 
                        (N93)? mem[1993] : 
                        (N95)? mem[2042] : 
                        (N97)? mem[2091] : 
                        (N99)? mem[2140] : 
                        (N101)? mem[2189] : 
                        (N103)? mem[2238] : 
                        (N105)? mem[2287] : 
                        (N107)? mem[2336] : 
                        (N109)? mem[2385] : 
                        (N111)? mem[2434] : 
                        (N113)? mem[2483] : 
                        (N115)? mem[2532] : 
                        (N117)? mem[2581] : 
                        (N119)? mem[2630] : 
                        (N121)? mem[2679] : 
                        (N123)? mem[2728] : 
                        (N125)? mem[2777] : 
                        (N127)? mem[2826] : 
                        (N129)? mem[2875] : 
                        (N131)? mem[2924] : 
                        (N133)? mem[2973] : 
                        (N135)? mem[3022] : 
                        (N137)? mem[3071] : 
                        (N139)? mem[3120] : 1'b0;
  assign r_data_o[32] = (N76)? mem[32] : 
                        (N78)? mem[81] : 
                        (N80)? mem[130] : 
                        (N82)? mem[179] : 
                        (N84)? mem[228] : 
                        (N86)? mem[277] : 
                        (N88)? mem[326] : 
                        (N90)? mem[375] : 
                        (N92)? mem[424] : 
                        (N94)? mem[473] : 
                        (N96)? mem[522] : 
                        (N98)? mem[571] : 
                        (N100)? mem[620] : 
                        (N102)? mem[669] : 
                        (N104)? mem[718] : 
                        (N106)? mem[767] : 
                        (N108)? mem[816] : 
                        (N110)? mem[865] : 
                        (N112)? mem[914] : 
                        (N114)? mem[963] : 
                        (N116)? mem[1012] : 
                        (N118)? mem[1061] : 
                        (N120)? mem[1110] : 
                        (N122)? mem[1159] : 
                        (N124)? mem[1208] : 
                        (N126)? mem[1257] : 
                        (N128)? mem[1306] : 
                        (N130)? mem[1355] : 
                        (N132)? mem[1404] : 
                        (N134)? mem[1453] : 
                        (N136)? mem[1502] : 
                        (N138)? mem[1551] : 
                        (N77)? mem[1600] : 
                        (N79)? mem[1649] : 
                        (N81)? mem[1698] : 
                        (N83)? mem[1747] : 
                        (N85)? mem[1796] : 
                        (N87)? mem[1845] : 
                        (N89)? mem[1894] : 
                        (N91)? mem[1943] : 
                        (N93)? mem[1992] : 
                        (N95)? mem[2041] : 
                        (N97)? mem[2090] : 
                        (N99)? mem[2139] : 
                        (N101)? mem[2188] : 
                        (N103)? mem[2237] : 
                        (N105)? mem[2286] : 
                        (N107)? mem[2335] : 
                        (N109)? mem[2384] : 
                        (N111)? mem[2433] : 
                        (N113)? mem[2482] : 
                        (N115)? mem[2531] : 
                        (N117)? mem[2580] : 
                        (N119)? mem[2629] : 
                        (N121)? mem[2678] : 
                        (N123)? mem[2727] : 
                        (N125)? mem[2776] : 
                        (N127)? mem[2825] : 
                        (N129)? mem[2874] : 
                        (N131)? mem[2923] : 
                        (N133)? mem[2972] : 
                        (N135)? mem[3021] : 
                        (N137)? mem[3070] : 
                        (N139)? mem[3119] : 1'b0;
  assign r_data_o[31] = (N76)? mem[31] : 
                        (N78)? mem[80] : 
                        (N80)? mem[129] : 
                        (N82)? mem[178] : 
                        (N84)? mem[227] : 
                        (N86)? mem[276] : 
                        (N88)? mem[325] : 
                        (N90)? mem[374] : 
                        (N92)? mem[423] : 
                        (N94)? mem[472] : 
                        (N96)? mem[521] : 
                        (N98)? mem[570] : 
                        (N100)? mem[619] : 
                        (N102)? mem[668] : 
                        (N104)? mem[717] : 
                        (N106)? mem[766] : 
                        (N108)? mem[815] : 
                        (N110)? mem[864] : 
                        (N112)? mem[913] : 
                        (N114)? mem[962] : 
                        (N116)? mem[1011] : 
                        (N118)? mem[1060] : 
                        (N120)? mem[1109] : 
                        (N122)? mem[1158] : 
                        (N124)? mem[1207] : 
                        (N126)? mem[1256] : 
                        (N128)? mem[1305] : 
                        (N130)? mem[1354] : 
                        (N132)? mem[1403] : 
                        (N134)? mem[1452] : 
                        (N136)? mem[1501] : 
                        (N138)? mem[1550] : 
                        (N77)? mem[1599] : 
                        (N79)? mem[1648] : 
                        (N81)? mem[1697] : 
                        (N83)? mem[1746] : 
                        (N85)? mem[1795] : 
                        (N87)? mem[1844] : 
                        (N89)? mem[1893] : 
                        (N91)? mem[1942] : 
                        (N93)? mem[1991] : 
                        (N95)? mem[2040] : 
                        (N97)? mem[2089] : 
                        (N99)? mem[2138] : 
                        (N101)? mem[2187] : 
                        (N103)? mem[2236] : 
                        (N105)? mem[2285] : 
                        (N107)? mem[2334] : 
                        (N109)? mem[2383] : 
                        (N111)? mem[2432] : 
                        (N113)? mem[2481] : 
                        (N115)? mem[2530] : 
                        (N117)? mem[2579] : 
                        (N119)? mem[2628] : 
                        (N121)? mem[2677] : 
                        (N123)? mem[2726] : 
                        (N125)? mem[2775] : 
                        (N127)? mem[2824] : 
                        (N129)? mem[2873] : 
                        (N131)? mem[2922] : 
                        (N133)? mem[2971] : 
                        (N135)? mem[3020] : 
                        (N137)? mem[3069] : 
                        (N139)? mem[3118] : 1'b0;
  assign r_data_o[30] = (N76)? mem[30] : 
                        (N78)? mem[79] : 
                        (N80)? mem[128] : 
                        (N82)? mem[177] : 
                        (N84)? mem[226] : 
                        (N86)? mem[275] : 
                        (N88)? mem[324] : 
                        (N90)? mem[373] : 
                        (N92)? mem[422] : 
                        (N94)? mem[471] : 
                        (N96)? mem[520] : 
                        (N98)? mem[569] : 
                        (N100)? mem[618] : 
                        (N102)? mem[667] : 
                        (N104)? mem[716] : 
                        (N106)? mem[765] : 
                        (N108)? mem[814] : 
                        (N110)? mem[863] : 
                        (N112)? mem[912] : 
                        (N114)? mem[961] : 
                        (N116)? mem[1010] : 
                        (N118)? mem[1059] : 
                        (N120)? mem[1108] : 
                        (N122)? mem[1157] : 
                        (N124)? mem[1206] : 
                        (N126)? mem[1255] : 
                        (N128)? mem[1304] : 
                        (N130)? mem[1353] : 
                        (N132)? mem[1402] : 
                        (N134)? mem[1451] : 
                        (N136)? mem[1500] : 
                        (N138)? mem[1549] : 
                        (N77)? mem[1598] : 
                        (N79)? mem[1647] : 
                        (N81)? mem[1696] : 
                        (N83)? mem[1745] : 
                        (N85)? mem[1794] : 
                        (N87)? mem[1843] : 
                        (N89)? mem[1892] : 
                        (N91)? mem[1941] : 
                        (N93)? mem[1990] : 
                        (N95)? mem[2039] : 
                        (N97)? mem[2088] : 
                        (N99)? mem[2137] : 
                        (N101)? mem[2186] : 
                        (N103)? mem[2235] : 
                        (N105)? mem[2284] : 
                        (N107)? mem[2333] : 
                        (N109)? mem[2382] : 
                        (N111)? mem[2431] : 
                        (N113)? mem[2480] : 
                        (N115)? mem[2529] : 
                        (N117)? mem[2578] : 
                        (N119)? mem[2627] : 
                        (N121)? mem[2676] : 
                        (N123)? mem[2725] : 
                        (N125)? mem[2774] : 
                        (N127)? mem[2823] : 
                        (N129)? mem[2872] : 
                        (N131)? mem[2921] : 
                        (N133)? mem[2970] : 
                        (N135)? mem[3019] : 
                        (N137)? mem[3068] : 
                        (N139)? mem[3117] : 1'b0;
  assign r_data_o[29] = (N76)? mem[29] : 
                        (N78)? mem[78] : 
                        (N80)? mem[127] : 
                        (N82)? mem[176] : 
                        (N84)? mem[225] : 
                        (N86)? mem[274] : 
                        (N88)? mem[323] : 
                        (N90)? mem[372] : 
                        (N92)? mem[421] : 
                        (N94)? mem[470] : 
                        (N96)? mem[519] : 
                        (N98)? mem[568] : 
                        (N100)? mem[617] : 
                        (N102)? mem[666] : 
                        (N104)? mem[715] : 
                        (N106)? mem[764] : 
                        (N108)? mem[813] : 
                        (N110)? mem[862] : 
                        (N112)? mem[911] : 
                        (N114)? mem[960] : 
                        (N116)? mem[1009] : 
                        (N118)? mem[1058] : 
                        (N120)? mem[1107] : 
                        (N122)? mem[1156] : 
                        (N124)? mem[1205] : 
                        (N126)? mem[1254] : 
                        (N128)? mem[1303] : 
                        (N130)? mem[1352] : 
                        (N132)? mem[1401] : 
                        (N134)? mem[1450] : 
                        (N136)? mem[1499] : 
                        (N138)? mem[1548] : 
                        (N77)? mem[1597] : 
                        (N79)? mem[1646] : 
                        (N81)? mem[1695] : 
                        (N83)? mem[1744] : 
                        (N85)? mem[1793] : 
                        (N87)? mem[1842] : 
                        (N89)? mem[1891] : 
                        (N91)? mem[1940] : 
                        (N93)? mem[1989] : 
                        (N95)? mem[2038] : 
                        (N97)? mem[2087] : 
                        (N99)? mem[2136] : 
                        (N101)? mem[2185] : 
                        (N103)? mem[2234] : 
                        (N105)? mem[2283] : 
                        (N107)? mem[2332] : 
                        (N109)? mem[2381] : 
                        (N111)? mem[2430] : 
                        (N113)? mem[2479] : 
                        (N115)? mem[2528] : 
                        (N117)? mem[2577] : 
                        (N119)? mem[2626] : 
                        (N121)? mem[2675] : 
                        (N123)? mem[2724] : 
                        (N125)? mem[2773] : 
                        (N127)? mem[2822] : 
                        (N129)? mem[2871] : 
                        (N131)? mem[2920] : 
                        (N133)? mem[2969] : 
                        (N135)? mem[3018] : 
                        (N137)? mem[3067] : 
                        (N139)? mem[3116] : 1'b0;
  assign r_data_o[28] = (N76)? mem[28] : 
                        (N78)? mem[77] : 
                        (N80)? mem[126] : 
                        (N82)? mem[175] : 
                        (N84)? mem[224] : 
                        (N86)? mem[273] : 
                        (N88)? mem[322] : 
                        (N90)? mem[371] : 
                        (N92)? mem[420] : 
                        (N94)? mem[469] : 
                        (N96)? mem[518] : 
                        (N98)? mem[567] : 
                        (N100)? mem[616] : 
                        (N102)? mem[665] : 
                        (N104)? mem[714] : 
                        (N106)? mem[763] : 
                        (N108)? mem[812] : 
                        (N110)? mem[861] : 
                        (N112)? mem[910] : 
                        (N114)? mem[959] : 
                        (N116)? mem[1008] : 
                        (N118)? mem[1057] : 
                        (N120)? mem[1106] : 
                        (N122)? mem[1155] : 
                        (N124)? mem[1204] : 
                        (N126)? mem[1253] : 
                        (N128)? mem[1302] : 
                        (N130)? mem[1351] : 
                        (N132)? mem[1400] : 
                        (N134)? mem[1449] : 
                        (N136)? mem[1498] : 
                        (N138)? mem[1547] : 
                        (N77)? mem[1596] : 
                        (N79)? mem[1645] : 
                        (N81)? mem[1694] : 
                        (N83)? mem[1743] : 
                        (N85)? mem[1792] : 
                        (N87)? mem[1841] : 
                        (N89)? mem[1890] : 
                        (N91)? mem[1939] : 
                        (N93)? mem[1988] : 
                        (N95)? mem[2037] : 
                        (N97)? mem[2086] : 
                        (N99)? mem[2135] : 
                        (N101)? mem[2184] : 
                        (N103)? mem[2233] : 
                        (N105)? mem[2282] : 
                        (N107)? mem[2331] : 
                        (N109)? mem[2380] : 
                        (N111)? mem[2429] : 
                        (N113)? mem[2478] : 
                        (N115)? mem[2527] : 
                        (N117)? mem[2576] : 
                        (N119)? mem[2625] : 
                        (N121)? mem[2674] : 
                        (N123)? mem[2723] : 
                        (N125)? mem[2772] : 
                        (N127)? mem[2821] : 
                        (N129)? mem[2870] : 
                        (N131)? mem[2919] : 
                        (N133)? mem[2968] : 
                        (N135)? mem[3017] : 
                        (N137)? mem[3066] : 
                        (N139)? mem[3115] : 1'b0;
  assign r_data_o[27] = (N76)? mem[27] : 
                        (N78)? mem[76] : 
                        (N80)? mem[125] : 
                        (N82)? mem[174] : 
                        (N84)? mem[223] : 
                        (N86)? mem[272] : 
                        (N88)? mem[321] : 
                        (N90)? mem[370] : 
                        (N92)? mem[419] : 
                        (N94)? mem[468] : 
                        (N96)? mem[517] : 
                        (N98)? mem[566] : 
                        (N100)? mem[615] : 
                        (N102)? mem[664] : 
                        (N104)? mem[713] : 
                        (N106)? mem[762] : 
                        (N108)? mem[811] : 
                        (N110)? mem[860] : 
                        (N112)? mem[909] : 
                        (N114)? mem[958] : 
                        (N116)? mem[1007] : 
                        (N118)? mem[1056] : 
                        (N120)? mem[1105] : 
                        (N122)? mem[1154] : 
                        (N124)? mem[1203] : 
                        (N126)? mem[1252] : 
                        (N128)? mem[1301] : 
                        (N130)? mem[1350] : 
                        (N132)? mem[1399] : 
                        (N134)? mem[1448] : 
                        (N136)? mem[1497] : 
                        (N138)? mem[1546] : 
                        (N77)? mem[1595] : 
                        (N79)? mem[1644] : 
                        (N81)? mem[1693] : 
                        (N83)? mem[1742] : 
                        (N85)? mem[1791] : 
                        (N87)? mem[1840] : 
                        (N89)? mem[1889] : 
                        (N91)? mem[1938] : 
                        (N93)? mem[1987] : 
                        (N95)? mem[2036] : 
                        (N97)? mem[2085] : 
                        (N99)? mem[2134] : 
                        (N101)? mem[2183] : 
                        (N103)? mem[2232] : 
                        (N105)? mem[2281] : 
                        (N107)? mem[2330] : 
                        (N109)? mem[2379] : 
                        (N111)? mem[2428] : 
                        (N113)? mem[2477] : 
                        (N115)? mem[2526] : 
                        (N117)? mem[2575] : 
                        (N119)? mem[2624] : 
                        (N121)? mem[2673] : 
                        (N123)? mem[2722] : 
                        (N125)? mem[2771] : 
                        (N127)? mem[2820] : 
                        (N129)? mem[2869] : 
                        (N131)? mem[2918] : 
                        (N133)? mem[2967] : 
                        (N135)? mem[3016] : 
                        (N137)? mem[3065] : 
                        (N139)? mem[3114] : 1'b0;
  assign r_data_o[26] = (N76)? mem[26] : 
                        (N78)? mem[75] : 
                        (N80)? mem[124] : 
                        (N82)? mem[173] : 
                        (N84)? mem[222] : 
                        (N86)? mem[271] : 
                        (N88)? mem[320] : 
                        (N90)? mem[369] : 
                        (N92)? mem[418] : 
                        (N94)? mem[467] : 
                        (N96)? mem[516] : 
                        (N98)? mem[565] : 
                        (N100)? mem[614] : 
                        (N102)? mem[663] : 
                        (N104)? mem[712] : 
                        (N106)? mem[761] : 
                        (N108)? mem[810] : 
                        (N110)? mem[859] : 
                        (N112)? mem[908] : 
                        (N114)? mem[957] : 
                        (N116)? mem[1006] : 
                        (N118)? mem[1055] : 
                        (N120)? mem[1104] : 
                        (N122)? mem[1153] : 
                        (N124)? mem[1202] : 
                        (N126)? mem[1251] : 
                        (N128)? mem[1300] : 
                        (N130)? mem[1349] : 
                        (N132)? mem[1398] : 
                        (N134)? mem[1447] : 
                        (N136)? mem[1496] : 
                        (N138)? mem[1545] : 
                        (N77)? mem[1594] : 
                        (N79)? mem[1643] : 
                        (N81)? mem[1692] : 
                        (N83)? mem[1741] : 
                        (N85)? mem[1790] : 
                        (N87)? mem[1839] : 
                        (N89)? mem[1888] : 
                        (N91)? mem[1937] : 
                        (N93)? mem[1986] : 
                        (N95)? mem[2035] : 
                        (N97)? mem[2084] : 
                        (N99)? mem[2133] : 
                        (N101)? mem[2182] : 
                        (N103)? mem[2231] : 
                        (N105)? mem[2280] : 
                        (N107)? mem[2329] : 
                        (N109)? mem[2378] : 
                        (N111)? mem[2427] : 
                        (N113)? mem[2476] : 
                        (N115)? mem[2525] : 
                        (N117)? mem[2574] : 
                        (N119)? mem[2623] : 
                        (N121)? mem[2672] : 
                        (N123)? mem[2721] : 
                        (N125)? mem[2770] : 
                        (N127)? mem[2819] : 
                        (N129)? mem[2868] : 
                        (N131)? mem[2917] : 
                        (N133)? mem[2966] : 
                        (N135)? mem[3015] : 
                        (N137)? mem[3064] : 
                        (N139)? mem[3113] : 1'b0;
  assign r_data_o[25] = (N76)? mem[25] : 
                        (N78)? mem[74] : 
                        (N80)? mem[123] : 
                        (N82)? mem[172] : 
                        (N84)? mem[221] : 
                        (N86)? mem[270] : 
                        (N88)? mem[319] : 
                        (N90)? mem[368] : 
                        (N92)? mem[417] : 
                        (N94)? mem[466] : 
                        (N96)? mem[515] : 
                        (N98)? mem[564] : 
                        (N100)? mem[613] : 
                        (N102)? mem[662] : 
                        (N104)? mem[711] : 
                        (N106)? mem[760] : 
                        (N108)? mem[809] : 
                        (N110)? mem[858] : 
                        (N112)? mem[907] : 
                        (N114)? mem[956] : 
                        (N116)? mem[1005] : 
                        (N118)? mem[1054] : 
                        (N120)? mem[1103] : 
                        (N122)? mem[1152] : 
                        (N124)? mem[1201] : 
                        (N126)? mem[1250] : 
                        (N128)? mem[1299] : 
                        (N130)? mem[1348] : 
                        (N132)? mem[1397] : 
                        (N134)? mem[1446] : 
                        (N136)? mem[1495] : 
                        (N138)? mem[1544] : 
                        (N77)? mem[1593] : 
                        (N79)? mem[1642] : 
                        (N81)? mem[1691] : 
                        (N83)? mem[1740] : 
                        (N85)? mem[1789] : 
                        (N87)? mem[1838] : 
                        (N89)? mem[1887] : 
                        (N91)? mem[1936] : 
                        (N93)? mem[1985] : 
                        (N95)? mem[2034] : 
                        (N97)? mem[2083] : 
                        (N99)? mem[2132] : 
                        (N101)? mem[2181] : 
                        (N103)? mem[2230] : 
                        (N105)? mem[2279] : 
                        (N107)? mem[2328] : 
                        (N109)? mem[2377] : 
                        (N111)? mem[2426] : 
                        (N113)? mem[2475] : 
                        (N115)? mem[2524] : 
                        (N117)? mem[2573] : 
                        (N119)? mem[2622] : 
                        (N121)? mem[2671] : 
                        (N123)? mem[2720] : 
                        (N125)? mem[2769] : 
                        (N127)? mem[2818] : 
                        (N129)? mem[2867] : 
                        (N131)? mem[2916] : 
                        (N133)? mem[2965] : 
                        (N135)? mem[3014] : 
                        (N137)? mem[3063] : 
                        (N139)? mem[3112] : 1'b0;
  assign r_data_o[24] = (N76)? mem[24] : 
                        (N78)? mem[73] : 
                        (N80)? mem[122] : 
                        (N82)? mem[171] : 
                        (N84)? mem[220] : 
                        (N86)? mem[269] : 
                        (N88)? mem[318] : 
                        (N90)? mem[367] : 
                        (N92)? mem[416] : 
                        (N94)? mem[465] : 
                        (N96)? mem[514] : 
                        (N98)? mem[563] : 
                        (N100)? mem[612] : 
                        (N102)? mem[661] : 
                        (N104)? mem[710] : 
                        (N106)? mem[759] : 
                        (N108)? mem[808] : 
                        (N110)? mem[857] : 
                        (N112)? mem[906] : 
                        (N114)? mem[955] : 
                        (N116)? mem[1004] : 
                        (N118)? mem[1053] : 
                        (N120)? mem[1102] : 
                        (N122)? mem[1151] : 
                        (N124)? mem[1200] : 
                        (N126)? mem[1249] : 
                        (N128)? mem[1298] : 
                        (N130)? mem[1347] : 
                        (N132)? mem[1396] : 
                        (N134)? mem[1445] : 
                        (N136)? mem[1494] : 
                        (N138)? mem[1543] : 
                        (N77)? mem[1592] : 
                        (N79)? mem[1641] : 
                        (N81)? mem[1690] : 
                        (N83)? mem[1739] : 
                        (N85)? mem[1788] : 
                        (N87)? mem[1837] : 
                        (N89)? mem[1886] : 
                        (N91)? mem[1935] : 
                        (N93)? mem[1984] : 
                        (N95)? mem[2033] : 
                        (N97)? mem[2082] : 
                        (N99)? mem[2131] : 
                        (N101)? mem[2180] : 
                        (N103)? mem[2229] : 
                        (N105)? mem[2278] : 
                        (N107)? mem[2327] : 
                        (N109)? mem[2376] : 
                        (N111)? mem[2425] : 
                        (N113)? mem[2474] : 
                        (N115)? mem[2523] : 
                        (N117)? mem[2572] : 
                        (N119)? mem[2621] : 
                        (N121)? mem[2670] : 
                        (N123)? mem[2719] : 
                        (N125)? mem[2768] : 
                        (N127)? mem[2817] : 
                        (N129)? mem[2866] : 
                        (N131)? mem[2915] : 
                        (N133)? mem[2964] : 
                        (N135)? mem[3013] : 
                        (N137)? mem[3062] : 
                        (N139)? mem[3111] : 1'b0;
  assign r_data_o[23] = (N76)? mem[23] : 
                        (N78)? mem[72] : 
                        (N80)? mem[121] : 
                        (N82)? mem[170] : 
                        (N84)? mem[219] : 
                        (N86)? mem[268] : 
                        (N88)? mem[317] : 
                        (N90)? mem[366] : 
                        (N92)? mem[415] : 
                        (N94)? mem[464] : 
                        (N96)? mem[513] : 
                        (N98)? mem[562] : 
                        (N100)? mem[611] : 
                        (N102)? mem[660] : 
                        (N104)? mem[709] : 
                        (N106)? mem[758] : 
                        (N108)? mem[807] : 
                        (N110)? mem[856] : 
                        (N112)? mem[905] : 
                        (N114)? mem[954] : 
                        (N116)? mem[1003] : 
                        (N118)? mem[1052] : 
                        (N120)? mem[1101] : 
                        (N122)? mem[1150] : 
                        (N124)? mem[1199] : 
                        (N126)? mem[1248] : 
                        (N128)? mem[1297] : 
                        (N130)? mem[1346] : 
                        (N132)? mem[1395] : 
                        (N134)? mem[1444] : 
                        (N136)? mem[1493] : 
                        (N138)? mem[1542] : 
                        (N77)? mem[1591] : 
                        (N79)? mem[1640] : 
                        (N81)? mem[1689] : 
                        (N83)? mem[1738] : 
                        (N85)? mem[1787] : 
                        (N87)? mem[1836] : 
                        (N89)? mem[1885] : 
                        (N91)? mem[1934] : 
                        (N93)? mem[1983] : 
                        (N95)? mem[2032] : 
                        (N97)? mem[2081] : 
                        (N99)? mem[2130] : 
                        (N101)? mem[2179] : 
                        (N103)? mem[2228] : 
                        (N105)? mem[2277] : 
                        (N107)? mem[2326] : 
                        (N109)? mem[2375] : 
                        (N111)? mem[2424] : 
                        (N113)? mem[2473] : 
                        (N115)? mem[2522] : 
                        (N117)? mem[2571] : 
                        (N119)? mem[2620] : 
                        (N121)? mem[2669] : 
                        (N123)? mem[2718] : 
                        (N125)? mem[2767] : 
                        (N127)? mem[2816] : 
                        (N129)? mem[2865] : 
                        (N131)? mem[2914] : 
                        (N133)? mem[2963] : 
                        (N135)? mem[3012] : 
                        (N137)? mem[3061] : 
                        (N139)? mem[3110] : 1'b0;
  assign r_data_o[22] = (N76)? mem[22] : 
                        (N78)? mem[71] : 
                        (N80)? mem[120] : 
                        (N82)? mem[169] : 
                        (N84)? mem[218] : 
                        (N86)? mem[267] : 
                        (N88)? mem[316] : 
                        (N90)? mem[365] : 
                        (N92)? mem[414] : 
                        (N94)? mem[463] : 
                        (N96)? mem[512] : 
                        (N98)? mem[561] : 
                        (N100)? mem[610] : 
                        (N102)? mem[659] : 
                        (N104)? mem[708] : 
                        (N106)? mem[757] : 
                        (N108)? mem[806] : 
                        (N110)? mem[855] : 
                        (N112)? mem[904] : 
                        (N114)? mem[953] : 
                        (N116)? mem[1002] : 
                        (N118)? mem[1051] : 
                        (N120)? mem[1100] : 
                        (N122)? mem[1149] : 
                        (N124)? mem[1198] : 
                        (N126)? mem[1247] : 
                        (N128)? mem[1296] : 
                        (N130)? mem[1345] : 
                        (N132)? mem[1394] : 
                        (N134)? mem[1443] : 
                        (N136)? mem[1492] : 
                        (N138)? mem[1541] : 
                        (N77)? mem[1590] : 
                        (N79)? mem[1639] : 
                        (N81)? mem[1688] : 
                        (N83)? mem[1737] : 
                        (N85)? mem[1786] : 
                        (N87)? mem[1835] : 
                        (N89)? mem[1884] : 
                        (N91)? mem[1933] : 
                        (N93)? mem[1982] : 
                        (N95)? mem[2031] : 
                        (N97)? mem[2080] : 
                        (N99)? mem[2129] : 
                        (N101)? mem[2178] : 
                        (N103)? mem[2227] : 
                        (N105)? mem[2276] : 
                        (N107)? mem[2325] : 
                        (N109)? mem[2374] : 
                        (N111)? mem[2423] : 
                        (N113)? mem[2472] : 
                        (N115)? mem[2521] : 
                        (N117)? mem[2570] : 
                        (N119)? mem[2619] : 
                        (N121)? mem[2668] : 
                        (N123)? mem[2717] : 
                        (N125)? mem[2766] : 
                        (N127)? mem[2815] : 
                        (N129)? mem[2864] : 
                        (N131)? mem[2913] : 
                        (N133)? mem[2962] : 
                        (N135)? mem[3011] : 
                        (N137)? mem[3060] : 
                        (N139)? mem[3109] : 1'b0;
  assign r_data_o[21] = (N76)? mem[21] : 
                        (N78)? mem[70] : 
                        (N80)? mem[119] : 
                        (N82)? mem[168] : 
                        (N84)? mem[217] : 
                        (N86)? mem[266] : 
                        (N88)? mem[315] : 
                        (N90)? mem[364] : 
                        (N92)? mem[413] : 
                        (N94)? mem[462] : 
                        (N96)? mem[511] : 
                        (N98)? mem[560] : 
                        (N100)? mem[609] : 
                        (N102)? mem[658] : 
                        (N104)? mem[707] : 
                        (N106)? mem[756] : 
                        (N108)? mem[805] : 
                        (N110)? mem[854] : 
                        (N112)? mem[903] : 
                        (N114)? mem[952] : 
                        (N116)? mem[1001] : 
                        (N118)? mem[1050] : 
                        (N120)? mem[1099] : 
                        (N122)? mem[1148] : 
                        (N124)? mem[1197] : 
                        (N126)? mem[1246] : 
                        (N128)? mem[1295] : 
                        (N130)? mem[1344] : 
                        (N132)? mem[1393] : 
                        (N134)? mem[1442] : 
                        (N136)? mem[1491] : 
                        (N138)? mem[1540] : 
                        (N77)? mem[1589] : 
                        (N79)? mem[1638] : 
                        (N81)? mem[1687] : 
                        (N83)? mem[1736] : 
                        (N85)? mem[1785] : 
                        (N87)? mem[1834] : 
                        (N89)? mem[1883] : 
                        (N91)? mem[1932] : 
                        (N93)? mem[1981] : 
                        (N95)? mem[2030] : 
                        (N97)? mem[2079] : 
                        (N99)? mem[2128] : 
                        (N101)? mem[2177] : 
                        (N103)? mem[2226] : 
                        (N105)? mem[2275] : 
                        (N107)? mem[2324] : 
                        (N109)? mem[2373] : 
                        (N111)? mem[2422] : 
                        (N113)? mem[2471] : 
                        (N115)? mem[2520] : 
                        (N117)? mem[2569] : 
                        (N119)? mem[2618] : 
                        (N121)? mem[2667] : 
                        (N123)? mem[2716] : 
                        (N125)? mem[2765] : 
                        (N127)? mem[2814] : 
                        (N129)? mem[2863] : 
                        (N131)? mem[2912] : 
                        (N133)? mem[2961] : 
                        (N135)? mem[3010] : 
                        (N137)? mem[3059] : 
                        (N139)? mem[3108] : 1'b0;
  assign r_data_o[20] = (N76)? mem[20] : 
                        (N78)? mem[69] : 
                        (N80)? mem[118] : 
                        (N82)? mem[167] : 
                        (N84)? mem[216] : 
                        (N86)? mem[265] : 
                        (N88)? mem[314] : 
                        (N90)? mem[363] : 
                        (N92)? mem[412] : 
                        (N94)? mem[461] : 
                        (N96)? mem[510] : 
                        (N98)? mem[559] : 
                        (N100)? mem[608] : 
                        (N102)? mem[657] : 
                        (N104)? mem[706] : 
                        (N106)? mem[755] : 
                        (N108)? mem[804] : 
                        (N110)? mem[853] : 
                        (N112)? mem[902] : 
                        (N114)? mem[951] : 
                        (N116)? mem[1000] : 
                        (N118)? mem[1049] : 
                        (N120)? mem[1098] : 
                        (N122)? mem[1147] : 
                        (N124)? mem[1196] : 
                        (N126)? mem[1245] : 
                        (N128)? mem[1294] : 
                        (N130)? mem[1343] : 
                        (N132)? mem[1392] : 
                        (N134)? mem[1441] : 
                        (N136)? mem[1490] : 
                        (N138)? mem[1539] : 
                        (N77)? mem[1588] : 
                        (N79)? mem[1637] : 
                        (N81)? mem[1686] : 
                        (N83)? mem[1735] : 
                        (N85)? mem[1784] : 
                        (N87)? mem[1833] : 
                        (N89)? mem[1882] : 
                        (N91)? mem[1931] : 
                        (N93)? mem[1980] : 
                        (N95)? mem[2029] : 
                        (N97)? mem[2078] : 
                        (N99)? mem[2127] : 
                        (N101)? mem[2176] : 
                        (N103)? mem[2225] : 
                        (N105)? mem[2274] : 
                        (N107)? mem[2323] : 
                        (N109)? mem[2372] : 
                        (N111)? mem[2421] : 
                        (N113)? mem[2470] : 
                        (N115)? mem[2519] : 
                        (N117)? mem[2568] : 
                        (N119)? mem[2617] : 
                        (N121)? mem[2666] : 
                        (N123)? mem[2715] : 
                        (N125)? mem[2764] : 
                        (N127)? mem[2813] : 
                        (N129)? mem[2862] : 
                        (N131)? mem[2911] : 
                        (N133)? mem[2960] : 
                        (N135)? mem[3009] : 
                        (N137)? mem[3058] : 
                        (N139)? mem[3107] : 1'b0;
  assign r_data_o[19] = (N76)? mem[19] : 
                        (N78)? mem[68] : 
                        (N80)? mem[117] : 
                        (N82)? mem[166] : 
                        (N84)? mem[215] : 
                        (N86)? mem[264] : 
                        (N88)? mem[313] : 
                        (N90)? mem[362] : 
                        (N92)? mem[411] : 
                        (N94)? mem[460] : 
                        (N96)? mem[509] : 
                        (N98)? mem[558] : 
                        (N100)? mem[607] : 
                        (N102)? mem[656] : 
                        (N104)? mem[705] : 
                        (N106)? mem[754] : 
                        (N108)? mem[803] : 
                        (N110)? mem[852] : 
                        (N112)? mem[901] : 
                        (N114)? mem[950] : 
                        (N116)? mem[999] : 
                        (N118)? mem[1048] : 
                        (N120)? mem[1097] : 
                        (N122)? mem[1146] : 
                        (N124)? mem[1195] : 
                        (N126)? mem[1244] : 
                        (N128)? mem[1293] : 
                        (N130)? mem[1342] : 
                        (N132)? mem[1391] : 
                        (N134)? mem[1440] : 
                        (N136)? mem[1489] : 
                        (N138)? mem[1538] : 
                        (N77)? mem[1587] : 
                        (N79)? mem[1636] : 
                        (N81)? mem[1685] : 
                        (N83)? mem[1734] : 
                        (N85)? mem[1783] : 
                        (N87)? mem[1832] : 
                        (N89)? mem[1881] : 
                        (N91)? mem[1930] : 
                        (N93)? mem[1979] : 
                        (N95)? mem[2028] : 
                        (N97)? mem[2077] : 
                        (N99)? mem[2126] : 
                        (N101)? mem[2175] : 
                        (N103)? mem[2224] : 
                        (N105)? mem[2273] : 
                        (N107)? mem[2322] : 
                        (N109)? mem[2371] : 
                        (N111)? mem[2420] : 
                        (N113)? mem[2469] : 
                        (N115)? mem[2518] : 
                        (N117)? mem[2567] : 
                        (N119)? mem[2616] : 
                        (N121)? mem[2665] : 
                        (N123)? mem[2714] : 
                        (N125)? mem[2763] : 
                        (N127)? mem[2812] : 
                        (N129)? mem[2861] : 
                        (N131)? mem[2910] : 
                        (N133)? mem[2959] : 
                        (N135)? mem[3008] : 
                        (N137)? mem[3057] : 
                        (N139)? mem[3106] : 1'b0;
  assign r_data_o[18] = (N76)? mem[18] : 
                        (N78)? mem[67] : 
                        (N80)? mem[116] : 
                        (N82)? mem[165] : 
                        (N84)? mem[214] : 
                        (N86)? mem[263] : 
                        (N88)? mem[312] : 
                        (N90)? mem[361] : 
                        (N92)? mem[410] : 
                        (N94)? mem[459] : 
                        (N96)? mem[508] : 
                        (N98)? mem[557] : 
                        (N100)? mem[606] : 
                        (N102)? mem[655] : 
                        (N104)? mem[704] : 
                        (N106)? mem[753] : 
                        (N108)? mem[802] : 
                        (N110)? mem[851] : 
                        (N112)? mem[900] : 
                        (N114)? mem[949] : 
                        (N116)? mem[998] : 
                        (N118)? mem[1047] : 
                        (N120)? mem[1096] : 
                        (N122)? mem[1145] : 
                        (N124)? mem[1194] : 
                        (N126)? mem[1243] : 
                        (N128)? mem[1292] : 
                        (N130)? mem[1341] : 
                        (N132)? mem[1390] : 
                        (N134)? mem[1439] : 
                        (N136)? mem[1488] : 
                        (N138)? mem[1537] : 
                        (N77)? mem[1586] : 
                        (N79)? mem[1635] : 
                        (N81)? mem[1684] : 
                        (N83)? mem[1733] : 
                        (N85)? mem[1782] : 
                        (N87)? mem[1831] : 
                        (N89)? mem[1880] : 
                        (N91)? mem[1929] : 
                        (N93)? mem[1978] : 
                        (N95)? mem[2027] : 
                        (N97)? mem[2076] : 
                        (N99)? mem[2125] : 
                        (N101)? mem[2174] : 
                        (N103)? mem[2223] : 
                        (N105)? mem[2272] : 
                        (N107)? mem[2321] : 
                        (N109)? mem[2370] : 
                        (N111)? mem[2419] : 
                        (N113)? mem[2468] : 
                        (N115)? mem[2517] : 
                        (N117)? mem[2566] : 
                        (N119)? mem[2615] : 
                        (N121)? mem[2664] : 
                        (N123)? mem[2713] : 
                        (N125)? mem[2762] : 
                        (N127)? mem[2811] : 
                        (N129)? mem[2860] : 
                        (N131)? mem[2909] : 
                        (N133)? mem[2958] : 
                        (N135)? mem[3007] : 
                        (N137)? mem[3056] : 
                        (N139)? mem[3105] : 1'b0;
  assign r_data_o[17] = (N76)? mem[17] : 
                        (N78)? mem[66] : 
                        (N80)? mem[115] : 
                        (N82)? mem[164] : 
                        (N84)? mem[213] : 
                        (N86)? mem[262] : 
                        (N88)? mem[311] : 
                        (N90)? mem[360] : 
                        (N92)? mem[409] : 
                        (N94)? mem[458] : 
                        (N96)? mem[507] : 
                        (N98)? mem[556] : 
                        (N100)? mem[605] : 
                        (N102)? mem[654] : 
                        (N104)? mem[703] : 
                        (N106)? mem[752] : 
                        (N108)? mem[801] : 
                        (N110)? mem[850] : 
                        (N112)? mem[899] : 
                        (N114)? mem[948] : 
                        (N116)? mem[997] : 
                        (N118)? mem[1046] : 
                        (N120)? mem[1095] : 
                        (N122)? mem[1144] : 
                        (N124)? mem[1193] : 
                        (N126)? mem[1242] : 
                        (N128)? mem[1291] : 
                        (N130)? mem[1340] : 
                        (N132)? mem[1389] : 
                        (N134)? mem[1438] : 
                        (N136)? mem[1487] : 
                        (N138)? mem[1536] : 
                        (N77)? mem[1585] : 
                        (N79)? mem[1634] : 
                        (N81)? mem[1683] : 
                        (N83)? mem[1732] : 
                        (N85)? mem[1781] : 
                        (N87)? mem[1830] : 
                        (N89)? mem[1879] : 
                        (N91)? mem[1928] : 
                        (N93)? mem[1977] : 
                        (N95)? mem[2026] : 
                        (N97)? mem[2075] : 
                        (N99)? mem[2124] : 
                        (N101)? mem[2173] : 
                        (N103)? mem[2222] : 
                        (N105)? mem[2271] : 
                        (N107)? mem[2320] : 
                        (N109)? mem[2369] : 
                        (N111)? mem[2418] : 
                        (N113)? mem[2467] : 
                        (N115)? mem[2516] : 
                        (N117)? mem[2565] : 
                        (N119)? mem[2614] : 
                        (N121)? mem[2663] : 
                        (N123)? mem[2712] : 
                        (N125)? mem[2761] : 
                        (N127)? mem[2810] : 
                        (N129)? mem[2859] : 
                        (N131)? mem[2908] : 
                        (N133)? mem[2957] : 
                        (N135)? mem[3006] : 
                        (N137)? mem[3055] : 
                        (N139)? mem[3104] : 1'b0;
  assign r_data_o[16] = (N76)? mem[16] : 
                        (N78)? mem[65] : 
                        (N80)? mem[114] : 
                        (N82)? mem[163] : 
                        (N84)? mem[212] : 
                        (N86)? mem[261] : 
                        (N88)? mem[310] : 
                        (N90)? mem[359] : 
                        (N92)? mem[408] : 
                        (N94)? mem[457] : 
                        (N96)? mem[506] : 
                        (N98)? mem[555] : 
                        (N100)? mem[604] : 
                        (N102)? mem[653] : 
                        (N104)? mem[702] : 
                        (N106)? mem[751] : 
                        (N108)? mem[800] : 
                        (N110)? mem[849] : 
                        (N112)? mem[898] : 
                        (N114)? mem[947] : 
                        (N116)? mem[996] : 
                        (N118)? mem[1045] : 
                        (N120)? mem[1094] : 
                        (N122)? mem[1143] : 
                        (N124)? mem[1192] : 
                        (N126)? mem[1241] : 
                        (N128)? mem[1290] : 
                        (N130)? mem[1339] : 
                        (N132)? mem[1388] : 
                        (N134)? mem[1437] : 
                        (N136)? mem[1486] : 
                        (N138)? mem[1535] : 
                        (N77)? mem[1584] : 
                        (N79)? mem[1633] : 
                        (N81)? mem[1682] : 
                        (N83)? mem[1731] : 
                        (N85)? mem[1780] : 
                        (N87)? mem[1829] : 
                        (N89)? mem[1878] : 
                        (N91)? mem[1927] : 
                        (N93)? mem[1976] : 
                        (N95)? mem[2025] : 
                        (N97)? mem[2074] : 
                        (N99)? mem[2123] : 
                        (N101)? mem[2172] : 
                        (N103)? mem[2221] : 
                        (N105)? mem[2270] : 
                        (N107)? mem[2319] : 
                        (N109)? mem[2368] : 
                        (N111)? mem[2417] : 
                        (N113)? mem[2466] : 
                        (N115)? mem[2515] : 
                        (N117)? mem[2564] : 
                        (N119)? mem[2613] : 
                        (N121)? mem[2662] : 
                        (N123)? mem[2711] : 
                        (N125)? mem[2760] : 
                        (N127)? mem[2809] : 
                        (N129)? mem[2858] : 
                        (N131)? mem[2907] : 
                        (N133)? mem[2956] : 
                        (N135)? mem[3005] : 
                        (N137)? mem[3054] : 
                        (N139)? mem[3103] : 1'b0;
  assign r_data_o[15] = (N76)? mem[15] : 
                        (N78)? mem[64] : 
                        (N80)? mem[113] : 
                        (N82)? mem[162] : 
                        (N84)? mem[211] : 
                        (N86)? mem[260] : 
                        (N88)? mem[309] : 
                        (N90)? mem[358] : 
                        (N92)? mem[407] : 
                        (N94)? mem[456] : 
                        (N96)? mem[505] : 
                        (N98)? mem[554] : 
                        (N100)? mem[603] : 
                        (N102)? mem[652] : 
                        (N104)? mem[701] : 
                        (N106)? mem[750] : 
                        (N108)? mem[799] : 
                        (N110)? mem[848] : 
                        (N112)? mem[897] : 
                        (N114)? mem[946] : 
                        (N116)? mem[995] : 
                        (N118)? mem[1044] : 
                        (N120)? mem[1093] : 
                        (N122)? mem[1142] : 
                        (N124)? mem[1191] : 
                        (N126)? mem[1240] : 
                        (N128)? mem[1289] : 
                        (N130)? mem[1338] : 
                        (N132)? mem[1387] : 
                        (N134)? mem[1436] : 
                        (N136)? mem[1485] : 
                        (N138)? mem[1534] : 
                        (N77)? mem[1583] : 
                        (N79)? mem[1632] : 
                        (N81)? mem[1681] : 
                        (N83)? mem[1730] : 
                        (N85)? mem[1779] : 
                        (N87)? mem[1828] : 
                        (N89)? mem[1877] : 
                        (N91)? mem[1926] : 
                        (N93)? mem[1975] : 
                        (N95)? mem[2024] : 
                        (N97)? mem[2073] : 
                        (N99)? mem[2122] : 
                        (N101)? mem[2171] : 
                        (N103)? mem[2220] : 
                        (N105)? mem[2269] : 
                        (N107)? mem[2318] : 
                        (N109)? mem[2367] : 
                        (N111)? mem[2416] : 
                        (N113)? mem[2465] : 
                        (N115)? mem[2514] : 
                        (N117)? mem[2563] : 
                        (N119)? mem[2612] : 
                        (N121)? mem[2661] : 
                        (N123)? mem[2710] : 
                        (N125)? mem[2759] : 
                        (N127)? mem[2808] : 
                        (N129)? mem[2857] : 
                        (N131)? mem[2906] : 
                        (N133)? mem[2955] : 
                        (N135)? mem[3004] : 
                        (N137)? mem[3053] : 
                        (N139)? mem[3102] : 1'b0;
  assign r_data_o[14] = (N76)? mem[14] : 
                        (N78)? mem[63] : 
                        (N80)? mem[112] : 
                        (N82)? mem[161] : 
                        (N84)? mem[210] : 
                        (N86)? mem[259] : 
                        (N88)? mem[308] : 
                        (N90)? mem[357] : 
                        (N92)? mem[406] : 
                        (N94)? mem[455] : 
                        (N96)? mem[504] : 
                        (N98)? mem[553] : 
                        (N100)? mem[602] : 
                        (N102)? mem[651] : 
                        (N104)? mem[700] : 
                        (N106)? mem[749] : 
                        (N108)? mem[798] : 
                        (N110)? mem[847] : 
                        (N112)? mem[896] : 
                        (N114)? mem[945] : 
                        (N116)? mem[994] : 
                        (N118)? mem[1043] : 
                        (N120)? mem[1092] : 
                        (N122)? mem[1141] : 
                        (N124)? mem[1190] : 
                        (N126)? mem[1239] : 
                        (N128)? mem[1288] : 
                        (N130)? mem[1337] : 
                        (N132)? mem[1386] : 
                        (N134)? mem[1435] : 
                        (N136)? mem[1484] : 
                        (N138)? mem[1533] : 
                        (N77)? mem[1582] : 
                        (N79)? mem[1631] : 
                        (N81)? mem[1680] : 
                        (N83)? mem[1729] : 
                        (N85)? mem[1778] : 
                        (N87)? mem[1827] : 
                        (N89)? mem[1876] : 
                        (N91)? mem[1925] : 
                        (N93)? mem[1974] : 
                        (N95)? mem[2023] : 
                        (N97)? mem[2072] : 
                        (N99)? mem[2121] : 
                        (N101)? mem[2170] : 
                        (N103)? mem[2219] : 
                        (N105)? mem[2268] : 
                        (N107)? mem[2317] : 
                        (N109)? mem[2366] : 
                        (N111)? mem[2415] : 
                        (N113)? mem[2464] : 
                        (N115)? mem[2513] : 
                        (N117)? mem[2562] : 
                        (N119)? mem[2611] : 
                        (N121)? mem[2660] : 
                        (N123)? mem[2709] : 
                        (N125)? mem[2758] : 
                        (N127)? mem[2807] : 
                        (N129)? mem[2856] : 
                        (N131)? mem[2905] : 
                        (N133)? mem[2954] : 
                        (N135)? mem[3003] : 
                        (N137)? mem[3052] : 
                        (N139)? mem[3101] : 1'b0;
  assign r_data_o[13] = (N76)? mem[13] : 
                        (N78)? mem[62] : 
                        (N80)? mem[111] : 
                        (N82)? mem[160] : 
                        (N84)? mem[209] : 
                        (N86)? mem[258] : 
                        (N88)? mem[307] : 
                        (N90)? mem[356] : 
                        (N92)? mem[405] : 
                        (N94)? mem[454] : 
                        (N96)? mem[503] : 
                        (N98)? mem[552] : 
                        (N100)? mem[601] : 
                        (N102)? mem[650] : 
                        (N104)? mem[699] : 
                        (N106)? mem[748] : 
                        (N108)? mem[797] : 
                        (N110)? mem[846] : 
                        (N112)? mem[895] : 
                        (N114)? mem[944] : 
                        (N116)? mem[993] : 
                        (N118)? mem[1042] : 
                        (N120)? mem[1091] : 
                        (N122)? mem[1140] : 
                        (N124)? mem[1189] : 
                        (N126)? mem[1238] : 
                        (N128)? mem[1287] : 
                        (N130)? mem[1336] : 
                        (N132)? mem[1385] : 
                        (N134)? mem[1434] : 
                        (N136)? mem[1483] : 
                        (N138)? mem[1532] : 
                        (N77)? mem[1581] : 
                        (N79)? mem[1630] : 
                        (N81)? mem[1679] : 
                        (N83)? mem[1728] : 
                        (N85)? mem[1777] : 
                        (N87)? mem[1826] : 
                        (N89)? mem[1875] : 
                        (N91)? mem[1924] : 
                        (N93)? mem[1973] : 
                        (N95)? mem[2022] : 
                        (N97)? mem[2071] : 
                        (N99)? mem[2120] : 
                        (N101)? mem[2169] : 
                        (N103)? mem[2218] : 
                        (N105)? mem[2267] : 
                        (N107)? mem[2316] : 
                        (N109)? mem[2365] : 
                        (N111)? mem[2414] : 
                        (N113)? mem[2463] : 
                        (N115)? mem[2512] : 
                        (N117)? mem[2561] : 
                        (N119)? mem[2610] : 
                        (N121)? mem[2659] : 
                        (N123)? mem[2708] : 
                        (N125)? mem[2757] : 
                        (N127)? mem[2806] : 
                        (N129)? mem[2855] : 
                        (N131)? mem[2904] : 
                        (N133)? mem[2953] : 
                        (N135)? mem[3002] : 
                        (N137)? mem[3051] : 
                        (N139)? mem[3100] : 1'b0;
  assign r_data_o[12] = (N76)? mem[12] : 
                        (N78)? mem[61] : 
                        (N80)? mem[110] : 
                        (N82)? mem[159] : 
                        (N84)? mem[208] : 
                        (N86)? mem[257] : 
                        (N88)? mem[306] : 
                        (N90)? mem[355] : 
                        (N92)? mem[404] : 
                        (N94)? mem[453] : 
                        (N96)? mem[502] : 
                        (N98)? mem[551] : 
                        (N100)? mem[600] : 
                        (N102)? mem[649] : 
                        (N104)? mem[698] : 
                        (N106)? mem[747] : 
                        (N108)? mem[796] : 
                        (N110)? mem[845] : 
                        (N112)? mem[894] : 
                        (N114)? mem[943] : 
                        (N116)? mem[992] : 
                        (N118)? mem[1041] : 
                        (N120)? mem[1090] : 
                        (N122)? mem[1139] : 
                        (N124)? mem[1188] : 
                        (N126)? mem[1237] : 
                        (N128)? mem[1286] : 
                        (N130)? mem[1335] : 
                        (N132)? mem[1384] : 
                        (N134)? mem[1433] : 
                        (N136)? mem[1482] : 
                        (N138)? mem[1531] : 
                        (N77)? mem[1580] : 
                        (N79)? mem[1629] : 
                        (N81)? mem[1678] : 
                        (N83)? mem[1727] : 
                        (N85)? mem[1776] : 
                        (N87)? mem[1825] : 
                        (N89)? mem[1874] : 
                        (N91)? mem[1923] : 
                        (N93)? mem[1972] : 
                        (N95)? mem[2021] : 
                        (N97)? mem[2070] : 
                        (N99)? mem[2119] : 
                        (N101)? mem[2168] : 
                        (N103)? mem[2217] : 
                        (N105)? mem[2266] : 
                        (N107)? mem[2315] : 
                        (N109)? mem[2364] : 
                        (N111)? mem[2413] : 
                        (N113)? mem[2462] : 
                        (N115)? mem[2511] : 
                        (N117)? mem[2560] : 
                        (N119)? mem[2609] : 
                        (N121)? mem[2658] : 
                        (N123)? mem[2707] : 
                        (N125)? mem[2756] : 
                        (N127)? mem[2805] : 
                        (N129)? mem[2854] : 
                        (N131)? mem[2903] : 
                        (N133)? mem[2952] : 
                        (N135)? mem[3001] : 
                        (N137)? mem[3050] : 
                        (N139)? mem[3099] : 1'b0;
  assign r_data_o[11] = (N76)? mem[11] : 
                        (N78)? mem[60] : 
                        (N80)? mem[109] : 
                        (N82)? mem[158] : 
                        (N84)? mem[207] : 
                        (N86)? mem[256] : 
                        (N88)? mem[305] : 
                        (N90)? mem[354] : 
                        (N92)? mem[403] : 
                        (N94)? mem[452] : 
                        (N96)? mem[501] : 
                        (N98)? mem[550] : 
                        (N100)? mem[599] : 
                        (N102)? mem[648] : 
                        (N104)? mem[697] : 
                        (N106)? mem[746] : 
                        (N108)? mem[795] : 
                        (N110)? mem[844] : 
                        (N112)? mem[893] : 
                        (N114)? mem[942] : 
                        (N116)? mem[991] : 
                        (N118)? mem[1040] : 
                        (N120)? mem[1089] : 
                        (N122)? mem[1138] : 
                        (N124)? mem[1187] : 
                        (N126)? mem[1236] : 
                        (N128)? mem[1285] : 
                        (N130)? mem[1334] : 
                        (N132)? mem[1383] : 
                        (N134)? mem[1432] : 
                        (N136)? mem[1481] : 
                        (N138)? mem[1530] : 
                        (N77)? mem[1579] : 
                        (N79)? mem[1628] : 
                        (N81)? mem[1677] : 
                        (N83)? mem[1726] : 
                        (N85)? mem[1775] : 
                        (N87)? mem[1824] : 
                        (N89)? mem[1873] : 
                        (N91)? mem[1922] : 
                        (N93)? mem[1971] : 
                        (N95)? mem[2020] : 
                        (N97)? mem[2069] : 
                        (N99)? mem[2118] : 
                        (N101)? mem[2167] : 
                        (N103)? mem[2216] : 
                        (N105)? mem[2265] : 
                        (N107)? mem[2314] : 
                        (N109)? mem[2363] : 
                        (N111)? mem[2412] : 
                        (N113)? mem[2461] : 
                        (N115)? mem[2510] : 
                        (N117)? mem[2559] : 
                        (N119)? mem[2608] : 
                        (N121)? mem[2657] : 
                        (N123)? mem[2706] : 
                        (N125)? mem[2755] : 
                        (N127)? mem[2804] : 
                        (N129)? mem[2853] : 
                        (N131)? mem[2902] : 
                        (N133)? mem[2951] : 
                        (N135)? mem[3000] : 
                        (N137)? mem[3049] : 
                        (N139)? mem[3098] : 1'b0;
  assign r_data_o[10] = (N76)? mem[10] : 
                        (N78)? mem[59] : 
                        (N80)? mem[108] : 
                        (N82)? mem[157] : 
                        (N84)? mem[206] : 
                        (N86)? mem[255] : 
                        (N88)? mem[304] : 
                        (N90)? mem[353] : 
                        (N92)? mem[402] : 
                        (N94)? mem[451] : 
                        (N96)? mem[500] : 
                        (N98)? mem[549] : 
                        (N100)? mem[598] : 
                        (N102)? mem[647] : 
                        (N104)? mem[696] : 
                        (N106)? mem[745] : 
                        (N108)? mem[794] : 
                        (N110)? mem[843] : 
                        (N112)? mem[892] : 
                        (N114)? mem[941] : 
                        (N116)? mem[990] : 
                        (N118)? mem[1039] : 
                        (N120)? mem[1088] : 
                        (N122)? mem[1137] : 
                        (N124)? mem[1186] : 
                        (N126)? mem[1235] : 
                        (N128)? mem[1284] : 
                        (N130)? mem[1333] : 
                        (N132)? mem[1382] : 
                        (N134)? mem[1431] : 
                        (N136)? mem[1480] : 
                        (N138)? mem[1529] : 
                        (N77)? mem[1578] : 
                        (N79)? mem[1627] : 
                        (N81)? mem[1676] : 
                        (N83)? mem[1725] : 
                        (N85)? mem[1774] : 
                        (N87)? mem[1823] : 
                        (N89)? mem[1872] : 
                        (N91)? mem[1921] : 
                        (N93)? mem[1970] : 
                        (N95)? mem[2019] : 
                        (N97)? mem[2068] : 
                        (N99)? mem[2117] : 
                        (N101)? mem[2166] : 
                        (N103)? mem[2215] : 
                        (N105)? mem[2264] : 
                        (N107)? mem[2313] : 
                        (N109)? mem[2362] : 
                        (N111)? mem[2411] : 
                        (N113)? mem[2460] : 
                        (N115)? mem[2509] : 
                        (N117)? mem[2558] : 
                        (N119)? mem[2607] : 
                        (N121)? mem[2656] : 
                        (N123)? mem[2705] : 
                        (N125)? mem[2754] : 
                        (N127)? mem[2803] : 
                        (N129)? mem[2852] : 
                        (N131)? mem[2901] : 
                        (N133)? mem[2950] : 
                        (N135)? mem[2999] : 
                        (N137)? mem[3048] : 
                        (N139)? mem[3097] : 1'b0;
  assign r_data_o[9] = (N76)? mem[9] : 
                       (N78)? mem[58] : 
                       (N80)? mem[107] : 
                       (N82)? mem[156] : 
                       (N84)? mem[205] : 
                       (N86)? mem[254] : 
                       (N88)? mem[303] : 
                       (N90)? mem[352] : 
                       (N92)? mem[401] : 
                       (N94)? mem[450] : 
                       (N96)? mem[499] : 
                       (N98)? mem[548] : 
                       (N100)? mem[597] : 
                       (N102)? mem[646] : 
                       (N104)? mem[695] : 
                       (N106)? mem[744] : 
                       (N108)? mem[793] : 
                       (N110)? mem[842] : 
                       (N112)? mem[891] : 
                       (N114)? mem[940] : 
                       (N116)? mem[989] : 
                       (N118)? mem[1038] : 
                       (N120)? mem[1087] : 
                       (N122)? mem[1136] : 
                       (N124)? mem[1185] : 
                       (N126)? mem[1234] : 
                       (N128)? mem[1283] : 
                       (N130)? mem[1332] : 
                       (N132)? mem[1381] : 
                       (N134)? mem[1430] : 
                       (N136)? mem[1479] : 
                       (N138)? mem[1528] : 
                       (N77)? mem[1577] : 
                       (N79)? mem[1626] : 
                       (N81)? mem[1675] : 
                       (N83)? mem[1724] : 
                       (N85)? mem[1773] : 
                       (N87)? mem[1822] : 
                       (N89)? mem[1871] : 
                       (N91)? mem[1920] : 
                       (N93)? mem[1969] : 
                       (N95)? mem[2018] : 
                       (N97)? mem[2067] : 
                       (N99)? mem[2116] : 
                       (N101)? mem[2165] : 
                       (N103)? mem[2214] : 
                       (N105)? mem[2263] : 
                       (N107)? mem[2312] : 
                       (N109)? mem[2361] : 
                       (N111)? mem[2410] : 
                       (N113)? mem[2459] : 
                       (N115)? mem[2508] : 
                       (N117)? mem[2557] : 
                       (N119)? mem[2606] : 
                       (N121)? mem[2655] : 
                       (N123)? mem[2704] : 
                       (N125)? mem[2753] : 
                       (N127)? mem[2802] : 
                       (N129)? mem[2851] : 
                       (N131)? mem[2900] : 
                       (N133)? mem[2949] : 
                       (N135)? mem[2998] : 
                       (N137)? mem[3047] : 
                       (N139)? mem[3096] : 1'b0;
  assign r_data_o[8] = (N76)? mem[8] : 
                       (N78)? mem[57] : 
                       (N80)? mem[106] : 
                       (N82)? mem[155] : 
                       (N84)? mem[204] : 
                       (N86)? mem[253] : 
                       (N88)? mem[302] : 
                       (N90)? mem[351] : 
                       (N92)? mem[400] : 
                       (N94)? mem[449] : 
                       (N96)? mem[498] : 
                       (N98)? mem[547] : 
                       (N100)? mem[596] : 
                       (N102)? mem[645] : 
                       (N104)? mem[694] : 
                       (N106)? mem[743] : 
                       (N108)? mem[792] : 
                       (N110)? mem[841] : 
                       (N112)? mem[890] : 
                       (N114)? mem[939] : 
                       (N116)? mem[988] : 
                       (N118)? mem[1037] : 
                       (N120)? mem[1086] : 
                       (N122)? mem[1135] : 
                       (N124)? mem[1184] : 
                       (N126)? mem[1233] : 
                       (N128)? mem[1282] : 
                       (N130)? mem[1331] : 
                       (N132)? mem[1380] : 
                       (N134)? mem[1429] : 
                       (N136)? mem[1478] : 
                       (N138)? mem[1527] : 
                       (N77)? mem[1576] : 
                       (N79)? mem[1625] : 
                       (N81)? mem[1674] : 
                       (N83)? mem[1723] : 
                       (N85)? mem[1772] : 
                       (N87)? mem[1821] : 
                       (N89)? mem[1870] : 
                       (N91)? mem[1919] : 
                       (N93)? mem[1968] : 
                       (N95)? mem[2017] : 
                       (N97)? mem[2066] : 
                       (N99)? mem[2115] : 
                       (N101)? mem[2164] : 
                       (N103)? mem[2213] : 
                       (N105)? mem[2262] : 
                       (N107)? mem[2311] : 
                       (N109)? mem[2360] : 
                       (N111)? mem[2409] : 
                       (N113)? mem[2458] : 
                       (N115)? mem[2507] : 
                       (N117)? mem[2556] : 
                       (N119)? mem[2605] : 
                       (N121)? mem[2654] : 
                       (N123)? mem[2703] : 
                       (N125)? mem[2752] : 
                       (N127)? mem[2801] : 
                       (N129)? mem[2850] : 
                       (N131)? mem[2899] : 
                       (N133)? mem[2948] : 
                       (N135)? mem[2997] : 
                       (N137)? mem[3046] : 
                       (N139)? mem[3095] : 1'b0;
  assign r_data_o[7] = (N76)? mem[7] : 
                       (N78)? mem[56] : 
                       (N80)? mem[105] : 
                       (N82)? mem[154] : 
                       (N84)? mem[203] : 
                       (N86)? mem[252] : 
                       (N88)? mem[301] : 
                       (N90)? mem[350] : 
                       (N92)? mem[399] : 
                       (N94)? mem[448] : 
                       (N96)? mem[497] : 
                       (N98)? mem[546] : 
                       (N100)? mem[595] : 
                       (N102)? mem[644] : 
                       (N104)? mem[693] : 
                       (N106)? mem[742] : 
                       (N108)? mem[791] : 
                       (N110)? mem[840] : 
                       (N112)? mem[889] : 
                       (N114)? mem[938] : 
                       (N116)? mem[987] : 
                       (N118)? mem[1036] : 
                       (N120)? mem[1085] : 
                       (N122)? mem[1134] : 
                       (N124)? mem[1183] : 
                       (N126)? mem[1232] : 
                       (N128)? mem[1281] : 
                       (N130)? mem[1330] : 
                       (N132)? mem[1379] : 
                       (N134)? mem[1428] : 
                       (N136)? mem[1477] : 
                       (N138)? mem[1526] : 
                       (N77)? mem[1575] : 
                       (N79)? mem[1624] : 
                       (N81)? mem[1673] : 
                       (N83)? mem[1722] : 
                       (N85)? mem[1771] : 
                       (N87)? mem[1820] : 
                       (N89)? mem[1869] : 
                       (N91)? mem[1918] : 
                       (N93)? mem[1967] : 
                       (N95)? mem[2016] : 
                       (N97)? mem[2065] : 
                       (N99)? mem[2114] : 
                       (N101)? mem[2163] : 
                       (N103)? mem[2212] : 
                       (N105)? mem[2261] : 
                       (N107)? mem[2310] : 
                       (N109)? mem[2359] : 
                       (N111)? mem[2408] : 
                       (N113)? mem[2457] : 
                       (N115)? mem[2506] : 
                       (N117)? mem[2555] : 
                       (N119)? mem[2604] : 
                       (N121)? mem[2653] : 
                       (N123)? mem[2702] : 
                       (N125)? mem[2751] : 
                       (N127)? mem[2800] : 
                       (N129)? mem[2849] : 
                       (N131)? mem[2898] : 
                       (N133)? mem[2947] : 
                       (N135)? mem[2996] : 
                       (N137)? mem[3045] : 
                       (N139)? mem[3094] : 1'b0;
  assign r_data_o[6] = (N76)? mem[6] : 
                       (N78)? mem[55] : 
                       (N80)? mem[104] : 
                       (N82)? mem[153] : 
                       (N84)? mem[202] : 
                       (N86)? mem[251] : 
                       (N88)? mem[300] : 
                       (N90)? mem[349] : 
                       (N92)? mem[398] : 
                       (N94)? mem[447] : 
                       (N96)? mem[496] : 
                       (N98)? mem[545] : 
                       (N100)? mem[594] : 
                       (N102)? mem[643] : 
                       (N104)? mem[692] : 
                       (N106)? mem[741] : 
                       (N108)? mem[790] : 
                       (N110)? mem[839] : 
                       (N112)? mem[888] : 
                       (N114)? mem[937] : 
                       (N116)? mem[986] : 
                       (N118)? mem[1035] : 
                       (N120)? mem[1084] : 
                       (N122)? mem[1133] : 
                       (N124)? mem[1182] : 
                       (N126)? mem[1231] : 
                       (N128)? mem[1280] : 
                       (N130)? mem[1329] : 
                       (N132)? mem[1378] : 
                       (N134)? mem[1427] : 
                       (N136)? mem[1476] : 
                       (N138)? mem[1525] : 
                       (N77)? mem[1574] : 
                       (N79)? mem[1623] : 
                       (N81)? mem[1672] : 
                       (N83)? mem[1721] : 
                       (N85)? mem[1770] : 
                       (N87)? mem[1819] : 
                       (N89)? mem[1868] : 
                       (N91)? mem[1917] : 
                       (N93)? mem[1966] : 
                       (N95)? mem[2015] : 
                       (N97)? mem[2064] : 
                       (N99)? mem[2113] : 
                       (N101)? mem[2162] : 
                       (N103)? mem[2211] : 
                       (N105)? mem[2260] : 
                       (N107)? mem[2309] : 
                       (N109)? mem[2358] : 
                       (N111)? mem[2407] : 
                       (N113)? mem[2456] : 
                       (N115)? mem[2505] : 
                       (N117)? mem[2554] : 
                       (N119)? mem[2603] : 
                       (N121)? mem[2652] : 
                       (N123)? mem[2701] : 
                       (N125)? mem[2750] : 
                       (N127)? mem[2799] : 
                       (N129)? mem[2848] : 
                       (N131)? mem[2897] : 
                       (N133)? mem[2946] : 
                       (N135)? mem[2995] : 
                       (N137)? mem[3044] : 
                       (N139)? mem[3093] : 1'b0;
  assign r_data_o[5] = (N76)? mem[5] : 
                       (N78)? mem[54] : 
                       (N80)? mem[103] : 
                       (N82)? mem[152] : 
                       (N84)? mem[201] : 
                       (N86)? mem[250] : 
                       (N88)? mem[299] : 
                       (N90)? mem[348] : 
                       (N92)? mem[397] : 
                       (N94)? mem[446] : 
                       (N96)? mem[495] : 
                       (N98)? mem[544] : 
                       (N100)? mem[593] : 
                       (N102)? mem[642] : 
                       (N104)? mem[691] : 
                       (N106)? mem[740] : 
                       (N108)? mem[789] : 
                       (N110)? mem[838] : 
                       (N112)? mem[887] : 
                       (N114)? mem[936] : 
                       (N116)? mem[985] : 
                       (N118)? mem[1034] : 
                       (N120)? mem[1083] : 
                       (N122)? mem[1132] : 
                       (N124)? mem[1181] : 
                       (N126)? mem[1230] : 
                       (N128)? mem[1279] : 
                       (N130)? mem[1328] : 
                       (N132)? mem[1377] : 
                       (N134)? mem[1426] : 
                       (N136)? mem[1475] : 
                       (N138)? mem[1524] : 
                       (N77)? mem[1573] : 
                       (N79)? mem[1622] : 
                       (N81)? mem[1671] : 
                       (N83)? mem[1720] : 
                       (N85)? mem[1769] : 
                       (N87)? mem[1818] : 
                       (N89)? mem[1867] : 
                       (N91)? mem[1916] : 
                       (N93)? mem[1965] : 
                       (N95)? mem[2014] : 
                       (N97)? mem[2063] : 
                       (N99)? mem[2112] : 
                       (N101)? mem[2161] : 
                       (N103)? mem[2210] : 
                       (N105)? mem[2259] : 
                       (N107)? mem[2308] : 
                       (N109)? mem[2357] : 
                       (N111)? mem[2406] : 
                       (N113)? mem[2455] : 
                       (N115)? mem[2504] : 
                       (N117)? mem[2553] : 
                       (N119)? mem[2602] : 
                       (N121)? mem[2651] : 
                       (N123)? mem[2700] : 
                       (N125)? mem[2749] : 
                       (N127)? mem[2798] : 
                       (N129)? mem[2847] : 
                       (N131)? mem[2896] : 
                       (N133)? mem[2945] : 
                       (N135)? mem[2994] : 
                       (N137)? mem[3043] : 
                       (N139)? mem[3092] : 1'b0;
  assign r_data_o[4] = (N76)? mem[4] : 
                       (N78)? mem[53] : 
                       (N80)? mem[102] : 
                       (N82)? mem[151] : 
                       (N84)? mem[200] : 
                       (N86)? mem[249] : 
                       (N88)? mem[298] : 
                       (N90)? mem[347] : 
                       (N92)? mem[396] : 
                       (N94)? mem[445] : 
                       (N96)? mem[494] : 
                       (N98)? mem[543] : 
                       (N100)? mem[592] : 
                       (N102)? mem[641] : 
                       (N104)? mem[690] : 
                       (N106)? mem[739] : 
                       (N108)? mem[788] : 
                       (N110)? mem[837] : 
                       (N112)? mem[886] : 
                       (N114)? mem[935] : 
                       (N116)? mem[984] : 
                       (N118)? mem[1033] : 
                       (N120)? mem[1082] : 
                       (N122)? mem[1131] : 
                       (N124)? mem[1180] : 
                       (N126)? mem[1229] : 
                       (N128)? mem[1278] : 
                       (N130)? mem[1327] : 
                       (N132)? mem[1376] : 
                       (N134)? mem[1425] : 
                       (N136)? mem[1474] : 
                       (N138)? mem[1523] : 
                       (N77)? mem[1572] : 
                       (N79)? mem[1621] : 
                       (N81)? mem[1670] : 
                       (N83)? mem[1719] : 
                       (N85)? mem[1768] : 
                       (N87)? mem[1817] : 
                       (N89)? mem[1866] : 
                       (N91)? mem[1915] : 
                       (N93)? mem[1964] : 
                       (N95)? mem[2013] : 
                       (N97)? mem[2062] : 
                       (N99)? mem[2111] : 
                       (N101)? mem[2160] : 
                       (N103)? mem[2209] : 
                       (N105)? mem[2258] : 
                       (N107)? mem[2307] : 
                       (N109)? mem[2356] : 
                       (N111)? mem[2405] : 
                       (N113)? mem[2454] : 
                       (N115)? mem[2503] : 
                       (N117)? mem[2552] : 
                       (N119)? mem[2601] : 
                       (N121)? mem[2650] : 
                       (N123)? mem[2699] : 
                       (N125)? mem[2748] : 
                       (N127)? mem[2797] : 
                       (N129)? mem[2846] : 
                       (N131)? mem[2895] : 
                       (N133)? mem[2944] : 
                       (N135)? mem[2993] : 
                       (N137)? mem[3042] : 
                       (N139)? mem[3091] : 1'b0;
  assign r_data_o[3] = (N76)? mem[3] : 
                       (N78)? mem[52] : 
                       (N80)? mem[101] : 
                       (N82)? mem[150] : 
                       (N84)? mem[199] : 
                       (N86)? mem[248] : 
                       (N88)? mem[297] : 
                       (N90)? mem[346] : 
                       (N92)? mem[395] : 
                       (N94)? mem[444] : 
                       (N96)? mem[493] : 
                       (N98)? mem[542] : 
                       (N100)? mem[591] : 
                       (N102)? mem[640] : 
                       (N104)? mem[689] : 
                       (N106)? mem[738] : 
                       (N108)? mem[787] : 
                       (N110)? mem[836] : 
                       (N112)? mem[885] : 
                       (N114)? mem[934] : 
                       (N116)? mem[983] : 
                       (N118)? mem[1032] : 
                       (N120)? mem[1081] : 
                       (N122)? mem[1130] : 
                       (N124)? mem[1179] : 
                       (N126)? mem[1228] : 
                       (N128)? mem[1277] : 
                       (N130)? mem[1326] : 
                       (N132)? mem[1375] : 
                       (N134)? mem[1424] : 
                       (N136)? mem[1473] : 
                       (N138)? mem[1522] : 
                       (N77)? mem[1571] : 
                       (N79)? mem[1620] : 
                       (N81)? mem[1669] : 
                       (N83)? mem[1718] : 
                       (N85)? mem[1767] : 
                       (N87)? mem[1816] : 
                       (N89)? mem[1865] : 
                       (N91)? mem[1914] : 
                       (N93)? mem[1963] : 
                       (N95)? mem[2012] : 
                       (N97)? mem[2061] : 
                       (N99)? mem[2110] : 
                       (N101)? mem[2159] : 
                       (N103)? mem[2208] : 
                       (N105)? mem[2257] : 
                       (N107)? mem[2306] : 
                       (N109)? mem[2355] : 
                       (N111)? mem[2404] : 
                       (N113)? mem[2453] : 
                       (N115)? mem[2502] : 
                       (N117)? mem[2551] : 
                       (N119)? mem[2600] : 
                       (N121)? mem[2649] : 
                       (N123)? mem[2698] : 
                       (N125)? mem[2747] : 
                       (N127)? mem[2796] : 
                       (N129)? mem[2845] : 
                       (N131)? mem[2894] : 
                       (N133)? mem[2943] : 
                       (N135)? mem[2992] : 
                       (N137)? mem[3041] : 
                       (N139)? mem[3090] : 1'b0;
  assign r_data_o[2] = (N76)? mem[2] : 
                       (N78)? mem[51] : 
                       (N80)? mem[100] : 
                       (N82)? mem[149] : 
                       (N84)? mem[198] : 
                       (N86)? mem[247] : 
                       (N88)? mem[296] : 
                       (N90)? mem[345] : 
                       (N92)? mem[394] : 
                       (N94)? mem[443] : 
                       (N96)? mem[492] : 
                       (N98)? mem[541] : 
                       (N100)? mem[590] : 
                       (N102)? mem[639] : 
                       (N104)? mem[688] : 
                       (N106)? mem[737] : 
                       (N108)? mem[786] : 
                       (N110)? mem[835] : 
                       (N112)? mem[884] : 
                       (N114)? mem[933] : 
                       (N116)? mem[982] : 
                       (N118)? mem[1031] : 
                       (N120)? mem[1080] : 
                       (N122)? mem[1129] : 
                       (N124)? mem[1178] : 
                       (N126)? mem[1227] : 
                       (N128)? mem[1276] : 
                       (N130)? mem[1325] : 
                       (N132)? mem[1374] : 
                       (N134)? mem[1423] : 
                       (N136)? mem[1472] : 
                       (N138)? mem[1521] : 
                       (N77)? mem[1570] : 
                       (N79)? mem[1619] : 
                       (N81)? mem[1668] : 
                       (N83)? mem[1717] : 
                       (N85)? mem[1766] : 
                       (N87)? mem[1815] : 
                       (N89)? mem[1864] : 
                       (N91)? mem[1913] : 
                       (N93)? mem[1962] : 
                       (N95)? mem[2011] : 
                       (N97)? mem[2060] : 
                       (N99)? mem[2109] : 
                       (N101)? mem[2158] : 
                       (N103)? mem[2207] : 
                       (N105)? mem[2256] : 
                       (N107)? mem[2305] : 
                       (N109)? mem[2354] : 
                       (N111)? mem[2403] : 
                       (N113)? mem[2452] : 
                       (N115)? mem[2501] : 
                       (N117)? mem[2550] : 
                       (N119)? mem[2599] : 
                       (N121)? mem[2648] : 
                       (N123)? mem[2697] : 
                       (N125)? mem[2746] : 
                       (N127)? mem[2795] : 
                       (N129)? mem[2844] : 
                       (N131)? mem[2893] : 
                       (N133)? mem[2942] : 
                       (N135)? mem[2991] : 
                       (N137)? mem[3040] : 
                       (N139)? mem[3089] : 1'b0;
  assign r_data_o[1] = (N76)? mem[1] : 
                       (N78)? mem[50] : 
                       (N80)? mem[99] : 
                       (N82)? mem[148] : 
                       (N84)? mem[197] : 
                       (N86)? mem[246] : 
                       (N88)? mem[295] : 
                       (N90)? mem[344] : 
                       (N92)? mem[393] : 
                       (N94)? mem[442] : 
                       (N96)? mem[491] : 
                       (N98)? mem[540] : 
                       (N100)? mem[589] : 
                       (N102)? mem[638] : 
                       (N104)? mem[687] : 
                       (N106)? mem[736] : 
                       (N108)? mem[785] : 
                       (N110)? mem[834] : 
                       (N112)? mem[883] : 
                       (N114)? mem[932] : 
                       (N116)? mem[981] : 
                       (N118)? mem[1030] : 
                       (N120)? mem[1079] : 
                       (N122)? mem[1128] : 
                       (N124)? mem[1177] : 
                       (N126)? mem[1226] : 
                       (N128)? mem[1275] : 
                       (N130)? mem[1324] : 
                       (N132)? mem[1373] : 
                       (N134)? mem[1422] : 
                       (N136)? mem[1471] : 
                       (N138)? mem[1520] : 
                       (N77)? mem[1569] : 
                       (N79)? mem[1618] : 
                       (N81)? mem[1667] : 
                       (N83)? mem[1716] : 
                       (N85)? mem[1765] : 
                       (N87)? mem[1814] : 
                       (N89)? mem[1863] : 
                       (N91)? mem[1912] : 
                       (N93)? mem[1961] : 
                       (N95)? mem[2010] : 
                       (N97)? mem[2059] : 
                       (N99)? mem[2108] : 
                       (N101)? mem[2157] : 
                       (N103)? mem[2206] : 
                       (N105)? mem[2255] : 
                       (N107)? mem[2304] : 
                       (N109)? mem[2353] : 
                       (N111)? mem[2402] : 
                       (N113)? mem[2451] : 
                       (N115)? mem[2500] : 
                       (N117)? mem[2549] : 
                       (N119)? mem[2598] : 
                       (N121)? mem[2647] : 
                       (N123)? mem[2696] : 
                       (N125)? mem[2745] : 
                       (N127)? mem[2794] : 
                       (N129)? mem[2843] : 
                       (N131)? mem[2892] : 
                       (N133)? mem[2941] : 
                       (N135)? mem[2990] : 
                       (N137)? mem[3039] : 
                       (N139)? mem[3088] : 1'b0;
  assign r_data_o[0] = (N76)? mem[0] : 
                       (N78)? mem[49] : 
                       (N80)? mem[98] : 
                       (N82)? mem[147] : 
                       (N84)? mem[196] : 
                       (N86)? mem[245] : 
                       (N88)? mem[294] : 
                       (N90)? mem[343] : 
                       (N92)? mem[392] : 
                       (N94)? mem[441] : 
                       (N96)? mem[490] : 
                       (N98)? mem[539] : 
                       (N100)? mem[588] : 
                       (N102)? mem[637] : 
                       (N104)? mem[686] : 
                       (N106)? mem[735] : 
                       (N108)? mem[784] : 
                       (N110)? mem[833] : 
                       (N112)? mem[882] : 
                       (N114)? mem[931] : 
                       (N116)? mem[980] : 
                       (N118)? mem[1029] : 
                       (N120)? mem[1078] : 
                       (N122)? mem[1127] : 
                       (N124)? mem[1176] : 
                       (N126)? mem[1225] : 
                       (N128)? mem[1274] : 
                       (N130)? mem[1323] : 
                       (N132)? mem[1372] : 
                       (N134)? mem[1421] : 
                       (N136)? mem[1470] : 
                       (N138)? mem[1519] : 
                       (N77)? mem[1568] : 
                       (N79)? mem[1617] : 
                       (N81)? mem[1666] : 
                       (N83)? mem[1715] : 
                       (N85)? mem[1764] : 
                       (N87)? mem[1813] : 
                       (N89)? mem[1862] : 
                       (N91)? mem[1911] : 
                       (N93)? mem[1960] : 
                       (N95)? mem[2009] : 
                       (N97)? mem[2058] : 
                       (N99)? mem[2107] : 
                       (N101)? mem[2156] : 
                       (N103)? mem[2205] : 
                       (N105)? mem[2254] : 
                       (N107)? mem[2303] : 
                       (N109)? mem[2352] : 
                       (N111)? mem[2401] : 
                       (N113)? mem[2450] : 
                       (N115)? mem[2499] : 
                       (N117)? mem[2548] : 
                       (N119)? mem[2597] : 
                       (N121)? mem[2646] : 
                       (N123)? mem[2695] : 
                       (N125)? mem[2744] : 
                       (N127)? mem[2793] : 
                       (N129)? mem[2842] : 
                       (N131)? mem[2891] : 
                       (N133)? mem[2940] : 
                       (N135)? mem[2989] : 
                       (N137)? mem[3038] : 
                       (N139)? mem[3087] : 1'b0;
  assign N269 = ~w_addr_i[5];
  assign N270 = w_addr_i[3] & w_addr_i[4];
  assign N271 = N0 & w_addr_i[4];
  assign N0 = ~w_addr_i[3];
  assign N272 = w_addr_i[3] & N1;
  assign N1 = ~w_addr_i[4];
  assign N273 = N2 & N3;
  assign N2 = ~w_addr_i[3];
  assign N3 = ~w_addr_i[4];
  assign N274 = w_addr_i[5] & N270;
  assign N275 = w_addr_i[5] & N271;
  assign N276 = w_addr_i[5] & N272;
  assign N277 = w_addr_i[5] & N273;
  assign N278 = N269 & N270;
  assign N279 = N269 & N271;
  assign N280 = N269 & N272;
  assign N281 = N269 & N273;
  assign N282 = ~w_addr_i[2];
  assign N283 = w_addr_i[0] & w_addr_i[1];
  assign N284 = N4 & w_addr_i[1];
  assign N4 = ~w_addr_i[0];
  assign N285 = w_addr_i[0] & N5;
  assign N5 = ~w_addr_i[1];
  assign N286 = N6 & N7;
  assign N6 = ~w_addr_i[0];
  assign N7 = ~w_addr_i[1];
  assign N287 = w_addr_i[2] & N283;
  assign N288 = w_addr_i[2] & N284;
  assign N289 = w_addr_i[2] & N285;
  assign N290 = w_addr_i[2] & N286;
  assign N291 = N282 & N283;
  assign N292 = N282 & N284;
  assign N293 = N282 & N285;
  assign N294 = N282 & N286;
  assign N204 = N274 & N287;
  assign N203 = N274 & N288;
  assign N202 = N274 & N289;
  assign N201 = N274 & N290;
  assign N200 = N274 & N291;
  assign N199 = N274 & N292;
  assign N198 = N274 & N293;
  assign N197 = N274 & N294;
  assign N196 = N275 & N287;
  assign N195 = N275 & N288;
  assign N194 = N275 & N289;
  assign N193 = N275 & N290;
  assign N192 = N275 & N291;
  assign N191 = N275 & N292;
  assign N190 = N275 & N293;
  assign N189 = N275 & N294;
  assign N188 = N276 & N287;
  assign N187 = N276 & N288;
  assign N186 = N276 & N289;
  assign N185 = N276 & N290;
  assign N184 = N276 & N291;
  assign N183 = N276 & N292;
  assign N182 = N276 & N293;
  assign N181 = N276 & N294;
  assign N180 = N277 & N287;
  assign N179 = N277 & N288;
  assign N178 = N277 & N289;
  assign N177 = N277 & N290;
  assign N176 = N277 & N291;
  assign N175 = N277 & N292;
  assign N174 = N277 & N293;
  assign N173 = N277 & N294;
  assign N172 = N278 & N287;
  assign N171 = N278 & N288;
  assign N170 = N278 & N289;
  assign N169 = N278 & N290;
  assign N168 = N278 & N291;
  assign N167 = N278 & N292;
  assign N166 = N278 & N293;
  assign N165 = N278 & N294;
  assign N164 = N279 & N287;
  assign N163 = N279 & N288;
  assign N162 = N279 & N289;
  assign N161 = N279 & N290;
  assign N160 = N279 & N291;
  assign N159 = N279 & N292;
  assign N158 = N279 & N293;
  assign N157 = N279 & N294;
  assign N156 = N280 & N287;
  assign N155 = N280 & N288;
  assign N154 = N280 & N289;
  assign N153 = N280 & N290;
  assign N152 = N280 & N291;
  assign N151 = N280 & N292;
  assign N150 = N280 & N293;
  assign N149 = N280 & N294;
  assign N148 = N281 & N287;
  assign N147 = N281 & N288;
  assign N146 = N281 & N289;
  assign N145 = N281 & N290;
  assign N144 = N281 & N291;
  assign N143 = N281 & N292;
  assign N142 = N281 & N293;
  assign N141 = N281 & N294;
  assign { N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205 } = (N8)? { N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N9)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N8 = w_v_i;
  assign N9 = N140;
  assign N10 = ~r_addr_i[0];
  assign N11 = ~r_addr_i[1];
  assign N12 = N10 & N11;
  assign N13 = N10 & r_addr_i[1];
  assign N14 = r_addr_i[0] & N11;
  assign N15 = r_addr_i[0] & r_addr_i[1];
  assign N16 = ~r_addr_i[2];
  assign N17 = N12 & N16;
  assign N18 = N12 & r_addr_i[2];
  assign N19 = N14 & N16;
  assign N20 = N14 & r_addr_i[2];
  assign N21 = N13 & N16;
  assign N22 = N13 & r_addr_i[2];
  assign N23 = N15 & N16;
  assign N24 = N15 & r_addr_i[2];
  assign N25 = ~r_addr_i[3];
  assign N26 = N17 & N25;
  assign N27 = N17 & r_addr_i[3];
  assign N28 = N19 & N25;
  assign N29 = N19 & r_addr_i[3];
  assign N30 = N21 & N25;
  assign N31 = N21 & r_addr_i[3];
  assign N32 = N23 & N25;
  assign N33 = N23 & r_addr_i[3];
  assign N34 = N18 & N25;
  assign N35 = N18 & r_addr_i[3];
  assign N36 = N20 & N25;
  assign N37 = N20 & r_addr_i[3];
  assign N38 = N22 & N25;
  assign N39 = N22 & r_addr_i[3];
  assign N40 = N24 & N25;
  assign N41 = N24 & r_addr_i[3];
  assign N42 = ~r_addr_i[4];
  assign N43 = N26 & N42;
  assign N44 = N26 & r_addr_i[4];
  assign N45 = N28 & N42;
  assign N46 = N28 & r_addr_i[4];
  assign N47 = N30 & N42;
  assign N48 = N30 & r_addr_i[4];
  assign N49 = N32 & N42;
  assign N50 = N32 & r_addr_i[4];
  assign N51 = N34 & N42;
  assign N52 = N34 & r_addr_i[4];
  assign N53 = N36 & N42;
  assign N54 = N36 & r_addr_i[4];
  assign N55 = N38 & N42;
  assign N56 = N38 & r_addr_i[4];
  assign N57 = N40 & N42;
  assign N58 = N40 & r_addr_i[4];
  assign N59 = N27 & N42;
  assign N60 = N27 & r_addr_i[4];
  assign N61 = N29 & N42;
  assign N62 = N29 & r_addr_i[4];
  assign N63 = N31 & N42;
  assign N64 = N31 & r_addr_i[4];
  assign N65 = N33 & N42;
  assign N66 = N33 & r_addr_i[4];
  assign N67 = N35 & N42;
  assign N68 = N35 & r_addr_i[4];
  assign N69 = N37 & N42;
  assign N70 = N37 & r_addr_i[4];
  assign N71 = N39 & N42;
  assign N72 = N39 & r_addr_i[4];
  assign N73 = N41 & N42;
  assign N74 = N41 & r_addr_i[4];
  assign N75 = ~r_addr_i[5];
  assign N76 = N43 & N75;
  assign N77 = N43 & r_addr_i[5];
  assign N78 = N45 & N75;
  assign N79 = N45 & r_addr_i[5];
  assign N80 = N47 & N75;
  assign N81 = N47 & r_addr_i[5];
  assign N82 = N49 & N75;
  assign N83 = N49 & r_addr_i[5];
  assign N84 = N51 & N75;
  assign N85 = N51 & r_addr_i[5];
  assign N86 = N53 & N75;
  assign N87 = N53 & r_addr_i[5];
  assign N88 = N55 & N75;
  assign N89 = N55 & r_addr_i[5];
  assign N90 = N57 & N75;
  assign N91 = N57 & r_addr_i[5];
  assign N92 = N59 & N75;
  assign N93 = N59 & r_addr_i[5];
  assign N94 = N61 & N75;
  assign N95 = N61 & r_addr_i[5];
  assign N96 = N63 & N75;
  assign N97 = N63 & r_addr_i[5];
  assign N98 = N65 & N75;
  assign N99 = N65 & r_addr_i[5];
  assign N100 = N67 & N75;
  assign N101 = N67 & r_addr_i[5];
  assign N102 = N69 & N75;
  assign N103 = N69 & r_addr_i[5];
  assign N104 = N71 & N75;
  assign N105 = N71 & r_addr_i[5];
  assign N106 = N73 & N75;
  assign N107 = N73 & r_addr_i[5];
  assign N108 = N44 & N75;
  assign N109 = N44 & r_addr_i[5];
  assign N110 = N46 & N75;
  assign N111 = N46 & r_addr_i[5];
  assign N112 = N48 & N75;
  assign N113 = N48 & r_addr_i[5];
  assign N114 = N50 & N75;
  assign N115 = N50 & r_addr_i[5];
  assign N116 = N52 & N75;
  assign N117 = N52 & r_addr_i[5];
  assign N118 = N54 & N75;
  assign N119 = N54 & r_addr_i[5];
  assign N120 = N56 & N75;
  assign N121 = N56 & r_addr_i[5];
  assign N122 = N58 & N75;
  assign N123 = N58 & r_addr_i[5];
  assign N124 = N60 & N75;
  assign N125 = N60 & r_addr_i[5];
  assign N126 = N62 & N75;
  assign N127 = N62 & r_addr_i[5];
  assign N128 = N64 & N75;
  assign N129 = N64 & r_addr_i[5];
  assign N130 = N66 & N75;
  assign N131 = N66 & r_addr_i[5];
  assign N132 = N68 & N75;
  assign N133 = N68 & r_addr_i[5];
  assign N134 = N70 & N75;
  assign N135 = N70 & r_addr_i[5];
  assign N136 = N72 & N75;
  assign N137 = N72 & r_addr_i[5];
  assign N138 = N74 & N75;
  assign N139 = N74 & r_addr_i[5];
  assign N140 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N268) begin
      { mem[3135:3087] } <= { w_data_i[48:0] };
    end 
    if(N267) begin
      { mem[3086:3038] } <= { w_data_i[48:0] };
    end 
    if(N266) begin
      { mem[3037:2989] } <= { w_data_i[48:0] };
    end 
    if(N265) begin
      { mem[2988:2940] } <= { w_data_i[48:0] };
    end 
    if(N264) begin
      { mem[2939:2891] } <= { w_data_i[48:0] };
    end 
    if(N263) begin
      { mem[2890:2842] } <= { w_data_i[48:0] };
    end 
    if(N262) begin
      { mem[2841:2793] } <= { w_data_i[48:0] };
    end 
    if(N261) begin
      { mem[2792:2744] } <= { w_data_i[48:0] };
    end 
    if(N260) begin
      { mem[2743:2695] } <= { w_data_i[48:0] };
    end 
    if(N259) begin
      { mem[2694:2646] } <= { w_data_i[48:0] };
    end 
    if(N258) begin
      { mem[2645:2597] } <= { w_data_i[48:0] };
    end 
    if(N257) begin
      { mem[2596:2548] } <= { w_data_i[48:0] };
    end 
    if(N256) begin
      { mem[2547:2499] } <= { w_data_i[48:0] };
    end 
    if(N255) begin
      { mem[2498:2450] } <= { w_data_i[48:0] };
    end 
    if(N254) begin
      { mem[2449:2401] } <= { w_data_i[48:0] };
    end 
    if(N253) begin
      { mem[2400:2352] } <= { w_data_i[48:0] };
    end 
    if(N252) begin
      { mem[2351:2303] } <= { w_data_i[48:0] };
    end 
    if(N251) begin
      { mem[2302:2254] } <= { w_data_i[48:0] };
    end 
    if(N250) begin
      { mem[2253:2205] } <= { w_data_i[48:0] };
    end 
    if(N249) begin
      { mem[2204:2156] } <= { w_data_i[48:0] };
    end 
    if(N248) begin
      { mem[2155:2107] } <= { w_data_i[48:0] };
    end 
    if(N247) begin
      { mem[2106:2058] } <= { w_data_i[48:0] };
    end 
    if(N246) begin
      { mem[2057:2009] } <= { w_data_i[48:0] };
    end 
    if(N245) begin
      { mem[2008:1960] } <= { w_data_i[48:0] };
    end 
    if(N244) begin
      { mem[1959:1911] } <= { w_data_i[48:0] };
    end 
    if(N243) begin
      { mem[1910:1862] } <= { w_data_i[48:0] };
    end 
    if(N242) begin
      { mem[1861:1813] } <= { w_data_i[48:0] };
    end 
    if(N241) begin
      { mem[1812:1764] } <= { w_data_i[48:0] };
    end 
    if(N240) begin
      { mem[1763:1715] } <= { w_data_i[48:0] };
    end 
    if(N239) begin
      { mem[1714:1666] } <= { w_data_i[48:0] };
    end 
    if(N238) begin
      { mem[1665:1617] } <= { w_data_i[48:0] };
    end 
    if(N237) begin
      { mem[1616:1568] } <= { w_data_i[48:0] };
    end 
    if(N236) begin
      { mem[1567:1519] } <= { w_data_i[48:0] };
    end 
    if(N235) begin
      { mem[1518:1470] } <= { w_data_i[48:0] };
    end 
    if(N234) begin
      { mem[1469:1421] } <= { w_data_i[48:0] };
    end 
    if(N233) begin
      { mem[1420:1372] } <= { w_data_i[48:0] };
    end 
    if(N232) begin
      { mem[1371:1323] } <= { w_data_i[48:0] };
    end 
    if(N231) begin
      { mem[1322:1274] } <= { w_data_i[48:0] };
    end 
    if(N230) begin
      { mem[1273:1225] } <= { w_data_i[48:0] };
    end 
    if(N229) begin
      { mem[1224:1176] } <= { w_data_i[48:0] };
    end 
    if(N228) begin
      { mem[1175:1127] } <= { w_data_i[48:0] };
    end 
    if(N227) begin
      { mem[1126:1078] } <= { w_data_i[48:0] };
    end 
    if(N226) begin
      { mem[1077:1029] } <= { w_data_i[48:0] };
    end 
    if(N225) begin
      { mem[1028:980] } <= { w_data_i[48:0] };
    end 
    if(N224) begin
      { mem[979:931] } <= { w_data_i[48:0] };
    end 
    if(N223) begin
      { mem[930:882] } <= { w_data_i[48:0] };
    end 
    if(N222) begin
      { mem[881:833] } <= { w_data_i[48:0] };
    end 
    if(N221) begin
      { mem[832:784] } <= { w_data_i[48:0] };
    end 
    if(N220) begin
      { mem[783:735] } <= { w_data_i[48:0] };
    end 
    if(N219) begin
      { mem[734:686] } <= { w_data_i[48:0] };
    end 
    if(N218) begin
      { mem[685:637] } <= { w_data_i[48:0] };
    end 
    if(N217) begin
      { mem[636:588] } <= { w_data_i[48:0] };
    end 
    if(N216) begin
      { mem[587:539] } <= { w_data_i[48:0] };
    end 
    if(N215) begin
      { mem[538:490] } <= { w_data_i[48:0] };
    end 
    if(N214) begin
      { mem[489:441] } <= { w_data_i[48:0] };
    end 
    if(N213) begin
      { mem[440:392] } <= { w_data_i[48:0] };
    end 
    if(N212) begin
      { mem[391:343] } <= { w_data_i[48:0] };
    end 
    if(N211) begin
      { mem[342:294] } <= { w_data_i[48:0] };
    end 
    if(N210) begin
      { mem[293:245] } <= { w_data_i[48:0] };
    end 
    if(N209) begin
      { mem[244:196] } <= { w_data_i[48:0] };
    end 
    if(N208) begin
      { mem[195:147] } <= { w_data_i[48:0] };
    end 
    if(N207) begin
      { mem[146:98] } <= { w_data_i[48:0] };
    end 
    if(N206) begin
      { mem[97:49] } <= { w_data_i[48:0] };
    end 
    if(N205) begin
      { mem[48:0] } <= { w_data_i[48:0] };
    end 
  end


endmodule



module bsg_mem_1r1w_width_p49_els_p64_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [5:0] w_addr_i;
  input [48:0] w_data_i;
  input [5:0] r_addr_i;
  output [48:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [48:0] r_data_o;

  bsg_mem_1r1w_synth_width_p49_els_p64_read_write_same_addr_p0_harden_p0
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_mem_1rw_sync_width_p49_els_p64
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_i,
  data_o
);

  input [48:0] data_i;
  input [5:0] addr_i;
  output [48:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire n_0_net_,n_1_net_,N0;
  wire [48:0] z_s1r1w_data_lo;
  reg [48:0] data_o;

  bsg_mem_1r1w_width_p49_els_p64_read_write_same_addr_p0
  z_s1r1w_mem
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(n_0_net_),
    .w_addr_i(addr_i),
    .w_data_i(data_i),
    .r_v_i(n_1_net_),
    .r_addr_i(addr_i),
    .r_data_o(z_s1r1w_data_lo)
  );

  assign n_1_net_ = v_i & N0;
  assign N0 = ~w_i;
  assign n_0_net_ = v_i & w_i;

  always @(posedge clk_i) begin
    if(1'b1) begin
      { data_o[48:0] } <= { z_s1r1w_data_lo[48:0] };
    end 
  end


endmodule



module bp_fe_btb_vaddr_width_p39_btb_tag_width_p10_btb_idx_width_p6
(
  clk_i,
  reset_i,
  r_addr_i,
  r_v_i,
  br_tgt_o,
  br_tgt_v_o,
  w_tag_i,
  w_idx_i,
  w_v_i,
  br_tgt_i
);

  input [38:0] r_addr_i;
  output [38:0] br_tgt_o;
  input [9:0] w_tag_i;
  input [5:0] w_idx_i;
  input [38:0] br_tgt_i;
  input clk_i;
  input reset_i;
  input r_v_i;
  input w_v_i;
  output br_tgt_v_o;
  wire [38:0] br_tgt_o;
  wire br_tgt_v_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,n_0_net_,N15,N16,
  N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,
  N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,
  N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,
  N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,
  N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,
  N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,
  N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,
  tag_mem_v_lo,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,
  N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,
  N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,
  N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,
  N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,
  N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,
  N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,
  N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,
  N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,
  N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,
  N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,
  N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,
  N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,
  N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,
  N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,
  N383,N384,N385,N386,N387,N388,N389,N390,N391,N392;
  wire [5:0] tag_mem_addr_li;
  wire [9:0] tag_mem_lo;
  reg [5:0] r_idx_r;
  reg r_v_r;
  reg [9:0] r_tag_r;
  reg [63:0] v_r;

  bsg_mem_1rw_sync_width_p49_els_p64
  tag_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i({ w_tag_i, br_tgt_i }),
    .addr_i(tag_mem_addr_li),
    .v_i(n_0_net_),
    .w_i(w_v_i),
    .data_o({ tag_mem_lo, br_tgt_o })
  );

  assign tag_mem_v_lo = (N81)? v_r[0] : 
                        (N83)? v_r[1] : 
                        (N85)? v_r[2] : 
                        (N87)? v_r[3] : 
                        (N89)? v_r[4] : 
                        (N91)? v_r[5] : 
                        (N93)? v_r[6] : 
                        (N95)? v_r[7] : 
                        (N97)? v_r[8] : 
                        (N99)? v_r[9] : 
                        (N101)? v_r[10] : 
                        (N103)? v_r[11] : 
                        (N105)? v_r[12] : 
                        (N107)? v_r[13] : 
                        (N109)? v_r[14] : 
                        (N111)? v_r[15] : 
                        (N113)? v_r[16] : 
                        (N115)? v_r[17] : 
                        (N117)? v_r[18] : 
                        (N119)? v_r[19] : 
                        (N121)? v_r[20] : 
                        (N123)? v_r[21] : 
                        (N125)? v_r[22] : 
                        (N127)? v_r[23] : 
                        (N129)? v_r[24] : 
                        (N131)? v_r[25] : 
                        (N133)? v_r[26] : 
                        (N135)? v_r[27] : 
                        (N137)? v_r[28] : 
                        (N139)? v_r[29] : 
                        (N141)? v_r[30] : 
                        (N143)? v_r[31] : 
                        (N82)? v_r[32] : 
                        (N84)? v_r[33] : 
                        (N86)? v_r[34] : 
                        (N88)? v_r[35] : 
                        (N90)? v_r[36] : 
                        (N92)? v_r[37] : 
                        (N94)? v_r[38] : 
                        (N96)? v_r[39] : 
                        (N98)? v_r[40] : 
                        (N100)? v_r[41] : 
                        (N102)? v_r[42] : 
                        (N104)? v_r[43] : 
                        (N106)? v_r[44] : 
                        (N108)? v_r[45] : 
                        (N110)? v_r[46] : 
                        (N112)? v_r[47] : 
                        (N114)? v_r[48] : 
                        (N116)? v_r[49] : 
                        (N118)? v_r[50] : 
                        (N120)? v_r[51] : 
                        (N122)? v_r[52] : 
                        (N124)? v_r[53] : 
                        (N126)? v_r[54] : 
                        (N128)? v_r[55] : 
                        (N130)? v_r[56] : 
                        (N132)? v_r[57] : 
                        (N134)? v_r[58] : 
                        (N136)? v_r[59] : 
                        (N138)? v_r[60] : 
                        (N140)? v_r[61] : 
                        (N142)? v_r[62] : 
                        (N144)? v_r[63] : 1'b0;
  assign N145 = tag_mem_lo == r_tag_r;
  assign N365 = ~tag_mem_addr_li[5];
  assign N366 = tag_mem_addr_li[3] & tag_mem_addr_li[4];
  assign N367 = N0 & tag_mem_addr_li[4];
  assign N0 = ~tag_mem_addr_li[3];
  assign N368 = tag_mem_addr_li[3] & N1;
  assign N1 = ~tag_mem_addr_li[4];
  assign N369 = N2 & N3;
  assign N2 = ~tag_mem_addr_li[3];
  assign N3 = ~tag_mem_addr_li[4];
  assign N370 = tag_mem_addr_li[5] & N366;
  assign N371 = tag_mem_addr_li[5] & N367;
  assign N372 = tag_mem_addr_li[5] & N368;
  assign N373 = tag_mem_addr_li[5] & N369;
  assign N374 = N365 & N366;
  assign N375 = N365 & N367;
  assign N376 = N365 & N368;
  assign N377 = N365 & N369;
  assign N378 = ~tag_mem_addr_li[2];
  assign N379 = tag_mem_addr_li[0] & tag_mem_addr_li[1];
  assign N380 = N4 & tag_mem_addr_li[1];
  assign N4 = ~tag_mem_addr_li[0];
  assign N381 = tag_mem_addr_li[0] & N5;
  assign N5 = ~tag_mem_addr_li[1];
  assign N382 = N6 & N7;
  assign N6 = ~tag_mem_addr_li[0];
  assign N7 = ~tag_mem_addr_li[1];
  assign N383 = tag_mem_addr_li[2] & N379;
  assign N384 = tag_mem_addr_li[2] & N380;
  assign N385 = tag_mem_addr_li[2] & N381;
  assign N386 = tag_mem_addr_li[2] & N382;
  assign N387 = N378 & N379;
  assign N388 = N378 & N380;
  assign N389 = N378 & N381;
  assign N390 = N378 & N382;
  assign N233 = N370 & N383;
  assign N232 = N370 & N384;
  assign N231 = N370 & N385;
  assign N230 = N370 & N386;
  assign N229 = N370 & N387;
  assign N228 = N370 & N388;
  assign N227 = N370 & N389;
  assign N226 = N370 & N390;
  assign N225 = N371 & N383;
  assign N224 = N371 & N384;
  assign N223 = N371 & N385;
  assign N222 = N371 & N386;
  assign N221 = N371 & N387;
  assign N220 = N371 & N388;
  assign N219 = N371 & N389;
  assign N218 = N371 & N390;
  assign N217 = N372 & N383;
  assign N216 = N372 & N384;
  assign N215 = N372 & N385;
  assign N214 = N372 & N386;
  assign N213 = N372 & N387;
  assign N212 = N372 & N388;
  assign N211 = N372 & N389;
  assign N210 = N372 & N390;
  assign N209 = N373 & N383;
  assign N208 = N373 & N384;
  assign N207 = N373 & N385;
  assign N206 = N373 & N386;
  assign N205 = N373 & N387;
  assign N204 = N373 & N388;
  assign N203 = N373 & N389;
  assign N202 = N373 & N390;
  assign N201 = N374 & N383;
  assign N200 = N374 & N384;
  assign N199 = N374 & N385;
  assign N198 = N374 & N386;
  assign N197 = N374 & N387;
  assign N196 = N374 & N388;
  assign N195 = N374 & N389;
  assign N194 = N374 & N390;
  assign N193 = N375 & N383;
  assign N192 = N375 & N384;
  assign N191 = N375 & N385;
  assign N190 = N375 & N386;
  assign N189 = N375 & N387;
  assign N188 = N375 & N388;
  assign N187 = N375 & N389;
  assign N186 = N375 & N390;
  assign N185 = N376 & N383;
  assign N184 = N376 & N384;
  assign N183 = N376 & N385;
  assign N182 = N376 & N386;
  assign N181 = N376 & N387;
  assign N180 = N376 & N388;
  assign N179 = N376 & N389;
  assign N178 = N376 & N390;
  assign N177 = N377 & N383;
  assign N176 = N377 & N384;
  assign N175 = N377 & N385;
  assign N174 = N377 & N386;
  assign N173 = N377 & N387;
  assign N172 = N377 & N388;
  assign N171 = N377 & N389;
  assign N170 = N377 & N390;
  assign tag_mem_addr_li = (N8)? w_idx_i : 
                           (N9)? r_addr_i[7:2] : 1'b0;
  assign N8 = N14;
  assign N9 = N13;
  assign N149 = (N10)? 1'b0 : 
                (N11)? N148 : 1'b0;
  assign N10 = N147;
  assign N11 = N146;
  assign { N159, N158, N157, N156, N155, N154, N153, N152, N151, N150 } = (N10)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                          (N11)? r_addr_i[17:8] : 1'b0;
  assign { N165, N164, N163, N162, N161, N160 } = (N10)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                  (N11)? r_addr_i[7:2] : 1'b0;
  assign { N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N234 } = (N12)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N300)? { N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N169)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign N12 = N166;
  assign N235 = (N12)? 1'b0 : 
                (N300)? 1'b1 : 1'b0;
  assign N13 = ~w_v_i;
  assign N14 = w_v_i;
  assign n_0_net_ = r_v_i | w_v_i;
  assign N15 = ~r_idx_r[0];
  assign N16 = ~r_idx_r[1];
  assign N17 = N15 & N16;
  assign N18 = N15 & r_idx_r[1];
  assign N19 = r_idx_r[0] & N16;
  assign N20 = r_idx_r[0] & r_idx_r[1];
  assign N21 = ~r_idx_r[2];
  assign N22 = N17 & N21;
  assign N23 = N17 & r_idx_r[2];
  assign N24 = N19 & N21;
  assign N25 = N19 & r_idx_r[2];
  assign N26 = N18 & N21;
  assign N27 = N18 & r_idx_r[2];
  assign N28 = N20 & N21;
  assign N29 = N20 & r_idx_r[2];
  assign N30 = ~r_idx_r[3];
  assign N31 = N22 & N30;
  assign N32 = N22 & r_idx_r[3];
  assign N33 = N24 & N30;
  assign N34 = N24 & r_idx_r[3];
  assign N35 = N26 & N30;
  assign N36 = N26 & r_idx_r[3];
  assign N37 = N28 & N30;
  assign N38 = N28 & r_idx_r[3];
  assign N39 = N23 & N30;
  assign N40 = N23 & r_idx_r[3];
  assign N41 = N25 & N30;
  assign N42 = N25 & r_idx_r[3];
  assign N43 = N27 & N30;
  assign N44 = N27 & r_idx_r[3];
  assign N45 = N29 & N30;
  assign N46 = N29 & r_idx_r[3];
  assign N47 = ~r_idx_r[4];
  assign N48 = N31 & N47;
  assign N49 = N31 & r_idx_r[4];
  assign N50 = N33 & N47;
  assign N51 = N33 & r_idx_r[4];
  assign N52 = N35 & N47;
  assign N53 = N35 & r_idx_r[4];
  assign N54 = N37 & N47;
  assign N55 = N37 & r_idx_r[4];
  assign N56 = N39 & N47;
  assign N57 = N39 & r_idx_r[4];
  assign N58 = N41 & N47;
  assign N59 = N41 & r_idx_r[4];
  assign N60 = N43 & N47;
  assign N61 = N43 & r_idx_r[4];
  assign N62 = N45 & N47;
  assign N63 = N45 & r_idx_r[4];
  assign N64 = N32 & N47;
  assign N65 = N32 & r_idx_r[4];
  assign N66 = N34 & N47;
  assign N67 = N34 & r_idx_r[4];
  assign N68 = N36 & N47;
  assign N69 = N36 & r_idx_r[4];
  assign N70 = N38 & N47;
  assign N71 = N38 & r_idx_r[4];
  assign N72 = N40 & N47;
  assign N73 = N40 & r_idx_r[4];
  assign N74 = N42 & N47;
  assign N75 = N42 & r_idx_r[4];
  assign N76 = N44 & N47;
  assign N77 = N44 & r_idx_r[4];
  assign N78 = N46 & N47;
  assign N79 = N46 & r_idx_r[4];
  assign N80 = ~r_idx_r[5];
  assign N81 = N48 & N80;
  assign N82 = N48 & r_idx_r[5];
  assign N83 = N50 & N80;
  assign N84 = N50 & r_idx_r[5];
  assign N85 = N52 & N80;
  assign N86 = N52 & r_idx_r[5];
  assign N87 = N54 & N80;
  assign N88 = N54 & r_idx_r[5];
  assign N89 = N56 & N80;
  assign N90 = N56 & r_idx_r[5];
  assign N91 = N58 & N80;
  assign N92 = N58 & r_idx_r[5];
  assign N93 = N60 & N80;
  assign N94 = N60 & r_idx_r[5];
  assign N95 = N62 & N80;
  assign N96 = N62 & r_idx_r[5];
  assign N97 = N64 & N80;
  assign N98 = N64 & r_idx_r[5];
  assign N99 = N66 & N80;
  assign N100 = N66 & r_idx_r[5];
  assign N101 = N68 & N80;
  assign N102 = N68 & r_idx_r[5];
  assign N103 = N70 & N80;
  assign N104 = N70 & r_idx_r[5];
  assign N105 = N72 & N80;
  assign N106 = N72 & r_idx_r[5];
  assign N107 = N74 & N80;
  assign N108 = N74 & r_idx_r[5];
  assign N109 = N76 & N80;
  assign N110 = N76 & r_idx_r[5];
  assign N111 = N78 & N80;
  assign N112 = N78 & r_idx_r[5];
  assign N113 = N49 & N80;
  assign N114 = N49 & r_idx_r[5];
  assign N115 = N51 & N80;
  assign N116 = N51 & r_idx_r[5];
  assign N117 = N53 & N80;
  assign N118 = N53 & r_idx_r[5];
  assign N119 = N55 & N80;
  assign N120 = N55 & r_idx_r[5];
  assign N121 = N57 & N80;
  assign N122 = N57 & r_idx_r[5];
  assign N123 = N59 & N80;
  assign N124 = N59 & r_idx_r[5];
  assign N125 = N61 & N80;
  assign N126 = N61 & r_idx_r[5];
  assign N127 = N63 & N80;
  assign N128 = N63 & r_idx_r[5];
  assign N129 = N65 & N80;
  assign N130 = N65 & r_idx_r[5];
  assign N131 = N67 & N80;
  assign N132 = N67 & r_idx_r[5];
  assign N133 = N69 & N80;
  assign N134 = N69 & r_idx_r[5];
  assign N135 = N71 & N80;
  assign N136 = N71 & r_idx_r[5];
  assign N137 = N73 & N80;
  assign N138 = N73 & r_idx_r[5];
  assign N139 = N75 & N80;
  assign N140 = N75 & r_idx_r[5];
  assign N141 = N77 & N80;
  assign N142 = N77 & r_idx_r[5];
  assign N143 = N79 & N80;
  assign N144 = N79 & r_idx_r[5];
  assign br_tgt_v_o = N391 & N145;
  assign N391 = tag_mem_v_lo & r_v_r;
  assign N146 = ~reset_i;
  assign N147 = reset_i;
  assign N148 = r_v_i & N392;
  assign N392 = ~w_v_i;
  assign N166 = reset_i;
  assign N167 = w_v_i;
  assign N168 = N167 | N166;
  assign N169 = ~N168;
  assign N299 = ~N166;
  assign N300 = N167 & N299;
  assign N301 = N298 & N168;
  assign N302 = N297 & N168;
  assign N303 = N296 & N168;
  assign N304 = N295 & N168;
  assign N305 = N294 & N168;
  assign N306 = N293 & N168;
  assign N307 = N292 & N168;
  assign N308 = N291 & N168;
  assign N309 = N290 & N168;
  assign N310 = N289 & N168;
  assign N311 = N288 & N168;
  assign N312 = N287 & N168;
  assign N313 = N286 & N168;
  assign N314 = N285 & N168;
  assign N315 = N284 & N168;
  assign N316 = N283 & N168;
  assign N317 = N282 & N168;
  assign N318 = N281 & N168;
  assign N319 = N280 & N168;
  assign N320 = N279 & N168;
  assign N321 = N278 & N168;
  assign N322 = N277 & N168;
  assign N323 = N276 & N168;
  assign N324 = N275 & N168;
  assign N325 = N274 & N168;
  assign N326 = N273 & N168;
  assign N327 = N272 & N168;
  assign N328 = N271 & N168;
  assign N329 = N270 & N168;
  assign N330 = N269 & N168;
  assign N331 = N268 & N168;
  assign N332 = N267 & N168;
  assign N333 = N266 & N168;
  assign N334 = N265 & N168;
  assign N335 = N264 & N168;
  assign N336 = N263 & N168;
  assign N337 = N262 & N168;
  assign N338 = N261 & N168;
  assign N339 = N260 & N168;
  assign N340 = N259 & N168;
  assign N341 = N258 & N168;
  assign N342 = N257 & N168;
  assign N343 = N256 & N168;
  assign N344 = N255 & N168;
  assign N345 = N254 & N168;
  assign N346 = N253 & N168;
  assign N347 = N252 & N168;
  assign N348 = N251 & N168;
  assign N349 = N250 & N168;
  assign N350 = N249 & N168;
  assign N351 = N248 & N168;
  assign N352 = N247 & N168;
  assign N353 = N246 & N168;
  assign N354 = N245 & N168;
  assign N355 = N244 & N168;
  assign N356 = N243 & N168;
  assign N357 = N242 & N168;
  assign N358 = N241 & N168;
  assign N359 = N240 & N168;
  assign N360 = N239 & N168;
  assign N361 = N238 & N168;
  assign N362 = N237 & N168;
  assign N363 = N236 & N168;
  assign N364 = N234 & N168;

  always @(posedge clk_i) begin
    if(1'b1) begin
      { r_idx_r[5:0] } <= { N165, N164, N163, N162, N161, N160 };
      r_v_r <= N149;
      { r_tag_r[9:0] } <= { N159, N158, N157, N156, N155, N154, N153, N152, N151, N150 };
    end 
    if(N301) begin
      { v_r[63:63] } <= { N235 };
    end 
    if(N302) begin
      { v_r[62:62] } <= { N235 };
    end 
    if(N303) begin
      { v_r[61:61] } <= { N235 };
    end 
    if(N304) begin
      { v_r[60:60] } <= { N235 };
    end 
    if(N305) begin
      { v_r[59:59] } <= { N235 };
    end 
    if(N306) begin
      { v_r[58:58] } <= { N235 };
    end 
    if(N307) begin
      { v_r[57:57] } <= { N235 };
    end 
    if(N308) begin
      { v_r[56:56] } <= { N235 };
    end 
    if(N309) begin
      { v_r[55:55] } <= { N235 };
    end 
    if(N310) begin
      { v_r[54:54] } <= { N235 };
    end 
    if(N311) begin
      { v_r[53:53] } <= { N235 };
    end 
    if(N312) begin
      { v_r[52:52] } <= { N235 };
    end 
    if(N313) begin
      { v_r[51:51] } <= { N235 };
    end 
    if(N314) begin
      { v_r[50:50] } <= { N235 };
    end 
    if(N315) begin
      { v_r[49:49] } <= { N235 };
    end 
    if(N316) begin
      { v_r[48:48] } <= { N235 };
    end 
    if(N317) begin
      { v_r[47:47] } <= { N235 };
    end 
    if(N318) begin
      { v_r[46:46] } <= { N235 };
    end 
    if(N319) begin
      { v_r[45:45] } <= { N235 };
    end 
    if(N320) begin
      { v_r[44:44] } <= { N235 };
    end 
    if(N321) begin
      { v_r[43:43] } <= { N235 };
    end 
    if(N322) begin
      { v_r[42:42] } <= { N235 };
    end 
    if(N323) begin
      { v_r[41:41] } <= { N235 };
    end 
    if(N324) begin
      { v_r[40:40] } <= { N235 };
    end 
    if(N325) begin
      { v_r[39:39] } <= { N235 };
    end 
    if(N326) begin
      { v_r[38:38] } <= { N235 };
    end 
    if(N327) begin
      { v_r[37:37] } <= { N235 };
    end 
    if(N328) begin
      { v_r[36:36] } <= { N235 };
    end 
    if(N329) begin
      { v_r[35:35] } <= { N235 };
    end 
    if(N330) begin
      { v_r[34:34] } <= { N235 };
    end 
    if(N331) begin
      { v_r[33:33] } <= { N235 };
    end 
    if(N332) begin
      { v_r[32:32] } <= { N235 };
    end 
    if(N333) begin
      { v_r[31:31] } <= { N235 };
    end 
    if(N334) begin
      { v_r[30:30] } <= { N235 };
    end 
    if(N335) begin
      { v_r[29:29] } <= { N235 };
    end 
    if(N336) begin
      { v_r[28:28] } <= { N235 };
    end 
    if(N337) begin
      { v_r[27:27] } <= { N235 };
    end 
    if(N338) begin
      { v_r[26:26] } <= { N235 };
    end 
    if(N339) begin
      { v_r[25:25] } <= { N235 };
    end 
    if(N340) begin
      { v_r[24:24] } <= { N235 };
    end 
    if(N341) begin
      { v_r[23:23] } <= { N235 };
    end 
    if(N342) begin
      { v_r[22:22] } <= { N235 };
    end 
    if(N343) begin
      { v_r[21:21] } <= { N235 };
    end 
    if(N344) begin
      { v_r[20:20] } <= { N235 };
    end 
    if(N345) begin
      { v_r[19:19] } <= { N235 };
    end 
    if(N346) begin
      { v_r[18:18] } <= { N235 };
    end 
    if(N347) begin
      { v_r[17:17] } <= { N235 };
    end 
    if(N348) begin
      { v_r[16:16] } <= { N235 };
    end 
    if(N349) begin
      { v_r[15:15] } <= { N235 };
    end 
    if(N350) begin
      { v_r[14:14] } <= { N235 };
    end 
    if(N351) begin
      { v_r[13:13] } <= { N235 };
    end 
    if(N352) begin
      { v_r[12:12] } <= { N235 };
    end 
    if(N353) begin
      { v_r[11:11] } <= { N235 };
    end 
    if(N354) begin
      { v_r[10:10] } <= { N235 };
    end 
    if(N355) begin
      { v_r[9:9] } <= { N235 };
    end 
    if(N356) begin
      { v_r[8:8] } <= { N235 };
    end 
    if(N357) begin
      { v_r[7:7] } <= { N235 };
    end 
    if(N358) begin
      { v_r[6:6] } <= { N235 };
    end 
    if(N359) begin
      { v_r[5:5] } <= { N235 };
    end 
    if(N360) begin
      { v_r[4:4] } <= { N235 };
    end 
    if(N361) begin
      { v_r[3:3] } <= { N235 };
    end 
    if(N362) begin
      { v_r[2:2] } <= { N235 };
    end 
    if(N363) begin
      { v_r[1:1] } <= { N235 };
    end 
    if(N364) begin
      { v_r[0:0] } <= { N235 };
    end 
  end


endmodule



module instr_scan_vaddr_width_p39_instr_width_p32
(
  instr_i,
  scan_o
);

  input [31:0] instr_i;
  output [68:0] scan_o;
  wire [68:0] scan_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,
  N23,N24,N25,N26,N27,N28,N29,N30;
  assign scan_o[66] = 1'b0;
  assign scan_o[67] = 1'b0;
  assign N7 = instr_i[0] & instr_i[1];
  assign scan_o[68] = ~N7;
  assign N9 = ~instr_i[6];
  assign N10 = ~instr_i[5];
  assign N11 = ~instr_i[3];
  assign N12 = ~instr_i[2];
  assign N13 = ~instr_i[1];
  assign N14 = ~instr_i[0];
  assign N15 = N10 | N9;
  assign N16 = instr_i[4] | N15;
  assign N17 = N11 | N16;
  assign N18 = N12 | N17;
  assign N19 = N13 | N18;
  assign N20 = N14 | N19;
  assign N21 = ~N20;
  assign N22 = instr_i[3] | N16;
  assign N23 = N12 | N22;
  assign N24 = N13 | N23;
  assign N25 = N14 | N24;
  assign N26 = ~N25;
  assign N27 = instr_i[2] | N22;
  assign N28 = N13 | N27;
  assign N29 = N14 | N28;
  assign N30 = ~N29;
  assign scan_o[65:64] = (N0)? { 1'b0, 1'b0 } : 
                         (N1)? { 1'b0, 1'b1 } : 
                         (N4)? { 1'b1, N20 } : 1'b0;
  assign N0 = N30;
  assign N1 = N26;
  assign scan_o[63:0] = (N0)? { instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[7:7], instr_i[30:25], instr_i[11:8], 1'b0 } : 
                        (N1)? { instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:20] } : 
                        (N2)? { instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[19:12], instr_i[20:20], instr_i[30:21], 1'b0 } : 
                        (N6)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N2 = N21;
  assign N3 = N26 | N30;
  assign N4 = ~N3;
  assign N5 = N21 | N3;
  assign N6 = ~N5;

endmodule



module bp_fe_pc_gen_02
(
  clk_i,
  reset_i,
  pc_gen_icache_o,
  pc_gen_icache_v_o,
  pc_gen_icache_ready_i,
  icache_pc_gen_i,
  icache_pc_gen_v_i,
  icache_pc_gen_ready_o,
  icache_miss_i,
  instr_access_fault_i,
  pc_gen_itlb_o,
  pc_gen_itlb_v_o,
  pc_gen_itlb_ready_i,
  pc_gen_fe_o,
  pc_gen_fe_v_o,
  pc_gen_fe_ready_i,
  fe_pc_gen_i,
  fe_pc_gen_v_i,
  fe_pc_gen_ready_o,
  itlb_miss_i
);

  output [38:0] pc_gen_icache_o;
  input [70:0] icache_pc_gen_i;
  output [38:0] pc_gen_itlb_o;
  output [168:0] pc_gen_fe_o;
  input [71:0] fe_pc_gen_i;
  input clk_i;
  input reset_i;
  input pc_gen_icache_ready_i;
  input icache_pc_gen_v_i;
  input icache_miss_i;
  input instr_access_fault_i;
  input pc_gen_itlb_ready_i;
  input pc_gen_fe_ready_i;
  input fe_pc_gen_v_i;
  input itlb_miss_i;
  output pc_gen_icache_v_o;
  output icache_pc_gen_ready_o;
  output pc_gen_itlb_v_o;
  output pc_gen_fe_v_o;
  output fe_pc_gen_ready_o;
  wire [38:0] pc_gen_icache_o,pc_gen_itlb_o,pc_resume_n,btb_br_tgt_lo,br_target;
  wire [168:0] pc_gen_fe_o;
  wire pc_gen_icache_v_o,icache_pc_gen_ready_o,pc_gen_itlb_v_o,pc_gen_fe_v_o,
  fe_pc_gen_ready_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,fe_pc_gen_v_i,state_reset_v,pc_redirect_v,
  icache_fence_v,itlb_fence_v,cmd_nonattaboy_v,misalign_exception,
  itlb_miss_exception,instr_access_fault_exception,fetch_fail,queue_miss,flush,fe_instr_v,
  fe_exception_v,N9,N10,N11,N12,N13,N14,N15,N16,pc_v_if1_n,N17,N18,N19,N20,N21,N22,N23,N24,
  N25,N26,N27,N28,N29,N30,btb_br_tgt_v_lo,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,
  N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,
  N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,
  N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,
  N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,
  N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,
  pc_v_if2_n,n_2_net_,scan_instr_is_compressed_,scan_instr_instr_scan_class__3_,
  scan_instr_instr_scan_class__2_,scan_instr_instr_scan_class__1_,
  scan_instr_instr_scan_class__0_,scan_instr_imm__63_,scan_instr_imm__62_,scan_instr_imm__61_,
  scan_instr_imm__60_,scan_instr_imm__59_,scan_instr_imm__58_,scan_instr_imm__57_,
  scan_instr_imm__56_,scan_instr_imm__55_,scan_instr_imm__54_,scan_instr_imm__53_,
  scan_instr_imm__52_,scan_instr_imm__51_,scan_instr_imm__50_,scan_instr_imm__49_,
  scan_instr_imm__48_,scan_instr_imm__47_,scan_instr_imm__46_,scan_instr_imm__45_,
  scan_instr_imm__44_,scan_instr_imm__43_,scan_instr_imm__42_,scan_instr_imm__41_,
  scan_instr_imm__40_,scan_instr_imm__39_,scan_instr_imm__38_,scan_instr_imm__37_,
  scan_instr_imm__36_,scan_instr_imm__35_,scan_instr_imm__34_,scan_instr_imm__33_,
  scan_instr_imm__32_,scan_instr_imm__31_,scan_instr_imm__30_,scan_instr_imm__29_,
  scan_instr_imm__28_,scan_instr_imm__27_,scan_instr_imm__26_,scan_instr_imm__25_,
  scan_instr_imm__24_,scan_instr_imm__23_,scan_instr_imm__22_,scan_instr_imm__21_,
  scan_instr_imm__20_,scan_instr_imm__19_,scan_instr_imm__18_,scan_instr_imm__17_,
  scan_instr_imm__16_,scan_instr_imm__15_,scan_instr_imm__14_,scan_instr_imm__13_,
  scan_instr_imm__12_,scan_instr_imm__11_,scan_instr_imm__10_,scan_instr_imm__9_,
  scan_instr_imm__8_,scan_instr_imm__7_,scan_instr_imm__6_,scan_instr_imm__5_,
  scan_instr_imm__4_,scan_instr_imm__3_,scan_instr_imm__2_,scan_instr_imm__1_,scan_instr_imm__0_,
  N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,
  N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159;
  wire [1:0] state_n;
  wire [26:0] fe_queue_branch_metadata_r;
  reg [38:0] pc_resume_r,pc_if2_r,pc_if1_r;
  reg [1:0] state_r;
  reg itlb_miss_if2_r,pc_v_if1_r,pc_v_if2_r;
  assign icache_pc_gen_ready_o = 1'b1;
  assign pc_gen_fe_o[0] = 1'b0;
  assign pc_gen_fe_o[99] = 1'b0;
  assign pc_gen_fe_o[100] = 1'b0;
  assign pc_gen_fe_o[101] = 1'b0;
  assign pc_gen_fe_o[102] = 1'b0;
  assign pc_gen_fe_o[103] = 1'b0;
  assign pc_gen_fe_o[104] = 1'b0;
  assign pc_gen_fe_o[105] = 1'b0;
  assign pc_gen_fe_o[106] = 1'b0;
  assign pc_gen_fe_o[107] = 1'b0;
  assign pc_gen_fe_o[108] = 1'b0;
  assign pc_gen_fe_o[109] = 1'b0;
  assign pc_gen_fe_o[110] = 1'b0;
  assign pc_gen_fe_o[111] = 1'b0;
  assign pc_gen_fe_o[112] = 1'b0;
  assign pc_gen_fe_o[113] = 1'b0;
  assign pc_gen_fe_o[114] = 1'b0;
  assign pc_gen_fe_o[115] = 1'b0;
  assign pc_gen_fe_o[116] = 1'b0;
  assign pc_gen_fe_o[117] = 1'b0;
  assign pc_gen_fe_o[118] = 1'b0;
  assign pc_gen_fe_o[119] = 1'b0;
  assign pc_gen_fe_o[120] = 1'b0;
  assign pc_gen_fe_o[121] = 1'b0;
  assign pc_gen_fe_o[122] = 1'b0;
  assign pc_gen_fe_o[123] = 1'b0;
  assign pc_gen_fe_o[124] = 1'b0;
  assign pc_gen_fe_o[125] = 1'b0;
  assign pc_gen_fe_o[126] = 1'b0;
  assign pc_gen_fe_o[127] = 1'b0;
  assign pc_gen_fe_o[128] = 1'b0;
  assign pc_gen_fe_o[129] = 1'b0;
  assign pc_gen_fe_o[130] = 1'b0;
  assign pc_gen_fe_o[131] = 1'b0;
  assign pc_gen_fe_o[132] = 1'b0;
  assign pc_gen_fe_o[133] = 1'b0;
  assign pc_gen_fe_o[134] = 1'b0;
  assign pc_gen_fe_o[135] = 1'b0;
  assign pc_gen_fe_o[136] = 1'b0;
  assign pc_gen_fe_o[137] = 1'b0;
  assign pc_gen_fe_o[138] = 1'b0;
  assign pc_gen_fe_o[139] = 1'b0;
  assign pc_gen_fe_o[140] = 1'b0;
  assign pc_gen_fe_o[141] = 1'b0;
  assign pc_gen_fe_o[142] = 1'b0;
  assign pc_gen_fe_o[143] = 1'b0;
  assign pc_gen_fe_o[144] = 1'b0;
  assign pc_gen_fe_o[145] = 1'b0;
  assign pc_gen_fe_o[146] = 1'b0;
  assign pc_gen_fe_o[147] = 1'b0;
  assign pc_gen_fe_o[148] = 1'b0;
  assign pc_gen_fe_o[149] = 1'b0;
  assign pc_gen_fe_o[150] = 1'b0;
  assign pc_gen_fe_o[151] = 1'b0;
  assign pc_gen_fe_o[152] = 1'b0;
  assign pc_gen_fe_o[153] = 1'b0;
  assign pc_gen_fe_o[154] = 1'b0;
  assign pc_gen_fe_o[155] = 1'b0;
  assign pc_gen_fe_o[156] = 1'b0;
  assign pc_gen_fe_o[157] = 1'b0;
  assign pc_gen_fe_o[158] = 1'b0;
  assign pc_gen_fe_o[159] = 1'b0;
  assign pc_gen_fe_o[160] = 1'b0;
  assign pc_gen_fe_o[161] = 1'b0;
  assign pc_gen_fe_o[162] = 1'b0;
  assign pc_gen_fe_o[163] = 1'b0;
  assign pc_gen_fe_o[164] = 1'b0;
  assign pc_gen_fe_o[165] = 1'b0;
  assign pc_gen_fe_o[166] = 1'b0;
  assign pc_gen_fe_o[167] = 1'b0;
  assign pc_gen_itlb_o[38] = pc_gen_icache_o[38];
  assign pc_gen_itlb_o[37] = pc_gen_icache_o[37];
  assign pc_gen_itlb_o[36] = pc_gen_icache_o[36];
  assign pc_gen_itlb_o[35] = pc_gen_icache_o[35];
  assign pc_gen_itlb_o[34] = pc_gen_icache_o[34];
  assign pc_gen_itlb_o[33] = pc_gen_icache_o[33];
  assign pc_gen_itlb_o[32] = pc_gen_icache_o[32];
  assign pc_gen_itlb_o[31] = pc_gen_icache_o[31];
  assign pc_gen_itlb_o[30] = pc_gen_icache_o[30];
  assign pc_gen_itlb_o[29] = pc_gen_icache_o[29];
  assign pc_gen_itlb_o[28] = pc_gen_icache_o[28];
  assign pc_gen_itlb_o[27] = pc_gen_icache_o[27];
  assign pc_gen_itlb_o[26] = pc_gen_icache_o[26];
  assign pc_gen_itlb_o[25] = pc_gen_icache_o[25];
  assign pc_gen_itlb_o[24] = pc_gen_icache_o[24];
  assign pc_gen_itlb_o[23] = pc_gen_icache_o[23];
  assign pc_gen_itlb_o[22] = pc_gen_icache_o[22];
  assign pc_gen_itlb_o[21] = pc_gen_icache_o[21];
  assign pc_gen_itlb_o[20] = pc_gen_icache_o[20];
  assign pc_gen_itlb_o[19] = pc_gen_icache_o[19];
  assign pc_gen_itlb_o[18] = pc_gen_icache_o[18];
  assign pc_gen_itlb_o[17] = pc_gen_icache_o[17];
  assign pc_gen_itlb_o[16] = pc_gen_icache_o[16];
  assign pc_gen_itlb_o[15] = pc_gen_icache_o[15];
  assign pc_gen_itlb_o[14] = pc_gen_icache_o[14];
  assign pc_gen_itlb_o[13] = pc_gen_icache_o[13];
  assign pc_gen_itlb_o[12] = pc_gen_icache_o[12];
  assign pc_gen_itlb_o[11] = pc_gen_icache_o[11];
  assign pc_gen_itlb_o[10] = pc_gen_icache_o[10];
  assign pc_gen_itlb_o[9] = pc_gen_icache_o[9];
  assign pc_gen_itlb_o[8] = pc_gen_icache_o[8];
  assign pc_gen_itlb_o[7] = pc_gen_icache_o[7];
  assign pc_gen_itlb_o[6] = pc_gen_icache_o[6];
  assign pc_gen_itlb_o[5] = pc_gen_icache_o[5];
  assign pc_gen_itlb_o[4] = pc_gen_icache_o[4];
  assign pc_gen_itlb_o[3] = pc_gen_icache_o[3];
  assign pc_gen_itlb_o[2] = pc_gen_icache_o[2];
  assign pc_gen_itlb_o[1] = pc_gen_icache_o[1];
  assign pc_gen_itlb_o[0] = pc_gen_icache_o[0];
  assign fe_pc_gen_ready_o = fe_pc_gen_v_i;
  assign N11 = N10 & N142;
  assign N12 = N10 | state_r[0];
  assign N14 = state_r[1] | N142;
  assign N16 = state_r[1] & state_r[0];

  bsg_dff_reset_en_width_p27
  branch_metadata_fwd_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(pc_gen_fe_v_o),
    .data_i({ icache_pc_gen_i[17:2], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }),
    .data_o(fe_queue_branch_metadata_r)
  );


  bp_fe_btb_vaddr_width_p39_btb_tag_width_p10_btb_idx_width_p6
  btb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .r_addr_i(pc_gen_icache_o),
    .r_v_i(pc_v_if1_n),
    .br_tgt_o(btb_br_tgt_lo),
    .br_tgt_v_o(btb_br_tgt_v_lo),
    .w_tag_i(fe_pc_gen_i[32:23]),
    .w_idx_i(fe_pc_gen_i[22:17]),
    .w_v_i(n_2_net_),
    .br_tgt_i(fe_pc_gen_i[71:33])
  );


  instr_scan_vaddr_width_p39_instr_width_p32
  instr_scan_1
  (
    .instr_i(icache_pc_gen_i[70:39]),
    .scan_o({ scan_instr_is_compressed_, scan_instr_instr_scan_class__3_, scan_instr_instr_scan_class__2_, scan_instr_instr_scan_class__1_, scan_instr_instr_scan_class__0_, scan_instr_imm__63_, scan_instr_imm__62_, scan_instr_imm__61_, scan_instr_imm__60_, scan_instr_imm__59_, scan_instr_imm__58_, scan_instr_imm__57_, scan_instr_imm__56_, scan_instr_imm__55_, scan_instr_imm__54_, scan_instr_imm__53_, scan_instr_imm__52_, scan_instr_imm__51_, scan_instr_imm__50_, scan_instr_imm__49_, scan_instr_imm__48_, scan_instr_imm__47_, scan_instr_imm__46_, scan_instr_imm__45_, scan_instr_imm__44_, scan_instr_imm__43_, scan_instr_imm__42_, scan_instr_imm__41_, scan_instr_imm__40_, scan_instr_imm__39_, scan_instr_imm__38_, scan_instr_imm__37_, scan_instr_imm__36_, scan_instr_imm__35_, scan_instr_imm__34_, scan_instr_imm__33_, scan_instr_imm__32_, scan_instr_imm__31_, scan_instr_imm__30_, scan_instr_imm__29_, scan_instr_imm__28_, scan_instr_imm__27_, scan_instr_imm__26_, scan_instr_imm__25_, scan_instr_imm__24_, scan_instr_imm__23_, scan_instr_imm__22_, scan_instr_imm__21_, scan_instr_imm__20_, scan_instr_imm__19_, scan_instr_imm__18_, scan_instr_imm__17_, scan_instr_imm__16_, scan_instr_imm__15_, scan_instr_imm__14_, scan_instr_imm__13_, scan_instr_imm__12_, scan_instr_imm__11_, scan_instr_imm__10_, scan_instr_imm__9_, scan_instr_imm__8_, scan_instr_imm__7_, scan_instr_imm__6_, scan_instr_imm__5_, scan_instr_imm__4_, scan_instr_imm__3_, scan_instr_imm__2_, scan_instr_imm__1_, scan_instr_imm__0_ })
  );

  assign N139 = ~state_n[0];
  assign N140 = N139 | state_n[1];
  assign N141 = ~N140;
  assign N142 = ~state_r[0];
  assign N143 = N142 | state_r[1];
  assign N144 = ~N143;
  assign N145 = state_r[0] | state_r[1];
  assign N146 = N142 | state_r[1];
  assign N147 = pc_if2_r[0] | pc_if2_r[1];
  assign br_target = icache_pc_gen_i[38:0] + icache_pc_gen_i[70:59];
  assign { N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79 } = pc_if1_r + { 1'b1, 1'b0, 1'b0 };
  assign { N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40 } = pc_if2_r + { 1'b1, 1'b0, 1'b0 };
  assign pc_resume_n = (N0)? fe_pc_gen_i[71:33] : 
                       (N25)? pc_if2_r : 1'b0;
  assign N0 = cmd_nonattaboy_v;
  assign { N23, N22 } = (N0)? { 1'b0, 1'b1 } : 
                        (N26)? { 1'b1, 1'b0 } : 
                        (N29)? { 1'b0, 1'b0 } : 
                        (N21)? { 1'b0, 1'b1 } : 1'b0;
  assign state_n = (N1)? { cmd_nonattaboy_v, 1'b0 } : 
                   (N2)? { N17, N18 } : 
                   (N3)? { N23, N22 } : 
                   (N4)? { 1'b0, 1'b0 } : 1'b0;
  assign N1 = N11;
  assign N2 = N13;
  assign N3 = N15;
  assign N4 = N16;
  assign pc_gen_icache_o = (N5)? fe_pc_gen_i[71:33] : 
                           (N119)? fe_pc_gen_i[71:33] : 
                           (N122)? pc_resume_r : 
                           (N125)? btb_br_tgt_lo : 
                           (N128)? br_target : 
                           (N131)? { N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40 } : 
                           (N38)? { N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79 } : 1'b0;
  assign N5 = state_reset_v;
  assign { N136, N135 } = (N6)? { 1'b0, 1'b0 } : 
                          (N138)? { 1'b0, 1'b1 } : 
                          (N134)? { 1'b1, 1'b1 } : 1'b0;
  assign N6 = misalign_exception;
  assign pc_gen_fe_o[98:1] = (N7)? { pc_if2_r, N136, N135, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                             (N8)? { icache_pc_gen_i[38:0], icache_pc_gen_i[70:39], fe_queue_branch_metadata_r } : 1'b0;
  assign N7 = pc_gen_fe_o[168];
  assign N8 = N132;
  assign state_reset_v = fe_pc_gen_v_i & fe_pc_gen_i[5];
  assign pc_redirect_v = fe_pc_gen_v_i & fe_pc_gen_i[4];
  assign icache_fence_v = fe_pc_gen_v_i & fe_pc_gen_i[1];
  assign itlb_fence_v = fe_pc_gen_v_i & fe_pc_gen_i[0];
  assign cmd_nonattaboy_v = fe_pc_gen_v_i & N148;
  assign N148 = ~fe_pc_gen_i[3];
  assign misalign_exception = pc_v_if2_r & N147;
  assign itlb_miss_exception = pc_v_if2_r & itlb_miss_if2_r;
  assign instr_access_fault_exception = pc_v_if2_r & instr_access_fault_i;
  assign fetch_fail = pc_v_if2_r & N149;
  assign N149 = ~pc_gen_fe_v_o;
  assign queue_miss = pc_v_if2_r & N150;
  assign N150 = ~pc_gen_fe_ready_i;
  assign flush = N152 | cmd_nonattaboy_v;
  assign N152 = N151 | queue_miss;
  assign N151 = itlb_miss_if2_r | icache_miss_i;
  assign fe_instr_v = pc_v_if2_r & N153;
  assign N153 = ~flush;
  assign fe_exception_v = pc_v_if2_r & N155;
  assign N155 = N154 | itlb_miss_exception;
  assign N154 = instr_access_fault_exception | misalign_exception;
  assign N9 = N144 | cmd_nonattaboy_v;
  assign N10 = ~state_r[1];
  assign N13 = ~N12;
  assign N15 = ~N14;
  assign N17 = ~pc_v_if1_n;
  assign N18 = pc_v_if1_n;
  assign N19 = fetch_fail | cmd_nonattaboy_v;
  assign N20 = fe_exception_v | N19;
  assign N21 = ~N20;
  assign N24 = ~cmd_nonattaboy_v;
  assign N25 = N144 & N24;
  assign N26 = fetch_fail & N24;
  assign N27 = ~fetch_fail;
  assign N28 = N24 & N27;
  assign N29 = fe_exception_v & N28;
  assign N30 = N156 | itlb_fence_v;
  assign N156 = pc_redirect_v | icache_fence_v;
  assign N31 = 1'b0;
  assign N32 = 1'b0;
  assign N33 = N30 | state_reset_v;
  assign N34 = N146 | N33;
  assign N35 = btb_br_tgt_v_lo | N34;
  assign N36 = N31 | N35;
  assign N37 = N32 | N36;
  assign N38 = ~N37;
  assign N39 = N131;
  assign N118 = ~state_reset_v;
  assign N119 = N30 & N118;
  assign N120 = ~N30;
  assign N121 = N118 & N120;
  assign N122 = N146 & N121;
  assign N123 = ~N146;
  assign N124 = N121 & N123;
  assign N125 = btb_br_tgt_v_lo & N124;
  assign N126 = ~btb_br_tgt_v_lo;
  assign N127 = N124 & N126;
  assign N128 = N31 & N127;
  assign N129 = ~N31;
  assign N130 = N127 & N129;
  assign N131 = N32 & N130;
  assign pc_v_if1_n = N158 & pc_gen_icache_ready_i;
  assign N158 = N157 & pc_gen_fe_ready_i;
  assign N157 = N145 & pc_gen_itlb_ready_i;
  assign pc_v_if2_n = pc_v_if1_r & N153;
  assign n_2_net_ = pc_redirect_v & fe_pc_gen_v_i;
  assign N132 = ~fe_exception_v;
  assign pc_gen_fe_o[168] = fe_exception_v;
  assign N133 = itlb_miss_exception | misalign_exception;
  assign N134 = ~N133;
  assign N137 = ~misalign_exception;
  assign N138 = itlb_miss_exception & N137;
  assign pc_gen_fe_v_o = pc_gen_fe_ready_i & N159;
  assign N159 = fe_instr_v | fe_exception_v;
  assign pc_gen_icache_v_o = pc_gen_icache_ready_i & pc_v_if1_n;
  assign pc_gen_itlb_v_o = pc_gen_itlb_ready_i & pc_v_if1_n;

  always @(posedge clk_i) begin
    if(N9) begin
      { pc_resume_r[38:0] } <= { pc_resume_n[38:0] };
    end 
    if(reset_i) begin
      { state_r[1:0] } <= { 1'b0, 1'b0 };
      itlb_miss_if2_r <= 1'b0;
      pc_v_if1_r <= 1'b0;
      pc_v_if2_r <= 1'b0;
    end else if(1'b1) begin
      { state_r[1:0] } <= { state_n[1:0] };
      itlb_miss_if2_r <= itlb_miss_i;
      pc_v_if1_r <= pc_v_if1_n;
      pc_v_if2_r <= pc_v_if2_n;
    end 
    if(reset_i) begin
      { pc_if2_r[38:0] } <= { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 };
      { pc_if1_r[38:0] } <= { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 };
    end else if(N141) begin
      { pc_if2_r[38:0] } <= { pc_if1_r[38:0] };
      { pc_if1_r[38:0] } <= { pc_gen_icache_o[38:0] };
    end 
  end


endmodule



module bsg_mem_1rw_sync_mask_write_bit_width_p232_els_p64
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_mask_i,
  w_i,
  data_o
);

  input [231:0] data_i;
  input [5:0] addr_i;
  input [231:0] w_mask_i;
  output [231:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [231:0] data_o;

  nangate45_120x64_1P_bit
  macro_mem0
  (
    .clk(clk_i),
    .we_in(w_i),
    .ce_in(v_i),
    .addr_in(addr_i),
    .wd_in(data_i[115:0]),
    .rd_out(data_o[115:0]),
    .w_mask_in(w_mask_i[115:0])
  );



  nangate45_120x64_1P_bit
  macro_mem1
  (
    .clk(clk_i),
    .we_in(w_i),
    .ce_in(v_i),
    .addr_in(addr_i),
    .wd_in(data_i[231:116]),
    .rd_out(data_o[231:116]),
    .w_mask_in(w_mask_i[231:116])
  );


endmodule



module bsg_mem_1rw_sync_mask_write_byte_els_p512_data_width_p64
(
  clk_i,
  reset_i,
  v_i,
  w_i,
  addr_i,
  data_i,
  write_mask_i,
  data_o
);

  input [8:0] addr_i;
  input [63:0] data_i;
  input [7:0] write_mask_i;
  output [63:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [63:0] data_o;

  nangate45_64x512_1P_BM
  macro_mem
  (
    .clk(clk_i),
    .we_in(w_i),
    .ce_in(v_i),
    .addr_in(addr_i),
    .wd_in(data_i),
    .rd_out(data_o),
    .w_mask_in(w_mask_i)
  );


endmodule



module bsg_scan_width_p8_or_p1_lo_to_hi_p1
(
  i,
  o
);

  input [7:0] i;
  output [7:0] o;
  wire [7:0] o;
  wire t_2__7_,t_2__6_,t_2__5_,t_2__4_,t_2__3_,t_2__2_,t_2__1_,t_2__0_,t_1__7_,t_1__6_,
  t_1__5_,t_1__4_,t_1__3_,t_1__2_,t_1__1_,t_1__0_;
  assign t_1__7_ = i[0] | 1'b0;
  assign t_1__6_ = i[1] | i[0];
  assign t_1__5_ = i[2] | i[1];
  assign t_1__4_ = i[3] | i[2];
  assign t_1__3_ = i[4] | i[3];
  assign t_1__2_ = i[5] | i[4];
  assign t_1__1_ = i[6] | i[5];
  assign t_1__0_ = i[7] | i[6];
  assign t_2__7_ = t_1__7_ | 1'b0;
  assign t_2__6_ = t_1__6_ | 1'b0;
  assign t_2__5_ = t_1__5_ | t_1__7_;
  assign t_2__4_ = t_1__4_ | t_1__6_;
  assign t_2__3_ = t_1__3_ | t_1__5_;
  assign t_2__2_ = t_1__2_ | t_1__4_;
  assign t_2__1_ = t_1__1_ | t_1__3_;
  assign t_2__0_ = t_1__0_ | t_1__2_;
  assign o[0] = t_2__7_ | 1'b0;
  assign o[1] = t_2__6_ | 1'b0;
  assign o[2] = t_2__5_ | 1'b0;
  assign o[3] = t_2__4_ | 1'b0;
  assign o[4] = t_2__3_ | t_2__7_;
  assign o[5] = t_2__2_ | t_2__6_;
  assign o[6] = t_2__1_ | t_2__5_;
  assign o[7] = t_2__0_ | t_2__4_;

endmodule



module bsg_priority_encode_one_hot_out_width_p8_lo_to_hi_p1
(
  i,
  o
);

  input [7:0] i;
  output [7:0] o;
  wire [7:0] o;
  wire N0,N1,N2,N3,N4,N5,N6;
  wire [7:1] scan_lo;

  bsg_scan_width_p8_or_p1_lo_to_hi_p1
  genblk1_scan
  (
    .i(i),
    .o({ scan_lo, o[0:0] })
  );

  assign o[7] = scan_lo[7] & N0;
  assign N0 = ~scan_lo[6];
  assign o[6] = scan_lo[6] & N1;
  assign N1 = ~scan_lo[5];
  assign o[5] = scan_lo[5] & N2;
  assign N2 = ~scan_lo[4];
  assign o[4] = scan_lo[4] & N3;
  assign N3 = ~scan_lo[3];
  assign o[3] = scan_lo[3] & N4;
  assign N4 = ~scan_lo[2];
  assign o[2] = scan_lo[2] & N5;
  assign N5 = ~scan_lo[1];
  assign o[1] = scan_lo[1] & N6;
  assign N6 = ~o[0];

endmodule



module bsg_encode_one_hot_width_p1
(
  i,
  addr_o,
  v_o
);

  input [0:0] i;
  output [0:0] addr_o;
  output v_o;
  wire [0:0] addr_o;
  wire v_o;
  assign v_o = i[0];
  assign addr_o[0] = 1'b0;

endmodule



module bsg_encode_one_hot_width_p2
(
  i,
  addr_o,
  v_o
);

  input [1:0] i;
  output [0:0] addr_o;
  output v_o;
  wire [0:0] addr_o,aligned_vs;
  wire v_o;
  wire [1:0] aligned_addrs;

  bsg_encode_one_hot_width_p1
  aligned_left
  (
    .i(i[0]),
    .addr_o(aligned_addrs[0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p1
  aligned_right
  (
    .i(i[1]),
    .addr_o(aligned_addrs[1]),
    .v_o(addr_o[0])
  );

  assign v_o = addr_o[0] | aligned_vs[0];

endmodule



module bsg_encode_one_hot_width_p4
(
  i,
  addr_o,
  v_o
);

  input [3:0] i;
  output [1:0] addr_o;
  output v_o;
  wire [1:0] addr_o,aligned_addrs;
  wire v_o;
  wire [0:0] aligned_vs;

  bsg_encode_one_hot_width_p2
  aligned_left
  (
    .i(i[1:0]),
    .addr_o(aligned_addrs[0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p2
  aligned_right
  (
    .i(i[3:2]),
    .addr_o(aligned_addrs[1]),
    .v_o(addr_o[1])
  );

  assign v_o = addr_o[1] | aligned_vs[0];
  assign addr_o[0] = aligned_addrs[0] | aligned_addrs[1];

endmodule



module bsg_encode_one_hot_width_p8_lo_to_hi_p1
(
  i,
  addr_o,
  v_o
);

  input [7:0] i;
  output [2:0] addr_o;
  output v_o;
  wire [2:0] addr_o;
  wire v_o;
  wire [3:0] aligned_addrs;
  wire [0:0] aligned_vs;

  bsg_encode_one_hot_width_p4
  aligned_left
  (
    .i(i[3:0]),
    .addr_o(aligned_addrs[1:0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p4
  aligned_right
  (
    .i(i[7:4]),
    .addr_o(aligned_addrs[3:2]),
    .v_o(addr_o[2])
  );

  assign v_o = addr_o[2] | aligned_vs[0];
  assign addr_o[1] = aligned_addrs[1] | aligned_addrs[3];
  assign addr_o[0] = aligned_addrs[0] | aligned_addrs[2];

endmodule



module bsg_priority_encode_width_p8_lo_to_hi_p1
(
  i,
  addr_o,
  v_o
);

  input [7:0] i;
  output [2:0] addr_o;
  output v_o;
  wire [2:0] addr_o;
  wire v_o;
  wire [7:0] enc_lo;

  bsg_priority_encode_one_hot_out_width_p8_lo_to_hi_p1
  a
  (
    .i(i),
    .o(enc_lo)
  );


  bsg_encode_one_hot_width_p8_lo_to_hi_p1
  b
  (
    .i(enc_lo),
    .addr_o(addr_o),
    .v_o(v_o)
  );


endmodule



module bsg_mem_1rw_sync_mask_write_bit_width_p7_els_p64
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_mask_i,
  w_i,
  data_o
);

  input [6:0] data_i;
  input [5:0] addr_i;
  input [6:0] w_mask_i;
  output [6:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [6:0] data_o;

  nangate45_8x64_1P_bit
  macro_mem
  (
    .clk(clk_i),
    .we_in(w_i),
    .ce_in(v_i),
    .addr_in(addr_i),
    .wd_in(data_i[6:0]),
    .rd_out(data_o[6:0]),
    .w_mask_in(w_mask_i[6:0])
  );


endmodule



module bsg_scan_7_1_1
(
  i,
  o
);

  input [6:0] i;
  output [6:0] o;
  wire [6:0] o;
  wire t_2__6_,t_2__5_,t_2__4_,t_2__3_,t_2__2_,t_2__1_,t_2__0_,t_1__6_,t_1__5_,t_1__4_,
  t_1__3_,t_1__2_,t_1__1_,t_1__0_;
  assign t_1__6_ = i[0] | 1'b0;
  assign t_1__5_ = i[1] | i[0];
  assign t_1__4_ = i[2] | i[1];
  assign t_1__3_ = i[3] | i[2];
  assign t_1__2_ = i[4] | i[3];
  assign t_1__1_ = i[5] | i[4];
  assign t_1__0_ = i[6] | i[5];
  assign t_2__6_ = t_1__6_ | 1'b0;
  assign t_2__5_ = t_1__5_ | 1'b0;
  assign t_2__4_ = t_1__4_ | t_1__6_;
  assign t_2__3_ = t_1__3_ | t_1__5_;
  assign t_2__2_ = t_1__2_ | t_1__4_;
  assign t_2__1_ = t_1__1_ | t_1__3_;
  assign t_2__0_ = t_1__0_ | t_1__2_;
  assign o[0] = t_2__6_ | 1'b0;
  assign o[1] = t_2__5_ | 1'b0;
  assign o[2] = t_2__4_ | 1'b0;
  assign o[3] = t_2__3_ | 1'b0;
  assign o[4] = t_2__2_ | t_2__6_;
  assign o[5] = t_2__1_ | t_2__5_;
  assign o[6] = t_2__0_ | t_2__4_;

endmodule



module bsg_priority_encode_one_hot_out_7_1
(
  i,
  o
);

  input [6:0] i;
  output [6:0] o;
  wire [6:0] o;
  wire N0,N1,N2,N3,N4,N5;
  wire [6:1] scan_lo;

  bsg_scan_7_1_1
  genblk1_scan
  (
    .i(i),
    .o({ scan_lo, o[0:0] })
  );

  assign o[6] = scan_lo[6] & N0;
  assign N0 = ~scan_lo[5];
  assign o[5] = scan_lo[5] & N1;
  assign N1 = ~scan_lo[4];
  assign o[4] = scan_lo[4] & N2;
  assign N2 = ~scan_lo[3];
  assign o[3] = scan_lo[3] & N3;
  assign N3 = ~scan_lo[2];
  assign o[2] = scan_lo[2] & N4;
  assign N4 = ~scan_lo[1];
  assign o[1] = scan_lo[1] & N5;
  assign N5 = ~o[0];

endmodule



module bsg_encode_one_hot_width_p8
(
  i,
  addr_o,
  v_o
);

  input [7:0] i;
  output [2:0] addr_o;
  output v_o;
  wire [2:0] addr_o;
  wire v_o;
  wire [3:0] aligned_addrs;
  wire [0:0] aligned_vs;

  bsg_encode_one_hot_width_p4
  aligned_left
  (
    .i(i[3:0]),
    .addr_o(aligned_addrs[1:0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p4
  aligned_right
  (
    .i(i[7:4]),
    .addr_o(aligned_addrs[3:2]),
    .v_o(addr_o[2])
  );

  assign v_o = addr_o[2] | aligned_vs[0];
  assign addr_o[1] = aligned_addrs[1] | aligned_addrs[3];
  assign addr_o[0] = aligned_addrs[0] | aligned_addrs[2];

endmodule



module bsg_encode_one_hot_7_1
(
  i,
  addr_o,
  v_o
);

  input [6:0] i;
  output [2:0] addr_o;
  output v_o;
  wire [2:0] addr_o;
  wire v_o;

  bsg_encode_one_hot_width_p8
  unaligned_align
  (
    .i({ 1'b0, i }),
    .addr_o(addr_o),
    .v_o(v_o)
  );


endmodule



module bsg_priority_encode_7_1
(
  i,
  addr_o,
  v_o
);

  input [6:0] i;
  output [2:0] addr_o;
  output v_o;
  wire [2:0] addr_o;
  wire v_o;
  wire [6:0] enc_lo;

  bsg_priority_encode_one_hot_out_7_1
  a
  (
    .i(i),
    .o(enc_lo)
  );


  bsg_encode_one_hot_7_1
  b
  (
    .i(enc_lo),
    .addr_o(addr_o),
    .v_o(v_o)
  );


endmodule



module bsg_lru_pseudo_tree_encode_ways_p8
(
  lru_i,
  way_id_o
);

  input [6:0] lru_i;
  output [2:0] way_id_o;
  wire [2:0] way_id_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,pe_o_2__2_,pe_o_2__1_,pe_o_2__0_,
  pe_o_1__2_,pe_o_1__1_,pe_o_1__0_,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,
  pe_i_2__6_,pe_i_2__5_,pe_i_2__4_,pe_i_2__3_,pe_i_2__2_,pe_i_2__1_,pe_i_2__0_,pe_i_1__6_,
  pe_i_1__5_,pe_i_1__4_,pe_i_1__3_,pe_i_1__2_,pe_i_1__1_,pe_i_1__0_,N44,N45,N46,
  N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,
  N67;
  wire [6:1] mask;

  bsg_priority_encode_7_1
  rof2_1__fi3_pe
  (
    .i({ pe_i_1__6_, pe_i_1__5_, pe_i_1__4_, pe_i_1__3_, pe_i_1__2_, pe_i_1__1_, pe_i_1__0_ }),
    .addr_o({ pe_o_1__2_, pe_o_1__1_, pe_o_1__0_ })
  );

  assign { N64, N63, N62, N61, N60, N59, N58 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << { pe_o_1__2_, pe_o_1__1_, pe_o_1__0_ };

  bsg_priority_encode_7_1
  rof2_2__fi3_pe
  (
    .i({ pe_i_2__6_, pe_i_2__5_, pe_i_2__4_, pe_i_2__3_, pe_i_2__2_, pe_i_2__1_, pe_i_2__0_ }),
    .addr_o({ pe_o_2__2_, pe_o_2__1_, pe_o_2__0_ })
  );

  assign N44 = N0 & N1 & N2;
  assign N0 = ~pe_o_1__2_;
  assign N1 = ~pe_o_1__0_;
  assign N2 = ~pe_o_1__1_;
  assign N45 = pe_o_1__2_ & N3 & N4;
  assign N3 = ~pe_o_1__0_;
  assign N4 = ~pe_o_1__1_;
  assign N46 = N5 & pe_o_1__0_ & N6;
  assign N5 = ~pe_o_1__2_;
  assign N6 = ~pe_o_1__1_;
  assign N48 = N7 & N8 & pe_o_1__1_;
  assign N7 = ~pe_o_1__2_;
  assign N8 = ~pe_o_1__0_;
  assign N50 = pe_o_1__0_ & pe_o_1__1_;
  assign N47 = pe_o_1__2_ & pe_o_1__0_;
  assign N49 = pe_o_1__2_ & pe_o_1__1_;
  assign N51 = N9 & N10 & N11;
  assign N9 = ~pe_o_2__2_;
  assign N10 = ~pe_o_2__0_;
  assign N11 = ~pe_o_2__1_;
  assign N52 = pe_o_2__2_ & N12 & N13;
  assign N12 = ~pe_o_2__0_;
  assign N13 = ~pe_o_2__1_;
  assign N53 = N14 & pe_o_2__0_ & N15;
  assign N14 = ~pe_o_2__2_;
  assign N15 = ~pe_o_2__1_;
  assign N55 = N16 & N17 & pe_o_2__1_;
  assign N16 = ~pe_o_2__2_;
  assign N17 = ~pe_o_2__0_;
  assign N57 = pe_o_2__0_ & pe_o_2__1_;
  assign N54 = pe_o_2__2_ & pe_o_2__0_;
  assign N56 = pe_o_2__2_ & pe_o_2__1_;
  assign way_id_o[1] = (N18)? lru_i[0] : 
                       (N19)? lru_i[1] : 
                       (N20)? lru_i[2] : 
                       (N21)? lru_i[3] : 
                       (N22)? lru_i[4] : 
                       (N23)? lru_i[5] : 
                       (N24)? lru_i[6] : 1'b0;
  assign N18 = N44;
  assign N19 = N46;
  assign N20 = N48;
  assign N21 = N50;
  assign N22 = N45;
  assign N23 = N47;
  assign N24 = N49;
  assign way_id_o[0] = (N25)? lru_i[0] : 
                       (N26)? lru_i[1] : 
                       (N27)? lru_i[2] : 
                       (N28)? lru_i[3] : 
                       (N29)? lru_i[4] : 
                       (N30)? lru_i[5] : 
                       (N31)? lru_i[6] : 1'b0;
  assign N25 = N51;
  assign N26 = N53;
  assign N27 = N55;
  assign N28 = N57;
  assign N29 = N52;
  assign N30 = N54;
  assign N31 = N56;
  assign way_id_o[2] = (N37)? lru_i[0] : 
                       (N39)? lru_i[1] : 
                       (N41)? lru_i[2] : 
                       (N43)? lru_i[3] : 
                       (N38)? lru_i[4] : 
                       (N40)? lru_i[5] : 
                       (N42)? lru_i[6] : 1'b0;
  assign mask[1] = 1'b1 & N65;
  assign N65 = ~lru_i[0];
  assign mask[2] = 1'b1 & lru_i[0];
  assign mask[3] = mask[1] & N66;
  assign N66 = ~lru_i[1];
  assign mask[4] = mask[1] & lru_i[1];
  assign mask[5] = mask[2] & N67;
  assign N67 = ~lru_i[2];
  assign mask[6] = mask[2] & lru_i[2];
  assign N32 = N36 & N36;
  assign N33 = N36 & 1'b0;
  assign N34 = 1'b0 & N36;
  assign N35 = 1'b0 & 1'b0;
  assign N36 = ~1'b0;
  assign N37 = N32 & N36;
  assign N38 = N32 & 1'b0;
  assign N39 = N34 & N36;
  assign N40 = N34 & 1'b0;
  assign N41 = N33 & N36;
  assign N42 = N33 & 1'b0;
  assign N43 = N35 & N36;
  assign pe_i_1__6_ = mask[6] ^ 1'b0;
  assign pe_i_1__5_ = mask[5] ^ 1'b0;
  assign pe_i_1__4_ = mask[4] ^ 1'b0;
  assign pe_i_1__3_ = mask[3] ^ 1'b0;
  assign pe_i_1__2_ = mask[2] ^ 1'b0;
  assign pe_i_1__1_ = mask[1] ^ 1'b0;
  assign pe_i_1__0_ = 1'b1 ^ 1'b1;
  assign pe_i_2__6_ = pe_i_1__6_ ^ N64;
  assign pe_i_2__5_ = pe_i_1__5_ ^ N63;
  assign pe_i_2__4_ = pe_i_1__4_ ^ N62;
  assign pe_i_2__3_ = pe_i_1__3_ ^ N61;
  assign pe_i_2__2_ = pe_i_1__2_ ^ N60;
  assign pe_i_2__1_ = pe_i_1__1_ ^ N59;
  assign pe_i_2__0_ = pe_i_1__0_ ^ N58;

endmodule



module bp_fe_lce_req_02
(
  clk_i,
  reset_i,
  id_i,
  miss_i,
  miss_addr_i,
  lru_way_i,
  uncached_req_i,
  cache_miss_o,
  miss_addr_o,
  tr_data_received_i,
  cce_data_received_i,
  uncached_data_received_i,
  set_tag_received_i,
  set_tag_wakeup_received_i,
  lce_req_o,
  lce_req_v_o,
  lce_req_ready_i,
  lce_resp_o,
  lce_resp_v_o,
  lce_resp_yumi_i
);

  input [0:0] id_i;
  input [38:0] miss_addr_i;
  input [2:0] lru_way_i;
  output [38:0] miss_addr_o;
  output [113:0] lce_req_o;
  output [42:0] lce_resp_o;
  input clk_i;
  input reset_i;
  input miss_i;
  input uncached_req_i;
  input tr_data_received_i;
  input cce_data_received_i;
  input uncached_data_received_i;
  input set_tag_received_i;
  input set_tag_wakeup_received_i;
  input lce_req_ready_i;
  input lce_resp_yumi_i;
  output cache_miss_o;
  output lce_req_v_o;
  output lce_resp_v_o;
  wire [113:0] lce_req_o;
  wire cache_miss_o,lce_req_v_o,lce_resp_v_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,
  tr_data_received_n,cce_data_received_n,set_tag_received_n,tr_data_received,
  cce_data_received,set_tag_received,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,
  N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,
  N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,
  N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,
  N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,
  N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114;
  wire [2:0] state_n;
  reg [42:0] lce_resp_o;
  reg [2:0] lru_way_r,state_r;
  reg lru_flopped_r,tr_data_received_r,cce_data_received_r,set_tag_received_r;
  reg [38:0] miss_addr_o;
  assign lce_resp_o[40] = 1'b1;
  assign lce_req_o[46] = 1'b1;
  assign lce_req_o[3] = 1'b0;
  assign lce_req_o[47] = 1'b0;
  assign lce_req_o[48] = 1'b0;
  assign lce_req_o[49] = 1'b0;
  assign lce_req_o[50] = 1'b0;
  assign lce_req_o[51] = 1'b0;
  assign lce_req_o[52] = 1'b0;
  assign lce_req_o[53] = 1'b0;
  assign lce_req_o[54] = 1'b0;
  assign lce_req_o[55] = 1'b0;
  assign lce_req_o[56] = 1'b0;
  assign lce_req_o[57] = 1'b0;
  assign lce_req_o[58] = 1'b0;
  assign lce_req_o[59] = 1'b0;
  assign lce_req_o[60] = 1'b0;
  assign lce_req_o[61] = 1'b0;
  assign lce_req_o[62] = 1'b0;
  assign lce_req_o[63] = 1'b0;
  assign lce_req_o[64] = 1'b0;
  assign lce_req_o[65] = 1'b0;
  assign lce_req_o[66] = 1'b0;
  assign lce_req_o[67] = 1'b0;
  assign lce_req_o[68] = 1'b0;
  assign lce_req_o[69] = 1'b0;
  assign lce_req_o[70] = 1'b0;
  assign lce_req_o[71] = 1'b0;
  assign lce_req_o[72] = 1'b0;
  assign lce_req_o[73] = 1'b0;
  assign lce_req_o[74] = 1'b0;
  assign lce_req_o[75] = 1'b0;
  assign lce_req_o[76] = 1'b0;
  assign lce_req_o[77] = 1'b0;
  assign lce_req_o[78] = 1'b0;
  assign lce_req_o[79] = 1'b0;
  assign lce_req_o[80] = 1'b0;
  assign lce_req_o[81] = 1'b0;
  assign lce_req_o[82] = 1'b0;
  assign lce_req_o[83] = 1'b0;
  assign lce_req_o[84] = 1'b0;
  assign lce_req_o[85] = 1'b0;
  assign lce_req_o[86] = 1'b0;
  assign lce_req_o[87] = 1'b0;
  assign lce_req_o[88] = 1'b0;
  assign lce_req_o[89] = 1'b0;
  assign lce_req_o[90] = 1'b0;
  assign lce_req_o[91] = 1'b0;
  assign lce_req_o[92] = 1'b0;
  assign lce_req_o[93] = 1'b0;
  assign lce_req_o[94] = 1'b0;
  assign lce_req_o[95] = 1'b0;
  assign lce_req_o[96] = 1'b0;
  assign lce_req_o[97] = 1'b0;
  assign lce_req_o[98] = 1'b0;
  assign lce_req_o[99] = 1'b0;
  assign lce_req_o[100] = 1'b0;
  assign lce_req_o[101] = 1'b0;
  assign lce_req_o[102] = 1'b0;
  assign lce_req_o[103] = 1'b0;
  assign lce_req_o[104] = 1'b0;
  assign lce_req_o[105] = 1'b0;
  assign lce_req_o[106] = 1'b0;
  assign lce_req_o[107] = 1'b0;
  assign lce_req_o[108] = 1'b0;
  assign lce_req_o[109] = 1'b0;
  assign lce_req_o[110] = 1'b0;
  assign lce_req_o[111] = 1'b0;
  assign lce_resp_o[38] = miss_addr_o[38];
  assign lce_req_o[45] = miss_addr_o[38];
  assign lce_resp_o[37] = miss_addr_o[37];
  assign lce_req_o[44] = miss_addr_o[37];
  assign lce_resp_o[36] = miss_addr_o[36];
  assign lce_req_o[43] = miss_addr_o[36];
  assign lce_resp_o[35] = miss_addr_o[35];
  assign lce_req_o[42] = miss_addr_o[35];
  assign lce_resp_o[34] = miss_addr_o[34];
  assign lce_req_o[41] = miss_addr_o[34];
  assign lce_resp_o[33] = miss_addr_o[33];
  assign lce_req_o[40] = miss_addr_o[33];
  assign lce_resp_o[32] = miss_addr_o[32];
  assign lce_req_o[39] = miss_addr_o[32];
  assign lce_resp_o[31] = miss_addr_o[31];
  assign lce_req_o[38] = miss_addr_o[31];
  assign lce_resp_o[30] = miss_addr_o[30];
  assign lce_req_o[37] = miss_addr_o[30];
  assign lce_resp_o[29] = miss_addr_o[29];
  assign lce_req_o[36] = miss_addr_o[29];
  assign lce_resp_o[28] = miss_addr_o[28];
  assign lce_req_o[35] = miss_addr_o[28];
  assign lce_resp_o[27] = miss_addr_o[27];
  assign lce_req_o[34] = miss_addr_o[27];
  assign lce_resp_o[26] = miss_addr_o[26];
  assign lce_req_o[33] = miss_addr_o[26];
  assign lce_resp_o[25] = miss_addr_o[25];
  assign lce_req_o[32] = miss_addr_o[25];
  assign lce_resp_o[24] = miss_addr_o[24];
  assign lce_req_o[31] = miss_addr_o[24];
  assign lce_resp_o[23] = miss_addr_o[23];
  assign lce_req_o[30] = miss_addr_o[23];
  assign lce_resp_o[22] = miss_addr_o[22];
  assign lce_req_o[29] = miss_addr_o[22];
  assign lce_resp_o[21] = miss_addr_o[21];
  assign lce_req_o[28] = miss_addr_o[21];
  assign lce_resp_o[20] = miss_addr_o[20];
  assign lce_req_o[27] = miss_addr_o[20];
  assign lce_resp_o[19] = miss_addr_o[19];
  assign lce_req_o[26] = miss_addr_o[19];
  assign lce_resp_o[18] = miss_addr_o[18];
  assign lce_req_o[25] = miss_addr_o[18];
  assign lce_resp_o[17] = miss_addr_o[17];
  assign lce_req_o[24] = miss_addr_o[17];
  assign lce_resp_o[16] = miss_addr_o[16];
  assign lce_req_o[23] = miss_addr_o[16];
  assign lce_resp_o[15] = miss_addr_o[15];
  assign lce_req_o[22] = miss_addr_o[15];
  assign lce_resp_o[14] = miss_addr_o[14];
  assign lce_req_o[21] = miss_addr_o[14];
  assign lce_resp_o[13] = miss_addr_o[13];
  assign lce_req_o[20] = miss_addr_o[13];
  assign lce_resp_o[12] = miss_addr_o[12];
  assign lce_req_o[19] = miss_addr_o[12];
  assign lce_resp_o[11] = miss_addr_o[11];
  assign lce_req_o[18] = miss_addr_o[11];
  assign lce_resp_o[10] = miss_addr_o[10];
  assign lce_req_o[17] = miss_addr_o[10];
  assign lce_resp_o[9] = miss_addr_o[9];
  assign lce_req_o[16] = miss_addr_o[9];
  assign lce_resp_o[8] = miss_addr_o[8];
  assign lce_req_o[15] = miss_addr_o[8];
  assign lce_resp_o[7] = miss_addr_o[7];
  assign lce_req_o[14] = miss_addr_o[7];
  assign lce_resp_o[6] = miss_addr_o[6];
  assign lce_req_o[13] = miss_addr_o[6];
  assign lce_resp_o[5] = miss_addr_o[5];
  assign lce_req_o[12] = miss_addr_o[5];
  assign lce_resp_o[4] = miss_addr_o[4];
  assign lce_req_o[11] = miss_addr_o[4];
  assign lce_resp_o[3] = miss_addr_o[3];
  assign lce_req_o[10] = miss_addr_o[3];
  assign lce_resp_o[2] = miss_addr_o[2];
  assign lce_resp_o[1] = miss_addr_o[1];
  assign lce_resp_o[0] = miss_addr_o[0];
  assign lce_resp_o[41] = id_i[0];
  assign lce_req_o[112] = id_i[0];
  assign lce_req_o[113] = lce_resp_o[42];
  assign N20 = N17 & N18;
  assign N21 = N20 & N19;
  assign N22 = state_r[2] | state_r[1];
  assign N23 = N22 | N19;
  assign N25 = N17 | state_r[1];
  assign N26 = N25 | state_r[0];
  assign N28 = N17 | state_r[1];
  assign N29 = N28 | N19;
  assign N31 = state_r[2] | N18;
  assign N32 = N31 | state_r[0];
  assign N34 = state_r[2] | N18;
  assign N35 = N34 | N19;
  assign N37 = state_r[2] & state_r[1];
  assign { N16, N15, N14 } = (N0)? lru_way_r : 
                             (N1)? lru_way_i : 1'b0;
  assign N0 = lru_flopped_r;
  assign N1 = N13;
  assign { N41, N40 } = (N2)? { 1'b0, 1'b1 } : 
                        (N59)? { 1'b1, 1'b0 } : 1'b0;
  assign N2 = miss_i;
  assign N42 = (N2)? 1'b1 : 
               (N59)? 1'b1 : 
               (N39)? 1'b0 : 1'b0;
  assign { N53, N52, N51 } = (N3)? { 1'b0, 1'b1, 1'b0 } : 
                             (N66)? { 1'b0, 1'b1, 1'b1 } : 
                             (N50)? { 1'b1, 1'b0, 1'b1 } : 1'b0;
  assign N3 = tr_data_received;
  assign { N56, N55, N54 } = (N4)? { 1'b0, 1'b1, 1'b1 } : 
                             (N61)? { 1'b0, 1'b0, 1'b0 } : 
                             (N64)? { N53, N52, N51 } : 
                             (N48)? { 1'b1, 1'b0, 1'b1 } : 1'b0;
  assign N4 = set_tag_wakeup_received_i;
  assign cache_miss_o = (N5)? N42 : 
                        (N6)? 1'b1 : 
                        (N7)? 1'b1 : 
                        (N8)? 1'b1 : 
                        (N9)? 1'b1 : 
                        (N10)? 1'b1 : 
                        (N11)? 1'b0 : 1'b0;
  assign N5 = N21;
  assign N6 = N24;
  assign N7 = N27;
  assign N8 = N30;
  assign N9 = N33;
  assign N10 = N36;
  assign N11 = N37;
  assign tr_data_received_n = (N5)? 1'b0 : 
                              (N8)? 1'b1 : 1'b0;
  assign cce_data_received_n = (N5)? 1'b0 : 
                               (N8)? 1'b1 : 1'b0;
  assign set_tag_received_n = (N5)? 1'b0 : 
                              (N8)? 1'b1 : 1'b0;
  assign state_n = (N5)? { N41, 1'b0, N40 } : 
                   (N6)? { lce_req_ready_i, 1'b0, 1'b1 } : 
                   (N7)? { 1'b1, 1'b0, lce_req_ready_i } : 
                   (N8)? { N56, N55, N54 } : 
                   (N9)? { 1'b0, N57, 1'b0 } : 
                   (N10)? { 1'b0, N57, N57 } : 
                   (N11)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign lce_req_v_o = (N5)? 1'b0 : 
                       (N6)? 1'b1 : 
                       (N7)? 1'b1 : 
                       (N8)? 1'b0 : 
                       (N9)? 1'b0 : 
                       (N10)? 1'b0 : 
                       (N11)? 1'b0 : 1'b0;
  assign { lce_req_o[9:4], lce_req_o[2:0] } = (N5)? { miss_addr_o[2:0], N16, N15, N14, 1'b0, 1'b0, 1'b0 } : 
                                              (N6)? { miss_addr_o[2:0], N16, N15, N14, 1'b0, 1'b0, 1'b0 } : 
                                              (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1 } : 
                                              (N8)? { miss_addr_o[2:0], N16, N15, N14, 1'b0, 1'b0, 1'b0 } : 
                                              (N9)? { miss_addr_o[2:0], N16, N15, N14, 1'b0, 1'b0, 1'b0 } : 
                                              (N10)? { miss_addr_o[2:0], N16, N15, N14, 1'b0, 1'b0, 1'b0 } : 
                                              (N11)? { miss_addr_o[2:0], N16, N15, N14, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign lce_resp_v_o = (N5)? 1'b0 : 
                        (N6)? 1'b0 : 
                        (N7)? 1'b0 : 
                        (N8)? 1'b0 : 
                        (N9)? 1'b1 : 
                        (N10)? 1'b1 : 
                        (N11)? 1'b0 : 1'b0;
  assign lce_resp_o[39] = (N5)? 1'b0 : 
                          (N6)? 1'b0 : 
                          (N7)? 1'b0 : 
                          (N8)? 1'b0 : 
                          (N9)? 1'b0 : 
                          (N10)? 1'b1 : 
                          (N11)? 1'b0 : 1'b0;
  assign N12 = 1'b0;
  assign tr_data_received = tr_data_received_r | tr_data_received_i;
  assign cce_data_received = cce_data_received_r | cce_data_received_i;
  assign set_tag_received = set_tag_received_r | set_tag_received_i;
  assign N13 = ~lru_flopped_r;
  assign N17 = ~state_r[2];
  assign N18 = ~state_r[1];
  assign N19 = ~state_r[0];
  assign N24 = ~N23;
  assign N27 = ~N26;
  assign N30 = ~N29;
  assign N33 = ~N32;
  assign N36 = ~N35;
  assign N38 = uncached_req_i | miss_i;
  assign N39 = ~N38;
  assign N43 = ~tr_data_received_i;
  assign N44 = ~cce_data_received_i;
  assign N45 = ~set_tag_received_i;
  assign N46 = uncached_data_received_i | set_tag_wakeup_received_i;
  assign N47 = set_tag_received | N46;
  assign N48 = ~N47;
  assign N49 = cce_data_received | tr_data_received;
  assign N50 = ~N49;
  assign N57 = ~lce_resp_yumi_i;
  assign N58 = ~miss_i;
  assign N59 = uncached_req_i & N58;
  assign N60 = ~set_tag_wakeup_received_i;
  assign N61 = uncached_data_received_i & N60;
  assign N62 = ~uncached_data_received_i;
  assign N63 = N60 & N62;
  assign N64 = set_tag_received & N63;
  assign N65 = ~tr_data_received;
  assign N66 = cce_data_received & N65;
  assign N67 = ~reset_i;
  assign N68 = N21 & N67;
  assign N69 = N24 & N67;
  assign N70 = lru_flopped_r & N69;
  assign N71 = N68 | N70;
  assign N72 = N27 & N67;
  assign N73 = N71 | N72;
  assign N74 = N30 & N67;
  assign N75 = N73 | N74;
  assign N76 = N33 & N67;
  assign N77 = N75 | N76;
  assign N78 = N36 & N67;
  assign N79 = N77 | N78;
  assign N80 = N37 & N67;
  assign N81 = N79 | N80;
  assign N82 = ~N81;
  assign N83 = N67 & N82;
  assign N84 = N39 & N21;
  assign N85 = ~N84;
  assign N86 = N84 | N24;
  assign N87 = N86 | N27;
  assign N88 = N43 & N30;
  assign N89 = N87 | N88;
  assign N90 = N89 | N33;
  assign N91 = N90 | N36;
  assign N92 = N91 | N37;
  assign N93 = ~N92;
  assign N94 = N44 & N30;
  assign N95 = N87 | N94;
  assign N96 = N95 | N33;
  assign N97 = N96 | N36;
  assign N98 = N97 | N37;
  assign N99 = ~N98;
  assign N100 = N45 & N30;
  assign N101 = N87 | N100;
  assign N102 = N101 | N33;
  assign N103 = N102 | N36;
  assign N104 = N103 | N37;
  assign N105 = ~N104;
  assign N106 = N39 & N68;
  assign N107 = N106 | N69;
  assign N108 = N107 | N72;
  assign N109 = N108 | N74;
  assign N110 = N109 | N76;
  assign N111 = N110 | N78;
  assign N112 = N111 | N80;
  assign N113 = ~N112;
  assign N114 = N67 & N113;

  always @(posedge clk_i) begin
    if(1'b1) begin
      { lce_resp_o[42:42] } <= { 1'b0 };
    end 
    if(N83) begin
      { lru_way_r[2:0] } <= { lru_way_i[2:0] };
    end 
    if(reset_i) begin
      { state_r[2:0] } <= { 1'b0, 1'b0, 1'b0 };
    end else if(N85) begin
      { state_r[2:0] } <= { state_n[2:0] };
    end 
    if(reset_i) begin
      lru_flopped_r <= 1'b0;
    end else begin
      lru_flopped_r <= N12;
    end
    if(reset_i) begin
      tr_data_received_r <= 1'b0;
    end else if(N93) begin
      tr_data_received_r <= tr_data_received_n;
    end 
    if(reset_i) begin
      cce_data_received_r <= 1'b0;
    end else if(N99) begin
      cce_data_received_r <= cce_data_received_n;
    end 
    if(reset_i) begin
      set_tag_received_r <= 1'b0;
    end else if(N105) begin
      set_tag_received_r <= set_tag_received_n;
    end 
    if(N114) begin
      { miss_addr_o[38:0] } <= { miss_addr_i[38:0] };
    end 
  end


endmodule



module bsg_mem_1r1w_synth_width_p53_els_p2_read_write_same_addr_p0_harden_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [52:0] w_data_i;
  input [0:0] r_addr_i;
  output [52:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [52:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N7,N8;
  reg [105:0] mem;
  assign r_data_o[52] = (N3)? mem[52] : 
                        (N0)? mem[105] : 1'b0;
  assign N0 = r_addr_i[0];
  assign r_data_o[51] = (N3)? mem[51] : 
                        (N0)? mem[104] : 1'b0;
  assign r_data_o[50] = (N3)? mem[50] : 
                        (N0)? mem[103] : 1'b0;
  assign r_data_o[49] = (N3)? mem[49] : 
                        (N0)? mem[102] : 1'b0;
  assign r_data_o[48] = (N3)? mem[48] : 
                        (N0)? mem[101] : 1'b0;
  assign r_data_o[47] = (N3)? mem[47] : 
                        (N0)? mem[100] : 1'b0;
  assign r_data_o[46] = (N3)? mem[46] : 
                        (N0)? mem[99] : 1'b0;
  assign r_data_o[45] = (N3)? mem[45] : 
                        (N0)? mem[98] : 1'b0;
  assign r_data_o[44] = (N3)? mem[44] : 
                        (N0)? mem[97] : 1'b0;
  assign r_data_o[43] = (N3)? mem[43] : 
                        (N0)? mem[96] : 1'b0;
  assign r_data_o[42] = (N3)? mem[42] : 
                        (N0)? mem[95] : 1'b0;
  assign r_data_o[41] = (N3)? mem[41] : 
                        (N0)? mem[94] : 1'b0;
  assign r_data_o[40] = (N3)? mem[40] : 
                        (N0)? mem[93] : 1'b0;
  assign r_data_o[39] = (N3)? mem[39] : 
                        (N0)? mem[92] : 1'b0;
  assign r_data_o[38] = (N3)? mem[38] : 
                        (N0)? mem[91] : 1'b0;
  assign r_data_o[37] = (N3)? mem[37] : 
                        (N0)? mem[90] : 1'b0;
  assign r_data_o[36] = (N3)? mem[36] : 
                        (N0)? mem[89] : 1'b0;
  assign r_data_o[35] = (N3)? mem[35] : 
                        (N0)? mem[88] : 1'b0;
  assign r_data_o[34] = (N3)? mem[34] : 
                        (N0)? mem[87] : 1'b0;
  assign r_data_o[33] = (N3)? mem[33] : 
                        (N0)? mem[86] : 1'b0;
  assign r_data_o[32] = (N3)? mem[32] : 
                        (N0)? mem[85] : 1'b0;
  assign r_data_o[31] = (N3)? mem[31] : 
                        (N0)? mem[84] : 1'b0;
  assign r_data_o[30] = (N3)? mem[30] : 
                        (N0)? mem[83] : 1'b0;
  assign r_data_o[29] = (N3)? mem[29] : 
                        (N0)? mem[82] : 1'b0;
  assign r_data_o[28] = (N3)? mem[28] : 
                        (N0)? mem[81] : 1'b0;
  assign r_data_o[27] = (N3)? mem[27] : 
                        (N0)? mem[80] : 1'b0;
  assign r_data_o[26] = (N3)? mem[26] : 
                        (N0)? mem[79] : 1'b0;
  assign r_data_o[25] = (N3)? mem[25] : 
                        (N0)? mem[78] : 1'b0;
  assign r_data_o[24] = (N3)? mem[24] : 
                        (N0)? mem[77] : 1'b0;
  assign r_data_o[23] = (N3)? mem[23] : 
                        (N0)? mem[76] : 1'b0;
  assign r_data_o[22] = (N3)? mem[22] : 
                        (N0)? mem[75] : 1'b0;
  assign r_data_o[21] = (N3)? mem[21] : 
                        (N0)? mem[74] : 1'b0;
  assign r_data_o[20] = (N3)? mem[20] : 
                        (N0)? mem[73] : 1'b0;
  assign r_data_o[19] = (N3)? mem[19] : 
                        (N0)? mem[72] : 1'b0;
  assign r_data_o[18] = (N3)? mem[18] : 
                        (N0)? mem[71] : 1'b0;
  assign r_data_o[17] = (N3)? mem[17] : 
                        (N0)? mem[70] : 1'b0;
  assign r_data_o[16] = (N3)? mem[16] : 
                        (N0)? mem[69] : 1'b0;
  assign r_data_o[15] = (N3)? mem[15] : 
                        (N0)? mem[68] : 1'b0;
  assign r_data_o[14] = (N3)? mem[14] : 
                        (N0)? mem[67] : 1'b0;
  assign r_data_o[13] = (N3)? mem[13] : 
                        (N0)? mem[66] : 1'b0;
  assign r_data_o[12] = (N3)? mem[12] : 
                        (N0)? mem[65] : 1'b0;
  assign r_data_o[11] = (N3)? mem[11] : 
                        (N0)? mem[64] : 1'b0;
  assign r_data_o[10] = (N3)? mem[10] : 
                        (N0)? mem[63] : 1'b0;
  assign r_data_o[9] = (N3)? mem[9] : 
                       (N0)? mem[62] : 1'b0;
  assign r_data_o[8] = (N3)? mem[8] : 
                       (N0)? mem[61] : 1'b0;
  assign r_data_o[7] = (N3)? mem[7] : 
                       (N0)? mem[60] : 1'b0;
  assign r_data_o[6] = (N3)? mem[6] : 
                       (N0)? mem[59] : 1'b0;
  assign r_data_o[5] = (N3)? mem[5] : 
                       (N0)? mem[58] : 1'b0;
  assign r_data_o[4] = (N3)? mem[4] : 
                       (N0)? mem[57] : 1'b0;
  assign r_data_o[3] = (N3)? mem[3] : 
                       (N0)? mem[56] : 1'b0;
  assign r_data_o[2] = (N3)? mem[2] : 
                       (N0)? mem[55] : 1'b0;
  assign r_data_o[1] = (N3)? mem[1] : 
                       (N0)? mem[54] : 1'b0;
  assign r_data_o[0] = (N3)? mem[0] : 
                       (N0)? mem[53] : 1'b0;
  assign N5 = ~w_addr_i[0];
  assign { N8, N7 } = (N1)? { w_addr_i[0:0], N5 } : 
                      (N2)? { 1'b0, 1'b0 } : 1'b0;
  assign N1 = w_v_i;
  assign N2 = N4;
  assign N3 = ~r_addr_i[0];
  assign N4 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N8) begin
      { mem[105:53] } <= { w_data_i[52:0] };
    end 
    if(N7) begin
      { mem[52:0] } <= { w_data_i[52:0] };
    end 
  end


endmodule



module bsg_mem_1r1w_width_p53_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [52:0] w_data_i;
  input [0:0] r_addr_i;
  output [52:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [52:0] r_data_o;

  bsg_mem_1r1w_synth_width_p53_els_p2_read_write_same_addr_p0_harden_p0
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i[0]),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i[0]),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_two_fifo_width_p53
(
  clk_i,
  reset_i,
  ready_o,
  data_i,
  v_i,
  v_o,
  data_o,
  yumi_i
);

  input [52:0] data_i;
  output [52:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [52:0] data_o;
  wire ready_o,v_o,N0,N1,enq_i,n_0_net_,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,
  N15,N16,N17,N18,N19,N20,N21,N22,N23,N24;
  reg full_r,tail_r,head_r,empty_r;

  bsg_mem_1r1w_width_p53_els_p2_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enq_i),
    .w_addr_i(tail_r),
    .w_data_i(data_i),
    .r_v_i(n_0_net_),
    .r_addr_i(head_r),
    .r_data_o(data_o)
  );

  assign N9 = (N0)? 1'b1 : 
              (N1)? N5 : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign N10 = (N0)? 1'b0 : 
               (N1)? N4 : 1'b0;
  assign N11 = (N0)? 1'b1 : 
               (N1)? yumi_i : 1'b0;
  assign N12 = (N0)? 1'b0 : 
               (N1)? N6 : 1'b0;
  assign N13 = (N0)? 1'b1 : 
               (N1)? N7 : 1'b0;
  assign N14 = (N0)? 1'b0 : 
               (N1)? N8 : 1'b0;
  assign n_0_net_ = ~empty_r;
  assign v_o = ~empty_r;
  assign ready_o = ~full_r;
  assign enq_i = v_i & N15;
  assign N15 = ~full_r;
  assign N2 = ~reset_i;
  assign N3 = reset_i;
  assign N5 = enq_i;
  assign N4 = ~tail_r;
  assign N6 = ~head_r;
  assign N7 = N17 | N19;
  assign N17 = empty_r & N16;
  assign N16 = ~enq_i;
  assign N19 = N18 & N16;
  assign N18 = N15 & yumi_i;
  assign N8 = N23 | N24;
  assign N23 = N21 & N22;
  assign N21 = N20 & enq_i;
  assign N20 = ~empty_r;
  assign N22 = ~yumi_i;
  assign N24 = full_r & N22;

  always @(posedge clk_i) begin
    if(1'b1) begin
      full_r <= N14;
      empty_r <= N13;
    end 
    if(N9) begin
      tail_r <= N10;
    end 
    if(N11) begin
      head_r <= N12;
    end 
  end


endmodule



module bp_fe_lce_cmd_02
(
  clk_i,
  reset_i,
  id_i,
  lce_ready_o,
  set_tag_received_o,
  set_tag_wakeup_received_o,
  data_mem_data_i,
  data_mem_pkt_o,
  data_mem_pkt_v_o,
  data_mem_pkt_yumi_i,
  tag_mem_pkt_o,
  tag_mem_pkt_v_o,
  tag_mem_pkt_yumi_i,
  stat_mem_pkt_v_o,
  stat_mem_pkt_o,
  stat_mem_pkt_yumi_i,
  lce_resp_o,
  lce_resp_v_o,
  lce_resp_yumi_i,
  lce_data_resp_o,
  lce_data_resp_v_o,
  lce_data_resp_ready_i,
  lce_cmd_i,
  lce_cmd_v_i,
  lce_cmd_ready_o,
  lce_data_cmd_o,
  lce_data_cmd_v_o,
  lce_data_cmd_ready_i
);

  input [0:0] id_i;
  input [511:0] data_mem_data_i;
  output [522:0] data_mem_pkt_o;
  output [39:0] tag_mem_pkt_o;
  output [9:0] stat_mem_pkt_o;
  output [42:0] lce_resp_o;
  output [553:0] lce_data_resp_o;
  input [52:0] lce_cmd_i;
  output [517:0] lce_data_cmd_o;
  input clk_i;
  input reset_i;
  input data_mem_pkt_yumi_i;
  input tag_mem_pkt_yumi_i;
  input stat_mem_pkt_yumi_i;
  input lce_resp_yumi_i;
  input lce_data_resp_ready_i;
  input lce_cmd_v_i;
  input lce_data_cmd_ready_i;
  output lce_ready_o;
  output set_tag_received_o;
  output set_tag_wakeup_received_o;
  output data_mem_pkt_v_o;
  output tag_mem_pkt_v_o;
  output stat_mem_pkt_v_o;
  output lce_resp_v_o;
  output lce_data_resp_v_o;
  output lce_cmd_ready_o;
  output lce_data_cmd_v_o;
  wire [522:0] data_mem_pkt_o;
  wire [39:0] tag_mem_pkt_o;
  wire [9:0] stat_mem_pkt_o;
  wire [42:0] lce_resp_o;
  wire [553:0] lce_data_resp_o;
  wire [517:0] lce_data_cmd_o;
  wire lce_ready_o,set_tag_received_o,set_tag_wakeup_received_o,data_mem_pkt_v_o,
  tag_mem_pkt_v_o,stat_mem_pkt_v_o,lce_resp_v_o,lce_data_resp_v_o,lce_cmd_ready_o,
  lce_data_cmd_v_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,
  N19,N20,N21,lce_cmd_li_dst_id__0_,lce_cmd_li_src_id__0_,lce_cmd_li_msg_type__2_,
  lce_cmd_li_msg_type__1_,lce_cmd_li_msg_type__0_,lce_cmd_li_addr__5_,
  lce_cmd_li_addr__4_,lce_cmd_li_addr__3_,lce_cmd_li_addr__2_,lce_cmd_li_addr__1_,
  lce_cmd_li_addr__0_,lce_cmd_li_way_id__2_,lce_cmd_li_way_id__1_,lce_cmd_li_way_id__0_,
  lce_cmd_li_state__1_,lce_cmd_li_state__0_,lce_cmd_li_target__0_,
  lce_cmd_li_target_way_id__2_,lce_cmd_li_target_way_id__1_,lce_cmd_li_target_way_id__0_,lce_cmd_yumi_lo,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,lce_cmd_v_li,N35,N36,N37,N38,
  N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,
  N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,
  N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,
  N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,
  N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,
  N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,
  N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,
  N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,
  N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,
  N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,
  N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,
  N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,
  N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,
  N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,
  N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,
  N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,
  N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,
  N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,
  N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,
  N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,
  N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,
  N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,
  N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,
  N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,
  N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,
  N451,N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,
  N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,
  N483,N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,
  N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,
  N515,N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,
  N531,N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,
  N547,N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,
  N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,
  N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,
  N595,N596,N597,N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,
  N611,N612,N613,N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,
  N627,N628,N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,
  N643,N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,
  N659,N660,N661,N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,
  N675,N676,N677,N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,
  N691,N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,
  N707,N708,N709,N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,
  N723,N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,
  N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,
  N755,N756,N757,N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,N769,N770,
  N771,N772,N773,N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,N785,N786,
  N787,N788,N789,N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,N801,N802,
  N803,N804,N805,N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,N817,N818,
  N819,N820,N821,N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,N833,N835,
  N836,N837,N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,N849,N850,N851,
  N852,N853,N854,N855,N856,N857,N858,N859;
  wire [5:0] lce_cmd_addr_index;
  wire [26:0] lce_cmd_addr_tag;
  wire [1:0] state_n;
  reg [511:0] data_r;
  reg [1:0] state_r;
  reg [0:0] syn_ack_cnt_r;
  reg flag_data_buffered_r,flag_invalidate_r;
  assign stat_mem_pkt_o[0] = 1'b0;
  assign stat_mem_pkt_o[1] = 1'b0;
  assign stat_mem_pkt_o[2] = 1'b0;
  assign stat_mem_pkt_o[3] = 1'b0;
  assign data_mem_pkt_o[1] = 1'b0;
  assign data_mem_pkt_o[2] = 1'b0;
  assign data_mem_pkt_o[3] = 1'b0;
  assign data_mem_pkt_o[4] = 1'b0;
  assign data_mem_pkt_o[5] = 1'b0;
  assign data_mem_pkt_o[6] = 1'b0;
  assign data_mem_pkt_o[7] = 1'b0;
  assign data_mem_pkt_o[8] = 1'b0;
  assign data_mem_pkt_o[9] = 1'b0;
  assign data_mem_pkt_o[10] = 1'b0;
  assign data_mem_pkt_o[11] = 1'b0;
  assign data_mem_pkt_o[12] = 1'b0;
  assign data_mem_pkt_o[13] = 1'b0;
  assign data_mem_pkt_o[14] = 1'b0;
  assign data_mem_pkt_o[15] = 1'b0;
  assign data_mem_pkt_o[16] = 1'b0;
  assign data_mem_pkt_o[17] = 1'b0;
  assign data_mem_pkt_o[18] = 1'b0;
  assign data_mem_pkt_o[19] = 1'b0;
  assign data_mem_pkt_o[20] = 1'b0;
  assign data_mem_pkt_o[21] = 1'b0;
  assign data_mem_pkt_o[22] = 1'b0;
  assign data_mem_pkt_o[23] = 1'b0;
  assign data_mem_pkt_o[24] = 1'b0;
  assign data_mem_pkt_o[25] = 1'b0;
  assign data_mem_pkt_o[26] = 1'b0;
  assign data_mem_pkt_o[27] = 1'b0;
  assign data_mem_pkt_o[28] = 1'b0;
  assign data_mem_pkt_o[29] = 1'b0;
  assign data_mem_pkt_o[30] = 1'b0;
  assign data_mem_pkt_o[31] = 1'b0;
  assign data_mem_pkt_o[32] = 1'b0;
  assign data_mem_pkt_o[33] = 1'b0;
  assign data_mem_pkt_o[34] = 1'b0;
  assign data_mem_pkt_o[35] = 1'b0;
  assign data_mem_pkt_o[36] = 1'b0;
  assign data_mem_pkt_o[37] = 1'b0;
  assign data_mem_pkt_o[38] = 1'b0;
  assign data_mem_pkt_o[39] = 1'b0;
  assign data_mem_pkt_o[40] = 1'b0;
  assign data_mem_pkt_o[41] = 1'b0;
  assign data_mem_pkt_o[42] = 1'b0;
  assign data_mem_pkt_o[43] = 1'b0;
  assign data_mem_pkt_o[44] = 1'b0;
  assign data_mem_pkt_o[45] = 1'b0;
  assign data_mem_pkt_o[46] = 1'b0;
  assign data_mem_pkt_o[47] = 1'b0;
  assign data_mem_pkt_o[48] = 1'b0;
  assign data_mem_pkt_o[49] = 1'b0;
  assign data_mem_pkt_o[50] = 1'b0;
  assign data_mem_pkt_o[51] = 1'b0;
  assign data_mem_pkt_o[52] = 1'b0;
  assign data_mem_pkt_o[53] = 1'b0;
  assign data_mem_pkt_o[54] = 1'b0;
  assign data_mem_pkt_o[55] = 1'b0;
  assign data_mem_pkt_o[56] = 1'b0;
  assign data_mem_pkt_o[57] = 1'b0;
  assign data_mem_pkt_o[58] = 1'b0;
  assign data_mem_pkt_o[59] = 1'b0;
  assign data_mem_pkt_o[60] = 1'b0;
  assign data_mem_pkt_o[61] = 1'b0;
  assign data_mem_pkt_o[62] = 1'b0;
  assign data_mem_pkt_o[63] = 1'b0;
  assign data_mem_pkt_o[64] = 1'b0;
  assign data_mem_pkt_o[65] = 1'b0;
  assign data_mem_pkt_o[66] = 1'b0;
  assign data_mem_pkt_o[67] = 1'b0;
  assign data_mem_pkt_o[68] = 1'b0;
  assign data_mem_pkt_o[69] = 1'b0;
  assign data_mem_pkt_o[70] = 1'b0;
  assign data_mem_pkt_o[71] = 1'b0;
  assign data_mem_pkt_o[72] = 1'b0;
  assign data_mem_pkt_o[73] = 1'b0;
  assign data_mem_pkt_o[74] = 1'b0;
  assign data_mem_pkt_o[75] = 1'b0;
  assign data_mem_pkt_o[76] = 1'b0;
  assign data_mem_pkt_o[77] = 1'b0;
  assign data_mem_pkt_o[78] = 1'b0;
  assign data_mem_pkt_o[79] = 1'b0;
  assign data_mem_pkt_o[80] = 1'b0;
  assign data_mem_pkt_o[81] = 1'b0;
  assign data_mem_pkt_o[82] = 1'b0;
  assign data_mem_pkt_o[83] = 1'b0;
  assign data_mem_pkt_o[84] = 1'b0;
  assign data_mem_pkt_o[85] = 1'b0;
  assign data_mem_pkt_o[86] = 1'b0;
  assign data_mem_pkt_o[87] = 1'b0;
  assign data_mem_pkt_o[88] = 1'b0;
  assign data_mem_pkt_o[89] = 1'b0;
  assign data_mem_pkt_o[90] = 1'b0;
  assign data_mem_pkt_o[91] = 1'b0;
  assign data_mem_pkt_o[92] = 1'b0;
  assign data_mem_pkt_o[93] = 1'b0;
  assign data_mem_pkt_o[94] = 1'b0;
  assign data_mem_pkt_o[95] = 1'b0;
  assign data_mem_pkt_o[96] = 1'b0;
  assign data_mem_pkt_o[97] = 1'b0;
  assign data_mem_pkt_o[98] = 1'b0;
  assign data_mem_pkt_o[99] = 1'b0;
  assign data_mem_pkt_o[100] = 1'b0;
  assign data_mem_pkt_o[101] = 1'b0;
  assign data_mem_pkt_o[102] = 1'b0;
  assign data_mem_pkt_o[103] = 1'b0;
  assign data_mem_pkt_o[104] = 1'b0;
  assign data_mem_pkt_o[105] = 1'b0;
  assign data_mem_pkt_o[106] = 1'b0;
  assign data_mem_pkt_o[107] = 1'b0;
  assign data_mem_pkt_o[108] = 1'b0;
  assign data_mem_pkt_o[109] = 1'b0;
  assign data_mem_pkt_o[110] = 1'b0;
  assign data_mem_pkt_o[111] = 1'b0;
  assign data_mem_pkt_o[112] = 1'b0;
  assign data_mem_pkt_o[113] = 1'b0;
  assign data_mem_pkt_o[114] = 1'b0;
  assign data_mem_pkt_o[115] = 1'b0;
  assign data_mem_pkt_o[116] = 1'b0;
  assign data_mem_pkt_o[117] = 1'b0;
  assign data_mem_pkt_o[118] = 1'b0;
  assign data_mem_pkt_o[119] = 1'b0;
  assign data_mem_pkt_o[120] = 1'b0;
  assign data_mem_pkt_o[121] = 1'b0;
  assign data_mem_pkt_o[122] = 1'b0;
  assign data_mem_pkt_o[123] = 1'b0;
  assign data_mem_pkt_o[124] = 1'b0;
  assign data_mem_pkt_o[125] = 1'b0;
  assign data_mem_pkt_o[126] = 1'b0;
  assign data_mem_pkt_o[127] = 1'b0;
  assign data_mem_pkt_o[128] = 1'b0;
  assign data_mem_pkt_o[129] = 1'b0;
  assign data_mem_pkt_o[130] = 1'b0;
  assign data_mem_pkt_o[131] = 1'b0;
  assign data_mem_pkt_o[132] = 1'b0;
  assign data_mem_pkt_o[133] = 1'b0;
  assign data_mem_pkt_o[134] = 1'b0;
  assign data_mem_pkt_o[135] = 1'b0;
  assign data_mem_pkt_o[136] = 1'b0;
  assign data_mem_pkt_o[137] = 1'b0;
  assign data_mem_pkt_o[138] = 1'b0;
  assign data_mem_pkt_o[139] = 1'b0;
  assign data_mem_pkt_o[140] = 1'b0;
  assign data_mem_pkt_o[141] = 1'b0;
  assign data_mem_pkt_o[142] = 1'b0;
  assign data_mem_pkt_o[143] = 1'b0;
  assign data_mem_pkt_o[144] = 1'b0;
  assign data_mem_pkt_o[145] = 1'b0;
  assign data_mem_pkt_o[146] = 1'b0;
  assign data_mem_pkt_o[147] = 1'b0;
  assign data_mem_pkt_o[148] = 1'b0;
  assign data_mem_pkt_o[149] = 1'b0;
  assign data_mem_pkt_o[150] = 1'b0;
  assign data_mem_pkt_o[151] = 1'b0;
  assign data_mem_pkt_o[152] = 1'b0;
  assign data_mem_pkt_o[153] = 1'b0;
  assign data_mem_pkt_o[154] = 1'b0;
  assign data_mem_pkt_o[155] = 1'b0;
  assign data_mem_pkt_o[156] = 1'b0;
  assign data_mem_pkt_o[157] = 1'b0;
  assign data_mem_pkt_o[158] = 1'b0;
  assign data_mem_pkt_o[159] = 1'b0;
  assign data_mem_pkt_o[160] = 1'b0;
  assign data_mem_pkt_o[161] = 1'b0;
  assign data_mem_pkt_o[162] = 1'b0;
  assign data_mem_pkt_o[163] = 1'b0;
  assign data_mem_pkt_o[164] = 1'b0;
  assign data_mem_pkt_o[165] = 1'b0;
  assign data_mem_pkt_o[166] = 1'b0;
  assign data_mem_pkt_o[167] = 1'b0;
  assign data_mem_pkt_o[168] = 1'b0;
  assign data_mem_pkt_o[169] = 1'b0;
  assign data_mem_pkt_o[170] = 1'b0;
  assign data_mem_pkt_o[171] = 1'b0;
  assign data_mem_pkt_o[172] = 1'b0;
  assign data_mem_pkt_o[173] = 1'b0;
  assign data_mem_pkt_o[174] = 1'b0;
  assign data_mem_pkt_o[175] = 1'b0;
  assign data_mem_pkt_o[176] = 1'b0;
  assign data_mem_pkt_o[177] = 1'b0;
  assign data_mem_pkt_o[178] = 1'b0;
  assign data_mem_pkt_o[179] = 1'b0;
  assign data_mem_pkt_o[180] = 1'b0;
  assign data_mem_pkt_o[181] = 1'b0;
  assign data_mem_pkt_o[182] = 1'b0;
  assign data_mem_pkt_o[183] = 1'b0;
  assign data_mem_pkt_o[184] = 1'b0;
  assign data_mem_pkt_o[185] = 1'b0;
  assign data_mem_pkt_o[186] = 1'b0;
  assign data_mem_pkt_o[187] = 1'b0;
  assign data_mem_pkt_o[188] = 1'b0;
  assign data_mem_pkt_o[189] = 1'b0;
  assign data_mem_pkt_o[190] = 1'b0;
  assign data_mem_pkt_o[191] = 1'b0;
  assign data_mem_pkt_o[192] = 1'b0;
  assign data_mem_pkt_o[193] = 1'b0;
  assign data_mem_pkt_o[194] = 1'b0;
  assign data_mem_pkt_o[195] = 1'b0;
  assign data_mem_pkt_o[196] = 1'b0;
  assign data_mem_pkt_o[197] = 1'b0;
  assign data_mem_pkt_o[198] = 1'b0;
  assign data_mem_pkt_o[199] = 1'b0;
  assign data_mem_pkt_o[200] = 1'b0;
  assign data_mem_pkt_o[201] = 1'b0;
  assign data_mem_pkt_o[202] = 1'b0;
  assign data_mem_pkt_o[203] = 1'b0;
  assign data_mem_pkt_o[204] = 1'b0;
  assign data_mem_pkt_o[205] = 1'b0;
  assign data_mem_pkt_o[206] = 1'b0;
  assign data_mem_pkt_o[207] = 1'b0;
  assign data_mem_pkt_o[208] = 1'b0;
  assign data_mem_pkt_o[209] = 1'b0;
  assign data_mem_pkt_o[210] = 1'b0;
  assign data_mem_pkt_o[211] = 1'b0;
  assign data_mem_pkt_o[212] = 1'b0;
  assign data_mem_pkt_o[213] = 1'b0;
  assign data_mem_pkt_o[214] = 1'b0;
  assign data_mem_pkt_o[215] = 1'b0;
  assign data_mem_pkt_o[216] = 1'b0;
  assign data_mem_pkt_o[217] = 1'b0;
  assign data_mem_pkt_o[218] = 1'b0;
  assign data_mem_pkt_o[219] = 1'b0;
  assign data_mem_pkt_o[220] = 1'b0;
  assign data_mem_pkt_o[221] = 1'b0;
  assign data_mem_pkt_o[222] = 1'b0;
  assign data_mem_pkt_o[223] = 1'b0;
  assign data_mem_pkt_o[224] = 1'b0;
  assign data_mem_pkt_o[225] = 1'b0;
  assign data_mem_pkt_o[226] = 1'b0;
  assign data_mem_pkt_o[227] = 1'b0;
  assign data_mem_pkt_o[228] = 1'b0;
  assign data_mem_pkt_o[229] = 1'b0;
  assign data_mem_pkt_o[230] = 1'b0;
  assign data_mem_pkt_o[231] = 1'b0;
  assign data_mem_pkt_o[232] = 1'b0;
  assign data_mem_pkt_o[233] = 1'b0;
  assign data_mem_pkt_o[234] = 1'b0;
  assign data_mem_pkt_o[235] = 1'b0;
  assign data_mem_pkt_o[236] = 1'b0;
  assign data_mem_pkt_o[237] = 1'b0;
  assign data_mem_pkt_o[238] = 1'b0;
  assign data_mem_pkt_o[239] = 1'b0;
  assign data_mem_pkt_o[240] = 1'b0;
  assign data_mem_pkt_o[241] = 1'b0;
  assign data_mem_pkt_o[242] = 1'b0;
  assign data_mem_pkt_o[243] = 1'b0;
  assign data_mem_pkt_o[244] = 1'b0;
  assign data_mem_pkt_o[245] = 1'b0;
  assign data_mem_pkt_o[246] = 1'b0;
  assign data_mem_pkt_o[247] = 1'b0;
  assign data_mem_pkt_o[248] = 1'b0;
  assign data_mem_pkt_o[249] = 1'b0;
  assign data_mem_pkt_o[250] = 1'b0;
  assign data_mem_pkt_o[251] = 1'b0;
  assign data_mem_pkt_o[252] = 1'b0;
  assign data_mem_pkt_o[253] = 1'b0;
  assign data_mem_pkt_o[254] = 1'b0;
  assign data_mem_pkt_o[255] = 1'b0;
  assign data_mem_pkt_o[256] = 1'b0;
  assign data_mem_pkt_o[257] = 1'b0;
  assign data_mem_pkt_o[258] = 1'b0;
  assign data_mem_pkt_o[259] = 1'b0;
  assign data_mem_pkt_o[260] = 1'b0;
  assign data_mem_pkt_o[261] = 1'b0;
  assign data_mem_pkt_o[262] = 1'b0;
  assign data_mem_pkt_o[263] = 1'b0;
  assign data_mem_pkt_o[264] = 1'b0;
  assign data_mem_pkt_o[265] = 1'b0;
  assign data_mem_pkt_o[266] = 1'b0;
  assign data_mem_pkt_o[267] = 1'b0;
  assign data_mem_pkt_o[268] = 1'b0;
  assign data_mem_pkt_o[269] = 1'b0;
  assign data_mem_pkt_o[270] = 1'b0;
  assign data_mem_pkt_o[271] = 1'b0;
  assign data_mem_pkt_o[272] = 1'b0;
  assign data_mem_pkt_o[273] = 1'b0;
  assign data_mem_pkt_o[274] = 1'b0;
  assign data_mem_pkt_o[275] = 1'b0;
  assign data_mem_pkt_o[276] = 1'b0;
  assign data_mem_pkt_o[277] = 1'b0;
  assign data_mem_pkt_o[278] = 1'b0;
  assign data_mem_pkt_o[279] = 1'b0;
  assign data_mem_pkt_o[280] = 1'b0;
  assign data_mem_pkt_o[281] = 1'b0;
  assign data_mem_pkt_o[282] = 1'b0;
  assign data_mem_pkt_o[283] = 1'b0;
  assign data_mem_pkt_o[284] = 1'b0;
  assign data_mem_pkt_o[285] = 1'b0;
  assign data_mem_pkt_o[286] = 1'b0;
  assign data_mem_pkt_o[287] = 1'b0;
  assign data_mem_pkt_o[288] = 1'b0;
  assign data_mem_pkt_o[289] = 1'b0;
  assign data_mem_pkt_o[290] = 1'b0;
  assign data_mem_pkt_o[291] = 1'b0;
  assign data_mem_pkt_o[292] = 1'b0;
  assign data_mem_pkt_o[293] = 1'b0;
  assign data_mem_pkt_o[294] = 1'b0;
  assign data_mem_pkt_o[295] = 1'b0;
  assign data_mem_pkt_o[296] = 1'b0;
  assign data_mem_pkt_o[297] = 1'b0;
  assign data_mem_pkt_o[298] = 1'b0;
  assign data_mem_pkt_o[299] = 1'b0;
  assign data_mem_pkt_o[300] = 1'b0;
  assign data_mem_pkt_o[301] = 1'b0;
  assign data_mem_pkt_o[302] = 1'b0;
  assign data_mem_pkt_o[303] = 1'b0;
  assign data_mem_pkt_o[304] = 1'b0;
  assign data_mem_pkt_o[305] = 1'b0;
  assign data_mem_pkt_o[306] = 1'b0;
  assign data_mem_pkt_o[307] = 1'b0;
  assign data_mem_pkt_o[308] = 1'b0;
  assign data_mem_pkt_o[309] = 1'b0;
  assign data_mem_pkt_o[310] = 1'b0;
  assign data_mem_pkt_o[311] = 1'b0;
  assign data_mem_pkt_o[312] = 1'b0;
  assign data_mem_pkt_o[313] = 1'b0;
  assign data_mem_pkt_o[314] = 1'b0;
  assign data_mem_pkt_o[315] = 1'b0;
  assign data_mem_pkt_o[316] = 1'b0;
  assign data_mem_pkt_o[317] = 1'b0;
  assign data_mem_pkt_o[318] = 1'b0;
  assign data_mem_pkt_o[319] = 1'b0;
  assign data_mem_pkt_o[320] = 1'b0;
  assign data_mem_pkt_o[321] = 1'b0;
  assign data_mem_pkt_o[322] = 1'b0;
  assign data_mem_pkt_o[323] = 1'b0;
  assign data_mem_pkt_o[324] = 1'b0;
  assign data_mem_pkt_o[325] = 1'b0;
  assign data_mem_pkt_o[326] = 1'b0;
  assign data_mem_pkt_o[327] = 1'b0;
  assign data_mem_pkt_o[328] = 1'b0;
  assign data_mem_pkt_o[329] = 1'b0;
  assign data_mem_pkt_o[330] = 1'b0;
  assign data_mem_pkt_o[331] = 1'b0;
  assign data_mem_pkt_o[332] = 1'b0;
  assign data_mem_pkt_o[333] = 1'b0;
  assign data_mem_pkt_o[334] = 1'b0;
  assign data_mem_pkt_o[335] = 1'b0;
  assign data_mem_pkt_o[336] = 1'b0;
  assign data_mem_pkt_o[337] = 1'b0;
  assign data_mem_pkt_o[338] = 1'b0;
  assign data_mem_pkt_o[339] = 1'b0;
  assign data_mem_pkt_o[340] = 1'b0;
  assign data_mem_pkt_o[341] = 1'b0;
  assign data_mem_pkt_o[342] = 1'b0;
  assign data_mem_pkt_o[343] = 1'b0;
  assign data_mem_pkt_o[344] = 1'b0;
  assign data_mem_pkt_o[345] = 1'b0;
  assign data_mem_pkt_o[346] = 1'b0;
  assign data_mem_pkt_o[347] = 1'b0;
  assign data_mem_pkt_o[348] = 1'b0;
  assign data_mem_pkt_o[349] = 1'b0;
  assign data_mem_pkt_o[350] = 1'b0;
  assign data_mem_pkt_o[351] = 1'b0;
  assign data_mem_pkt_o[352] = 1'b0;
  assign data_mem_pkt_o[353] = 1'b0;
  assign data_mem_pkt_o[354] = 1'b0;
  assign data_mem_pkt_o[355] = 1'b0;
  assign data_mem_pkt_o[356] = 1'b0;
  assign data_mem_pkt_o[357] = 1'b0;
  assign data_mem_pkt_o[358] = 1'b0;
  assign data_mem_pkt_o[359] = 1'b0;
  assign data_mem_pkt_o[360] = 1'b0;
  assign data_mem_pkt_o[361] = 1'b0;
  assign data_mem_pkt_o[362] = 1'b0;
  assign data_mem_pkt_o[363] = 1'b0;
  assign data_mem_pkt_o[364] = 1'b0;
  assign data_mem_pkt_o[365] = 1'b0;
  assign data_mem_pkt_o[366] = 1'b0;
  assign data_mem_pkt_o[367] = 1'b0;
  assign data_mem_pkt_o[368] = 1'b0;
  assign data_mem_pkt_o[369] = 1'b0;
  assign data_mem_pkt_o[370] = 1'b0;
  assign data_mem_pkt_o[371] = 1'b0;
  assign data_mem_pkt_o[372] = 1'b0;
  assign data_mem_pkt_o[373] = 1'b0;
  assign data_mem_pkt_o[374] = 1'b0;
  assign data_mem_pkt_o[375] = 1'b0;
  assign data_mem_pkt_o[376] = 1'b0;
  assign data_mem_pkt_o[377] = 1'b0;
  assign data_mem_pkt_o[378] = 1'b0;
  assign data_mem_pkt_o[379] = 1'b0;
  assign data_mem_pkt_o[380] = 1'b0;
  assign data_mem_pkt_o[381] = 1'b0;
  assign data_mem_pkt_o[382] = 1'b0;
  assign data_mem_pkt_o[383] = 1'b0;
  assign data_mem_pkt_o[384] = 1'b0;
  assign data_mem_pkt_o[385] = 1'b0;
  assign data_mem_pkt_o[386] = 1'b0;
  assign data_mem_pkt_o[387] = 1'b0;
  assign data_mem_pkt_o[388] = 1'b0;
  assign data_mem_pkt_o[389] = 1'b0;
  assign data_mem_pkt_o[390] = 1'b0;
  assign data_mem_pkt_o[391] = 1'b0;
  assign data_mem_pkt_o[392] = 1'b0;
  assign data_mem_pkt_o[393] = 1'b0;
  assign data_mem_pkt_o[394] = 1'b0;
  assign data_mem_pkt_o[395] = 1'b0;
  assign data_mem_pkt_o[396] = 1'b0;
  assign data_mem_pkt_o[397] = 1'b0;
  assign data_mem_pkt_o[398] = 1'b0;
  assign data_mem_pkt_o[399] = 1'b0;
  assign data_mem_pkt_o[400] = 1'b0;
  assign data_mem_pkt_o[401] = 1'b0;
  assign data_mem_pkt_o[402] = 1'b0;
  assign data_mem_pkt_o[403] = 1'b0;
  assign data_mem_pkt_o[404] = 1'b0;
  assign data_mem_pkt_o[405] = 1'b0;
  assign data_mem_pkt_o[406] = 1'b0;
  assign data_mem_pkt_o[407] = 1'b0;
  assign data_mem_pkt_o[408] = 1'b0;
  assign data_mem_pkt_o[409] = 1'b0;
  assign data_mem_pkt_o[410] = 1'b0;
  assign data_mem_pkt_o[411] = 1'b0;
  assign data_mem_pkt_o[412] = 1'b0;
  assign data_mem_pkt_o[413] = 1'b0;
  assign data_mem_pkt_o[414] = 1'b0;
  assign data_mem_pkt_o[415] = 1'b0;
  assign data_mem_pkt_o[416] = 1'b0;
  assign data_mem_pkt_o[417] = 1'b0;
  assign data_mem_pkt_o[418] = 1'b0;
  assign data_mem_pkt_o[419] = 1'b0;
  assign data_mem_pkt_o[420] = 1'b0;
  assign data_mem_pkt_o[421] = 1'b0;
  assign data_mem_pkt_o[422] = 1'b0;
  assign data_mem_pkt_o[423] = 1'b0;
  assign data_mem_pkt_o[424] = 1'b0;
  assign data_mem_pkt_o[425] = 1'b0;
  assign data_mem_pkt_o[426] = 1'b0;
  assign data_mem_pkt_o[427] = 1'b0;
  assign data_mem_pkt_o[428] = 1'b0;
  assign data_mem_pkt_o[429] = 1'b0;
  assign data_mem_pkt_o[430] = 1'b0;
  assign data_mem_pkt_o[431] = 1'b0;
  assign data_mem_pkt_o[432] = 1'b0;
  assign data_mem_pkt_o[433] = 1'b0;
  assign data_mem_pkt_o[434] = 1'b0;
  assign data_mem_pkt_o[435] = 1'b0;
  assign data_mem_pkt_o[436] = 1'b0;
  assign data_mem_pkt_o[437] = 1'b0;
  assign data_mem_pkt_o[438] = 1'b0;
  assign data_mem_pkt_o[439] = 1'b0;
  assign data_mem_pkt_o[440] = 1'b0;
  assign data_mem_pkt_o[441] = 1'b0;
  assign data_mem_pkt_o[442] = 1'b0;
  assign data_mem_pkt_o[443] = 1'b0;
  assign data_mem_pkt_o[444] = 1'b0;
  assign data_mem_pkt_o[445] = 1'b0;
  assign data_mem_pkt_o[446] = 1'b0;
  assign data_mem_pkt_o[447] = 1'b0;
  assign data_mem_pkt_o[448] = 1'b0;
  assign data_mem_pkt_o[449] = 1'b0;
  assign data_mem_pkt_o[450] = 1'b0;
  assign data_mem_pkt_o[451] = 1'b0;
  assign data_mem_pkt_o[452] = 1'b0;
  assign data_mem_pkt_o[453] = 1'b0;
  assign data_mem_pkt_o[454] = 1'b0;
  assign data_mem_pkt_o[455] = 1'b0;
  assign data_mem_pkt_o[456] = 1'b0;
  assign data_mem_pkt_o[457] = 1'b0;
  assign data_mem_pkt_o[458] = 1'b0;
  assign data_mem_pkt_o[459] = 1'b0;
  assign data_mem_pkt_o[460] = 1'b0;
  assign data_mem_pkt_o[461] = 1'b0;
  assign data_mem_pkt_o[462] = 1'b0;
  assign data_mem_pkt_o[463] = 1'b0;
  assign data_mem_pkt_o[464] = 1'b0;
  assign data_mem_pkt_o[465] = 1'b0;
  assign data_mem_pkt_o[466] = 1'b0;
  assign data_mem_pkt_o[467] = 1'b0;
  assign data_mem_pkt_o[468] = 1'b0;
  assign data_mem_pkt_o[469] = 1'b0;
  assign data_mem_pkt_o[470] = 1'b0;
  assign data_mem_pkt_o[471] = 1'b0;
  assign data_mem_pkt_o[472] = 1'b0;
  assign data_mem_pkt_o[473] = 1'b0;
  assign data_mem_pkt_o[474] = 1'b0;
  assign data_mem_pkt_o[475] = 1'b0;
  assign data_mem_pkt_o[476] = 1'b0;
  assign data_mem_pkt_o[477] = 1'b0;
  assign data_mem_pkt_o[478] = 1'b0;
  assign data_mem_pkt_o[479] = 1'b0;
  assign data_mem_pkt_o[480] = 1'b0;
  assign data_mem_pkt_o[481] = 1'b0;
  assign data_mem_pkt_o[482] = 1'b0;
  assign data_mem_pkt_o[483] = 1'b0;
  assign data_mem_pkt_o[484] = 1'b0;
  assign data_mem_pkt_o[485] = 1'b0;
  assign data_mem_pkt_o[486] = 1'b0;
  assign data_mem_pkt_o[487] = 1'b0;
  assign data_mem_pkt_o[488] = 1'b0;
  assign data_mem_pkt_o[489] = 1'b0;
  assign data_mem_pkt_o[490] = 1'b0;
  assign data_mem_pkt_o[491] = 1'b0;
  assign data_mem_pkt_o[492] = 1'b0;
  assign data_mem_pkt_o[493] = 1'b0;
  assign data_mem_pkt_o[494] = 1'b0;
  assign data_mem_pkt_o[495] = 1'b0;
  assign data_mem_pkt_o[496] = 1'b0;
  assign data_mem_pkt_o[497] = 1'b0;
  assign data_mem_pkt_o[498] = 1'b0;
  assign data_mem_pkt_o[499] = 1'b0;
  assign data_mem_pkt_o[500] = 1'b0;
  assign data_mem_pkt_o[501] = 1'b0;
  assign data_mem_pkt_o[502] = 1'b0;
  assign data_mem_pkt_o[503] = 1'b0;
  assign data_mem_pkt_o[504] = 1'b0;
  assign data_mem_pkt_o[505] = 1'b0;
  assign data_mem_pkt_o[506] = 1'b0;
  assign data_mem_pkt_o[507] = 1'b0;
  assign data_mem_pkt_o[508] = 1'b0;
  assign data_mem_pkt_o[509] = 1'b0;
  assign data_mem_pkt_o[510] = 1'b0;
  assign data_mem_pkt_o[511] = 1'b0;
  assign data_mem_pkt_o[512] = 1'b0;
  assign data_mem_pkt_o[513] = 1'b0;
  assign lce_data_cmd_o[3] = 1'b0;
  assign lce_data_cmd_o[4] = 1'b0;
  assign lce_data_resp_o[42] = 1'b0;
  assign lce_data_resp_o[43] = 1'b0;
  assign lce_data_resp_o[44] = 1'b0;
  assign lce_data_resp_o[45] = 1'b0;
  assign lce_data_resp_o[46] = 1'b0;
  assign lce_data_resp_o[47] = 1'b0;
  assign lce_data_resp_o[48] = 1'b0;
  assign lce_data_resp_o[49] = 1'b0;
  assign lce_data_resp_o[50] = 1'b0;
  assign lce_data_resp_o[51] = 1'b0;
  assign lce_data_resp_o[52] = 1'b0;
  assign lce_data_resp_o[53] = 1'b0;
  assign lce_data_resp_o[54] = 1'b0;
  assign lce_data_resp_o[55] = 1'b0;
  assign lce_data_resp_o[56] = 1'b0;
  assign lce_data_resp_o[57] = 1'b0;
  assign lce_data_resp_o[58] = 1'b0;
  assign lce_data_resp_o[59] = 1'b0;
  assign lce_data_resp_o[60] = 1'b0;
  assign lce_data_resp_o[61] = 1'b0;
  assign lce_data_resp_o[62] = 1'b0;
  assign lce_data_resp_o[63] = 1'b0;
  assign lce_data_resp_o[64] = 1'b0;
  assign lce_data_resp_o[65] = 1'b0;
  assign lce_data_resp_o[66] = 1'b0;
  assign lce_data_resp_o[67] = 1'b0;
  assign lce_data_resp_o[68] = 1'b0;
  assign lce_data_resp_o[69] = 1'b0;
  assign lce_data_resp_o[70] = 1'b0;
  assign lce_data_resp_o[71] = 1'b0;
  assign lce_data_resp_o[72] = 1'b0;
  assign lce_data_resp_o[73] = 1'b0;
  assign lce_data_resp_o[74] = 1'b0;
  assign lce_data_resp_o[75] = 1'b0;
  assign lce_data_resp_o[76] = 1'b0;
  assign lce_data_resp_o[77] = 1'b0;
  assign lce_data_resp_o[78] = 1'b0;
  assign lce_data_resp_o[79] = 1'b0;
  assign lce_data_resp_o[80] = 1'b0;
  assign lce_data_resp_o[81] = 1'b0;
  assign lce_data_resp_o[82] = 1'b0;
  assign lce_data_resp_o[83] = 1'b0;
  assign lce_data_resp_o[84] = 1'b0;
  assign lce_data_resp_o[85] = 1'b0;
  assign lce_data_resp_o[86] = 1'b0;
  assign lce_data_resp_o[87] = 1'b0;
  assign lce_data_resp_o[88] = 1'b0;
  assign lce_data_resp_o[89] = 1'b0;
  assign lce_data_resp_o[90] = 1'b0;
  assign lce_data_resp_o[91] = 1'b0;
  assign lce_data_resp_o[92] = 1'b0;
  assign lce_data_resp_o[93] = 1'b0;
  assign lce_data_resp_o[94] = 1'b0;
  assign lce_data_resp_o[95] = 1'b0;
  assign lce_data_resp_o[96] = 1'b0;
  assign lce_data_resp_o[97] = 1'b0;
  assign lce_data_resp_o[98] = 1'b0;
  assign lce_data_resp_o[99] = 1'b0;
  assign lce_data_resp_o[100] = 1'b0;
  assign lce_data_resp_o[101] = 1'b0;
  assign lce_data_resp_o[102] = 1'b0;
  assign lce_data_resp_o[103] = 1'b0;
  assign lce_data_resp_o[104] = 1'b0;
  assign lce_data_resp_o[105] = 1'b0;
  assign lce_data_resp_o[106] = 1'b0;
  assign lce_data_resp_o[107] = 1'b0;
  assign lce_data_resp_o[108] = 1'b0;
  assign lce_data_resp_o[109] = 1'b0;
  assign lce_data_resp_o[110] = 1'b0;
  assign lce_data_resp_o[111] = 1'b0;
  assign lce_data_resp_o[112] = 1'b0;
  assign lce_data_resp_o[113] = 1'b0;
  assign lce_data_resp_o[114] = 1'b0;
  assign lce_data_resp_o[115] = 1'b0;
  assign lce_data_resp_o[116] = 1'b0;
  assign lce_data_resp_o[117] = 1'b0;
  assign lce_data_resp_o[118] = 1'b0;
  assign lce_data_resp_o[119] = 1'b0;
  assign lce_data_resp_o[120] = 1'b0;
  assign lce_data_resp_o[121] = 1'b0;
  assign lce_data_resp_o[122] = 1'b0;
  assign lce_data_resp_o[123] = 1'b0;
  assign lce_data_resp_o[124] = 1'b0;
  assign lce_data_resp_o[125] = 1'b0;
  assign lce_data_resp_o[126] = 1'b0;
  assign lce_data_resp_o[127] = 1'b0;
  assign lce_data_resp_o[128] = 1'b0;
  assign lce_data_resp_o[129] = 1'b0;
  assign lce_data_resp_o[130] = 1'b0;
  assign lce_data_resp_o[131] = 1'b0;
  assign lce_data_resp_o[132] = 1'b0;
  assign lce_data_resp_o[133] = 1'b0;
  assign lce_data_resp_o[134] = 1'b0;
  assign lce_data_resp_o[135] = 1'b0;
  assign lce_data_resp_o[136] = 1'b0;
  assign lce_data_resp_o[137] = 1'b0;
  assign lce_data_resp_o[138] = 1'b0;
  assign lce_data_resp_o[139] = 1'b0;
  assign lce_data_resp_o[140] = 1'b0;
  assign lce_data_resp_o[141] = 1'b0;
  assign lce_data_resp_o[142] = 1'b0;
  assign lce_data_resp_o[143] = 1'b0;
  assign lce_data_resp_o[144] = 1'b0;
  assign lce_data_resp_o[145] = 1'b0;
  assign lce_data_resp_o[146] = 1'b0;
  assign lce_data_resp_o[147] = 1'b0;
  assign lce_data_resp_o[148] = 1'b0;
  assign lce_data_resp_o[149] = 1'b0;
  assign lce_data_resp_o[150] = 1'b0;
  assign lce_data_resp_o[151] = 1'b0;
  assign lce_data_resp_o[152] = 1'b0;
  assign lce_data_resp_o[153] = 1'b0;
  assign lce_data_resp_o[154] = 1'b0;
  assign lce_data_resp_o[155] = 1'b0;
  assign lce_data_resp_o[156] = 1'b0;
  assign lce_data_resp_o[157] = 1'b0;
  assign lce_data_resp_o[158] = 1'b0;
  assign lce_data_resp_o[159] = 1'b0;
  assign lce_data_resp_o[160] = 1'b0;
  assign lce_data_resp_o[161] = 1'b0;
  assign lce_data_resp_o[162] = 1'b0;
  assign lce_data_resp_o[163] = 1'b0;
  assign lce_data_resp_o[164] = 1'b0;
  assign lce_data_resp_o[165] = 1'b0;
  assign lce_data_resp_o[166] = 1'b0;
  assign lce_data_resp_o[167] = 1'b0;
  assign lce_data_resp_o[168] = 1'b0;
  assign lce_data_resp_o[169] = 1'b0;
  assign lce_data_resp_o[170] = 1'b0;
  assign lce_data_resp_o[171] = 1'b0;
  assign lce_data_resp_o[172] = 1'b0;
  assign lce_data_resp_o[173] = 1'b0;
  assign lce_data_resp_o[174] = 1'b0;
  assign lce_data_resp_o[175] = 1'b0;
  assign lce_data_resp_o[176] = 1'b0;
  assign lce_data_resp_o[177] = 1'b0;
  assign lce_data_resp_o[178] = 1'b0;
  assign lce_data_resp_o[179] = 1'b0;
  assign lce_data_resp_o[180] = 1'b0;
  assign lce_data_resp_o[181] = 1'b0;
  assign lce_data_resp_o[182] = 1'b0;
  assign lce_data_resp_o[183] = 1'b0;
  assign lce_data_resp_o[184] = 1'b0;
  assign lce_data_resp_o[185] = 1'b0;
  assign lce_data_resp_o[186] = 1'b0;
  assign lce_data_resp_o[187] = 1'b0;
  assign lce_data_resp_o[188] = 1'b0;
  assign lce_data_resp_o[189] = 1'b0;
  assign lce_data_resp_o[190] = 1'b0;
  assign lce_data_resp_o[191] = 1'b0;
  assign lce_data_resp_o[192] = 1'b0;
  assign lce_data_resp_o[193] = 1'b0;
  assign lce_data_resp_o[194] = 1'b0;
  assign lce_data_resp_o[195] = 1'b0;
  assign lce_data_resp_o[196] = 1'b0;
  assign lce_data_resp_o[197] = 1'b0;
  assign lce_data_resp_o[198] = 1'b0;
  assign lce_data_resp_o[199] = 1'b0;
  assign lce_data_resp_o[200] = 1'b0;
  assign lce_data_resp_o[201] = 1'b0;
  assign lce_data_resp_o[202] = 1'b0;
  assign lce_data_resp_o[203] = 1'b0;
  assign lce_data_resp_o[204] = 1'b0;
  assign lce_data_resp_o[205] = 1'b0;
  assign lce_data_resp_o[206] = 1'b0;
  assign lce_data_resp_o[207] = 1'b0;
  assign lce_data_resp_o[208] = 1'b0;
  assign lce_data_resp_o[209] = 1'b0;
  assign lce_data_resp_o[210] = 1'b0;
  assign lce_data_resp_o[211] = 1'b0;
  assign lce_data_resp_o[212] = 1'b0;
  assign lce_data_resp_o[213] = 1'b0;
  assign lce_data_resp_o[214] = 1'b0;
  assign lce_data_resp_o[215] = 1'b0;
  assign lce_data_resp_o[216] = 1'b0;
  assign lce_data_resp_o[217] = 1'b0;
  assign lce_data_resp_o[218] = 1'b0;
  assign lce_data_resp_o[219] = 1'b0;
  assign lce_data_resp_o[220] = 1'b0;
  assign lce_data_resp_o[221] = 1'b0;
  assign lce_data_resp_o[222] = 1'b0;
  assign lce_data_resp_o[223] = 1'b0;
  assign lce_data_resp_o[224] = 1'b0;
  assign lce_data_resp_o[225] = 1'b0;
  assign lce_data_resp_o[226] = 1'b0;
  assign lce_data_resp_o[227] = 1'b0;
  assign lce_data_resp_o[228] = 1'b0;
  assign lce_data_resp_o[229] = 1'b0;
  assign lce_data_resp_o[230] = 1'b0;
  assign lce_data_resp_o[231] = 1'b0;
  assign lce_data_resp_o[232] = 1'b0;
  assign lce_data_resp_o[233] = 1'b0;
  assign lce_data_resp_o[234] = 1'b0;
  assign lce_data_resp_o[235] = 1'b0;
  assign lce_data_resp_o[236] = 1'b0;
  assign lce_data_resp_o[237] = 1'b0;
  assign lce_data_resp_o[238] = 1'b0;
  assign lce_data_resp_o[239] = 1'b0;
  assign lce_data_resp_o[240] = 1'b0;
  assign lce_data_resp_o[241] = 1'b0;
  assign lce_data_resp_o[242] = 1'b0;
  assign lce_data_resp_o[243] = 1'b0;
  assign lce_data_resp_o[244] = 1'b0;
  assign lce_data_resp_o[245] = 1'b0;
  assign lce_data_resp_o[246] = 1'b0;
  assign lce_data_resp_o[247] = 1'b0;
  assign lce_data_resp_o[248] = 1'b0;
  assign lce_data_resp_o[249] = 1'b0;
  assign lce_data_resp_o[250] = 1'b0;
  assign lce_data_resp_o[251] = 1'b0;
  assign lce_data_resp_o[252] = 1'b0;
  assign lce_data_resp_o[253] = 1'b0;
  assign lce_data_resp_o[254] = 1'b0;
  assign lce_data_resp_o[255] = 1'b0;
  assign lce_data_resp_o[256] = 1'b0;
  assign lce_data_resp_o[257] = 1'b0;
  assign lce_data_resp_o[258] = 1'b0;
  assign lce_data_resp_o[259] = 1'b0;
  assign lce_data_resp_o[260] = 1'b0;
  assign lce_data_resp_o[261] = 1'b0;
  assign lce_data_resp_o[262] = 1'b0;
  assign lce_data_resp_o[263] = 1'b0;
  assign lce_data_resp_o[264] = 1'b0;
  assign lce_data_resp_o[265] = 1'b0;
  assign lce_data_resp_o[266] = 1'b0;
  assign lce_data_resp_o[267] = 1'b0;
  assign lce_data_resp_o[268] = 1'b0;
  assign lce_data_resp_o[269] = 1'b0;
  assign lce_data_resp_o[270] = 1'b0;
  assign lce_data_resp_o[271] = 1'b0;
  assign lce_data_resp_o[272] = 1'b0;
  assign lce_data_resp_o[273] = 1'b0;
  assign lce_data_resp_o[274] = 1'b0;
  assign lce_data_resp_o[275] = 1'b0;
  assign lce_data_resp_o[276] = 1'b0;
  assign lce_data_resp_o[277] = 1'b0;
  assign lce_data_resp_o[278] = 1'b0;
  assign lce_data_resp_o[279] = 1'b0;
  assign lce_data_resp_o[280] = 1'b0;
  assign lce_data_resp_o[281] = 1'b0;
  assign lce_data_resp_o[282] = 1'b0;
  assign lce_data_resp_o[283] = 1'b0;
  assign lce_data_resp_o[284] = 1'b0;
  assign lce_data_resp_o[285] = 1'b0;
  assign lce_data_resp_o[286] = 1'b0;
  assign lce_data_resp_o[287] = 1'b0;
  assign lce_data_resp_o[288] = 1'b0;
  assign lce_data_resp_o[289] = 1'b0;
  assign lce_data_resp_o[290] = 1'b0;
  assign lce_data_resp_o[291] = 1'b0;
  assign lce_data_resp_o[292] = 1'b0;
  assign lce_data_resp_o[293] = 1'b0;
  assign lce_data_resp_o[294] = 1'b0;
  assign lce_data_resp_o[295] = 1'b0;
  assign lce_data_resp_o[296] = 1'b0;
  assign lce_data_resp_o[297] = 1'b0;
  assign lce_data_resp_o[298] = 1'b0;
  assign lce_data_resp_o[299] = 1'b0;
  assign lce_data_resp_o[300] = 1'b0;
  assign lce_data_resp_o[301] = 1'b0;
  assign lce_data_resp_o[302] = 1'b0;
  assign lce_data_resp_o[303] = 1'b0;
  assign lce_data_resp_o[304] = 1'b0;
  assign lce_data_resp_o[305] = 1'b0;
  assign lce_data_resp_o[306] = 1'b0;
  assign lce_data_resp_o[307] = 1'b0;
  assign lce_data_resp_o[308] = 1'b0;
  assign lce_data_resp_o[309] = 1'b0;
  assign lce_data_resp_o[310] = 1'b0;
  assign lce_data_resp_o[311] = 1'b0;
  assign lce_data_resp_o[312] = 1'b0;
  assign lce_data_resp_o[313] = 1'b0;
  assign lce_data_resp_o[314] = 1'b0;
  assign lce_data_resp_o[315] = 1'b0;
  assign lce_data_resp_o[316] = 1'b0;
  assign lce_data_resp_o[317] = 1'b0;
  assign lce_data_resp_o[318] = 1'b0;
  assign lce_data_resp_o[319] = 1'b0;
  assign lce_data_resp_o[320] = 1'b0;
  assign lce_data_resp_o[321] = 1'b0;
  assign lce_data_resp_o[322] = 1'b0;
  assign lce_data_resp_o[323] = 1'b0;
  assign lce_data_resp_o[324] = 1'b0;
  assign lce_data_resp_o[325] = 1'b0;
  assign lce_data_resp_o[326] = 1'b0;
  assign lce_data_resp_o[327] = 1'b0;
  assign lce_data_resp_o[328] = 1'b0;
  assign lce_data_resp_o[329] = 1'b0;
  assign lce_data_resp_o[330] = 1'b0;
  assign lce_data_resp_o[331] = 1'b0;
  assign lce_data_resp_o[332] = 1'b0;
  assign lce_data_resp_o[333] = 1'b0;
  assign lce_data_resp_o[334] = 1'b0;
  assign lce_data_resp_o[335] = 1'b0;
  assign lce_data_resp_o[336] = 1'b0;
  assign lce_data_resp_o[337] = 1'b0;
  assign lce_data_resp_o[338] = 1'b0;
  assign lce_data_resp_o[339] = 1'b0;
  assign lce_data_resp_o[340] = 1'b0;
  assign lce_data_resp_o[341] = 1'b0;
  assign lce_data_resp_o[342] = 1'b0;
  assign lce_data_resp_o[343] = 1'b0;
  assign lce_data_resp_o[344] = 1'b0;
  assign lce_data_resp_o[345] = 1'b0;
  assign lce_data_resp_o[346] = 1'b0;
  assign lce_data_resp_o[347] = 1'b0;
  assign lce_data_resp_o[348] = 1'b0;
  assign lce_data_resp_o[349] = 1'b0;
  assign lce_data_resp_o[350] = 1'b0;
  assign lce_data_resp_o[351] = 1'b0;
  assign lce_data_resp_o[352] = 1'b0;
  assign lce_data_resp_o[353] = 1'b0;
  assign lce_data_resp_o[354] = 1'b0;
  assign lce_data_resp_o[355] = 1'b0;
  assign lce_data_resp_o[356] = 1'b0;
  assign lce_data_resp_o[357] = 1'b0;
  assign lce_data_resp_o[358] = 1'b0;
  assign lce_data_resp_o[359] = 1'b0;
  assign lce_data_resp_o[360] = 1'b0;
  assign lce_data_resp_o[361] = 1'b0;
  assign lce_data_resp_o[362] = 1'b0;
  assign lce_data_resp_o[363] = 1'b0;
  assign lce_data_resp_o[364] = 1'b0;
  assign lce_data_resp_o[365] = 1'b0;
  assign lce_data_resp_o[366] = 1'b0;
  assign lce_data_resp_o[367] = 1'b0;
  assign lce_data_resp_o[368] = 1'b0;
  assign lce_data_resp_o[369] = 1'b0;
  assign lce_data_resp_o[370] = 1'b0;
  assign lce_data_resp_o[371] = 1'b0;
  assign lce_data_resp_o[372] = 1'b0;
  assign lce_data_resp_o[373] = 1'b0;
  assign lce_data_resp_o[374] = 1'b0;
  assign lce_data_resp_o[375] = 1'b0;
  assign lce_data_resp_o[376] = 1'b0;
  assign lce_data_resp_o[377] = 1'b0;
  assign lce_data_resp_o[378] = 1'b0;
  assign lce_data_resp_o[379] = 1'b0;
  assign lce_data_resp_o[380] = 1'b0;
  assign lce_data_resp_o[381] = 1'b0;
  assign lce_data_resp_o[382] = 1'b0;
  assign lce_data_resp_o[383] = 1'b0;
  assign lce_data_resp_o[384] = 1'b0;
  assign lce_data_resp_o[385] = 1'b0;
  assign lce_data_resp_o[386] = 1'b0;
  assign lce_data_resp_o[387] = 1'b0;
  assign lce_data_resp_o[388] = 1'b0;
  assign lce_data_resp_o[389] = 1'b0;
  assign lce_data_resp_o[390] = 1'b0;
  assign lce_data_resp_o[391] = 1'b0;
  assign lce_data_resp_o[392] = 1'b0;
  assign lce_data_resp_o[393] = 1'b0;
  assign lce_data_resp_o[394] = 1'b0;
  assign lce_data_resp_o[395] = 1'b0;
  assign lce_data_resp_o[396] = 1'b0;
  assign lce_data_resp_o[397] = 1'b0;
  assign lce_data_resp_o[398] = 1'b0;
  assign lce_data_resp_o[399] = 1'b0;
  assign lce_data_resp_o[400] = 1'b0;
  assign lce_data_resp_o[401] = 1'b0;
  assign lce_data_resp_o[402] = 1'b0;
  assign lce_data_resp_o[403] = 1'b0;
  assign lce_data_resp_o[404] = 1'b0;
  assign lce_data_resp_o[405] = 1'b0;
  assign lce_data_resp_o[406] = 1'b0;
  assign lce_data_resp_o[407] = 1'b0;
  assign lce_data_resp_o[408] = 1'b0;
  assign lce_data_resp_o[409] = 1'b0;
  assign lce_data_resp_o[410] = 1'b0;
  assign lce_data_resp_o[411] = 1'b0;
  assign lce_data_resp_o[412] = 1'b0;
  assign lce_data_resp_o[413] = 1'b0;
  assign lce_data_resp_o[414] = 1'b0;
  assign lce_data_resp_o[415] = 1'b0;
  assign lce_data_resp_o[416] = 1'b0;
  assign lce_data_resp_o[417] = 1'b0;
  assign lce_data_resp_o[418] = 1'b0;
  assign lce_data_resp_o[419] = 1'b0;
  assign lce_data_resp_o[420] = 1'b0;
  assign lce_data_resp_o[421] = 1'b0;
  assign lce_data_resp_o[422] = 1'b0;
  assign lce_data_resp_o[423] = 1'b0;
  assign lce_data_resp_o[424] = 1'b0;
  assign lce_data_resp_o[425] = 1'b0;
  assign lce_data_resp_o[426] = 1'b0;
  assign lce_data_resp_o[427] = 1'b0;
  assign lce_data_resp_o[428] = 1'b0;
  assign lce_data_resp_o[429] = 1'b0;
  assign lce_data_resp_o[430] = 1'b0;
  assign lce_data_resp_o[431] = 1'b0;
  assign lce_data_resp_o[432] = 1'b0;
  assign lce_data_resp_o[433] = 1'b0;
  assign lce_data_resp_o[434] = 1'b0;
  assign lce_data_resp_o[435] = 1'b0;
  assign lce_data_resp_o[436] = 1'b0;
  assign lce_data_resp_o[437] = 1'b0;
  assign lce_data_resp_o[438] = 1'b0;
  assign lce_data_resp_o[439] = 1'b0;
  assign lce_data_resp_o[440] = 1'b0;
  assign lce_data_resp_o[441] = 1'b0;
  assign lce_data_resp_o[442] = 1'b0;
  assign lce_data_resp_o[443] = 1'b0;
  assign lce_data_resp_o[444] = 1'b0;
  assign lce_data_resp_o[445] = 1'b0;
  assign lce_data_resp_o[446] = 1'b0;
  assign lce_data_resp_o[447] = 1'b0;
  assign lce_data_resp_o[448] = 1'b0;
  assign lce_data_resp_o[449] = 1'b0;
  assign lce_data_resp_o[450] = 1'b0;
  assign lce_data_resp_o[451] = 1'b0;
  assign lce_data_resp_o[452] = 1'b0;
  assign lce_data_resp_o[453] = 1'b0;
  assign lce_data_resp_o[454] = 1'b0;
  assign lce_data_resp_o[455] = 1'b0;
  assign lce_data_resp_o[456] = 1'b0;
  assign lce_data_resp_o[457] = 1'b0;
  assign lce_data_resp_o[458] = 1'b0;
  assign lce_data_resp_o[459] = 1'b0;
  assign lce_data_resp_o[460] = 1'b0;
  assign lce_data_resp_o[461] = 1'b0;
  assign lce_data_resp_o[462] = 1'b0;
  assign lce_data_resp_o[463] = 1'b0;
  assign lce_data_resp_o[464] = 1'b0;
  assign lce_data_resp_o[465] = 1'b0;
  assign lce_data_resp_o[466] = 1'b0;
  assign lce_data_resp_o[467] = 1'b0;
  assign lce_data_resp_o[468] = 1'b0;
  assign lce_data_resp_o[469] = 1'b0;
  assign lce_data_resp_o[470] = 1'b0;
  assign lce_data_resp_o[471] = 1'b0;
  assign lce_data_resp_o[472] = 1'b0;
  assign lce_data_resp_o[473] = 1'b0;
  assign lce_data_resp_o[474] = 1'b0;
  assign lce_data_resp_o[475] = 1'b0;
  assign lce_data_resp_o[476] = 1'b0;
  assign lce_data_resp_o[477] = 1'b0;
  assign lce_data_resp_o[478] = 1'b0;
  assign lce_data_resp_o[479] = 1'b0;
  assign lce_data_resp_o[480] = 1'b0;
  assign lce_data_resp_o[481] = 1'b0;
  assign lce_data_resp_o[482] = 1'b0;
  assign lce_data_resp_o[483] = 1'b0;
  assign lce_data_resp_o[484] = 1'b0;
  assign lce_data_resp_o[485] = 1'b0;
  assign lce_data_resp_o[486] = 1'b0;
  assign lce_data_resp_o[487] = 1'b0;
  assign lce_data_resp_o[488] = 1'b0;
  assign lce_data_resp_o[489] = 1'b0;
  assign lce_data_resp_o[490] = 1'b0;
  assign lce_data_resp_o[491] = 1'b0;
  assign lce_data_resp_o[492] = 1'b0;
  assign lce_data_resp_o[493] = 1'b0;
  assign lce_data_resp_o[494] = 1'b0;
  assign lce_data_resp_o[495] = 1'b0;
  assign lce_data_resp_o[496] = 1'b0;
  assign lce_data_resp_o[497] = 1'b0;
  assign lce_data_resp_o[498] = 1'b0;
  assign lce_data_resp_o[499] = 1'b0;
  assign lce_data_resp_o[500] = 1'b0;
  assign lce_data_resp_o[501] = 1'b0;
  assign lce_data_resp_o[502] = 1'b0;
  assign lce_data_resp_o[503] = 1'b0;
  assign lce_data_resp_o[504] = 1'b0;
  assign lce_data_resp_o[505] = 1'b0;
  assign lce_data_resp_o[506] = 1'b0;
  assign lce_data_resp_o[507] = 1'b0;
  assign lce_data_resp_o[508] = 1'b0;
  assign lce_data_resp_o[509] = 1'b0;
  assign lce_data_resp_o[510] = 1'b0;
  assign lce_data_resp_o[511] = 1'b0;
  assign lce_data_resp_o[512] = 1'b0;
  assign lce_data_resp_o[513] = 1'b0;
  assign lce_data_resp_o[514] = 1'b0;
  assign lce_data_resp_o[515] = 1'b0;
  assign lce_data_resp_o[516] = 1'b0;
  assign lce_data_resp_o[517] = 1'b0;
  assign lce_data_resp_o[518] = 1'b0;
  assign lce_data_resp_o[519] = 1'b0;
  assign lce_data_resp_o[520] = 1'b0;
  assign lce_data_resp_o[521] = 1'b0;
  assign lce_data_resp_o[522] = 1'b0;
  assign lce_data_resp_o[523] = 1'b0;
  assign lce_data_resp_o[524] = 1'b0;
  assign lce_data_resp_o[525] = 1'b0;
  assign lce_data_resp_o[526] = 1'b0;
  assign lce_data_resp_o[527] = 1'b0;
  assign lce_data_resp_o[528] = 1'b0;
  assign lce_data_resp_o[529] = 1'b0;
  assign lce_data_resp_o[530] = 1'b0;
  assign lce_data_resp_o[531] = 1'b0;
  assign lce_data_resp_o[532] = 1'b0;
  assign lce_data_resp_o[533] = 1'b0;
  assign lce_data_resp_o[534] = 1'b0;
  assign lce_data_resp_o[535] = 1'b0;
  assign lce_data_resp_o[536] = 1'b0;
  assign lce_data_resp_o[537] = 1'b0;
  assign lce_data_resp_o[538] = 1'b0;
  assign lce_data_resp_o[539] = 1'b0;
  assign lce_data_resp_o[540] = 1'b0;
  assign lce_data_resp_o[541] = 1'b0;
  assign lce_data_resp_o[542] = 1'b0;
  assign lce_data_resp_o[543] = 1'b0;
  assign lce_data_resp_o[544] = 1'b0;
  assign lce_data_resp_o[545] = 1'b0;
  assign lce_data_resp_o[546] = 1'b0;
  assign lce_data_resp_o[547] = 1'b0;
  assign lce_data_resp_o[548] = 1'b0;
  assign lce_data_resp_o[549] = 1'b0;
  assign lce_data_resp_o[550] = 1'b0;
  assign lce_data_resp_o[551] = 1'b0;
  assign lce_data_resp_o[552] = 1'b0;
  assign lce_data_resp_o[553] = 1'b0;
  assign lce_resp_o[40] = 1'b0;
  assign lce_data_resp_o[40] = id_i[0];
  assign lce_resp_o[41] = id_i[0];
  assign N23 = state_r[1] | N22;
  assign N26 = N25 | state_r[0];
  assign N28 = N25 & N22;
  assign N29 = state_r[1] & state_r[0];

  bsg_two_fifo_width_p53
  rv_adapter
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(lce_cmd_ready_o),
    .data_i(lce_cmd_i),
    .v_i(lce_cmd_v_i),
    .v_o(lce_cmd_v_li),
    .data_o({ lce_cmd_li_dst_id__0_, lce_cmd_li_src_id__0_, lce_cmd_li_msg_type__2_, lce_cmd_li_msg_type__1_, lce_cmd_li_msg_type__0_, lce_cmd_addr_tag, lce_cmd_addr_index, lce_cmd_li_addr__5_, lce_cmd_li_addr__4_, lce_cmd_li_addr__3_, lce_cmd_li_addr__2_, lce_cmd_li_addr__1_, lce_cmd_li_addr__0_, lce_cmd_li_way_id__2_, lce_cmd_li_way_id__1_, lce_cmd_li_way_id__0_, lce_cmd_li_state__1_, lce_cmd_li_state__0_, lce_cmd_li_target__0_, lce_cmd_li_target_way_id__2_, lce_cmd_li_target_way_id__1_, lce_cmd_li_target_way_id__0_ }),
    .yumi_i(lce_cmd_yumi_lo)
  );

  assign lce_ready_o = state_r[0] | state_r[1];
  assign N835 = ~lce_cmd_li_msg_type__0_;
  assign N836 = lce_cmd_li_msg_type__1_ | lce_cmd_li_msg_type__2_;
  assign N837 = N835 | N836;
  assign N838 = ~N837;
  assign N839 = ~lce_cmd_li_msg_type__2_;
  assign N840 = ~lce_cmd_li_msg_type__1_;
  assign N841 = N840 | N839;
  assign N842 = lce_cmd_li_msg_type__0_ | N841;
  assign N843 = ~N842;
  assign N844 = ~syn_ack_cnt_r[0];
  assign N845 = lce_cmd_li_msg_type__1_ | N839;
  assign N846 = N835 | N845;
  assign N847 = ~N846;
  assign N848 = lce_cmd_li_msg_type__1_ | lce_cmd_li_msg_type__2_;
  assign N849 = lce_cmd_li_msg_type__0_ | N848;
  assign N850 = ~N849;
  assign N851 = lce_cmd_li_msg_type__1_ | N839;
  assign N852 = lce_cmd_li_msg_type__0_ | N851;
  assign N853 = ~N852;
  assign N854 = N840 | lce_cmd_li_msg_type__2_;
  assign N855 = N835 | N854;
  assign N856 = ~N855;
  assign N857 = N840 | lce_cmd_li_msg_type__2_;
  assign N858 = lce_cmd_li_msg_type__0_ | N857;
  assign N859 = ~N858;
  assign N705 = syn_ack_cnt_r[0] ^ 1'b1;
  assign N38 = (N0)? 1'b0 : 
               (N1)? lce_cmd_v_li : 1'b0;
  assign N0 = flag_invalidate_r;
  assign N1 = N37;
  assign N41 = (N2)? 1'b0 : 
               (N729)? 1'b1 : 
               (N40)? tag_mem_pkt_yumi_i : 1'b0;
  assign N2 = lce_resp_yumi_i;
  assign { N52, N51, N50, N49, N48, N47, N46, N45, N44, N43 } = (N3)? { lce_cmd_addr_index, lce_cmd_li_way_id__2_, lce_cmd_li_way_id__1_, lce_cmd_li_way_id__0_, 1'b1 } : 
                                                                (N4)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N3 = N859;
  assign N4 = N858;
  assign N5 = 1'b0;
  assign N53 = (N3)? lce_cmd_v_li : 
               (N4)? 1'b0 : 
               (N5)? 1'b0 : 
               (N5)? 1'b0 : 
               (N5)? 1'b0 : 
               (N5)? 1'b0 : 1'b0;
  assign { N55, N54 } = (N3)? { data_mem_pkt_yumi_i, N35 } : 
                        (N4)? state_r : 1'b0;
  assign { N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57 } = (N3)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                           (N6)? { lce_cmd_li_src_id__0_, 1'b1, lce_cmd_addr_tag, lce_cmd_addr_index, lce_cmd_li_addr__5_, lce_cmd_li_addr__4_, lce_cmd_li_addr__3_, lce_cmd_li_addr__2_, lce_cmd_li_addr__1_, lce_cmd_li_addr__0_ } : 
                                                                                                                                                                                                                           (N56)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                           (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                           (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                           (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N6 = N856;
  assign N98 = (N3)? 1'b0 : 
               (N6)? lce_cmd_v_li : 
               (N56)? 1'b0 : 
               (N5)? 1'b0 : 
               (N5)? 1'b0 : 
               (N5)? 1'b0 : 1'b0;
  assign N99 = (N3)? 1'b0 : 
               (N6)? N36 : 
               (N7)? tag_mem_pkt_yumi_i : 
               (N8)? tag_mem_pkt_yumi_i : 
               (N9)? lce_resp_yumi_i : 
               (N34)? 1'b0 : 1'b0;
  assign N7 = N853;
  assign N8 = N847;
  assign N9 = N843;
  assign { N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101 } = (N3)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                  (N6)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                  (N7)? { lce_cmd_li_state__1_, lce_cmd_li_state__0_, lce_cmd_addr_tag, 1'b1 } : 
                                                                                                                                                                                                  (N8)? { lce_cmd_li_state__1_, lce_cmd_li_state__0_, lce_cmd_addr_tag, 1'b1 } : 
                                                                                                                                                                                                  (N100)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                  (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { N139, N138, N137, N136, N135, N134, N133, N132, N131 } = (N3)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                    (N6)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                    (N7)? { lce_cmd_addr_index, lce_cmd_li_way_id__2_, lce_cmd_li_way_id__1_, lce_cmd_li_way_id__0_ } : 
                                                                    (N8)? { lce_cmd_addr_index, lce_cmd_li_way_id__2_, lce_cmd_li_way_id__1_, lce_cmd_li_way_id__0_ } : 
                                                                    (N9)? { lce_cmd_addr_index, lce_cmd_li_way_id__2_, lce_cmd_li_way_id__1_, lce_cmd_li_way_id__0_ } : 
                                                                    (N34)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N140 = (N3)? 1'b0 : 
                (N6)? 1'b0 : 
                (N7)? lce_cmd_v_li : 
                (N8)? lce_cmd_v_li : 
                (N9)? N38 : 
                (N34)? 1'b0 : 1'b0;
  assign N142 = (N3)? 1'b0 : 
                (N6)? 1'b0 : 
                (N7)? tag_mem_pkt_yumi_i : 
                (N141)? 1'b0 : 
                (N5)? 1'b0 : 
                (N5)? 1'b0 : 1'b0;
  assign N143 = (N3)? 1'b0 : 
                (N6)? 1'b0 : 
                (N7)? 1'b0 : 
                (N8)? tag_mem_pkt_yumi_i : 
                (N100)? 1'b0 : 
                (N5)? 1'b0 : 1'b0;
  assign N144 = (N3)? flag_invalidate_r : 
                (N6)? flag_invalidate_r : 
                (N7)? flag_invalidate_r : 
                (N8)? flag_invalidate_r : 
                (N9)? N41 : 
                (N34)? flag_invalidate_r : 1'b0;
  assign { N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145 } = (N3)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                    (N6)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                    (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                    (N8)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                    (N9)? { lce_cmd_li_src_id__0_, 1'b1, lce_cmd_addr_tag, lce_cmd_addr_index, lce_cmd_li_addr__5_, lce_cmd_li_addr__4_, lce_cmd_li_addr__3_, lce_cmd_li_addr__2_, lce_cmd_li_addr__1_, lce_cmd_li_addr__0_ } : 
                                                                                                                                                                                                                                                                    (N34)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N186 = (N3)? 1'b0 : 
                (N6)? 1'b0 : 
                (N7)? 1'b0 : 
                (N8)? 1'b0 : 
                (N9)? N42 : 
                (N34)? 1'b0 : 1'b0;
  assign { N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189 } = (N10)? data_r : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N11)? data_mem_data_i : 1'b0;
  assign N10 = flag_data_buffered_r;
  assign N11 = N188;
  assign N706 = (N2)? N705 : 
                (N12)? syn_ack_cnt_r[0] : 1'b0;
  assign N12 = N704;
  assign { N713, N712, N711, N710, N709, N708 } = (N13)? lce_cmd_addr_index : 
                                                  (N14)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                  (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N13 = N838;
  assign N14 = N837;
  assign N714 = (N13)? lce_cmd_v_li : 
                (N14)? 1'b0 : 
                (N5)? 1'b0 : 1'b0;
  assign { N720, N719, N718, N717, N716, N715 } = (N13)? lce_cmd_addr_index : 
                                                  (N14)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                  (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N721 = (N13)? lce_cmd_v_li : 
                (N14)? 1'b0 : 
                (N5)? 1'b0 : 1'b0;
  assign N722 = (N13)? N703 : 
                (N15)? lce_resp_yumi_i : 
                (N702)? 1'b0 : 1'b0;
  assign N15 = N850;
  assign N723 = (N13)? 1'b0 : 
                (N15)? lce_cmd_li_src_id__0_ : 
                (N702)? 1'b0 : 1'b0;
  assign N724 = (N13)? 1'b0 : 
                (N15)? lce_cmd_v_li : 
                (N702)? 1'b0 : 1'b0;
  assign N725 = (N13)? syn_ack_cnt_r[0] : 
                (N15)? N706 : 
                (N702)? syn_ack_cnt_r[0] : 1'b0;
  assign { N727, N726 } = (N13)? state_r : 
                          (N15)? { 1'b0, N707 } : 
                          (N702)? state_r : 1'b0;
  assign lce_resp_v_o = (N16)? N186 : 
                        (N17)? 1'b0 : 
                        (N18)? N724 : 
                        (N19)? 1'b0 : 1'b0;
  assign N16 = N24;
  assign N17 = N27;
  assign N18 = N28;
  assign N19 = N29;
  assign { data_mem_pkt_o[522:514], data_mem_pkt_o[0:0] } = (N16)? { N52, N51, N50, N49, N48, N47, N46, N45, N44, N43 } : 
                                                            (N17)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                            (N18)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                            (N19)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign data_mem_pkt_v_o = (N16)? N53 : 
                            (N17)? 1'b0 : 
                            (N18)? 1'b0 : 
                            (N19)? 1'b0 : 1'b0;
  assign state_n = (N16)? { N55, N54 } : 
                   (N17)? { N187, lce_data_cmd_ready_i } : 
                   (N18)? { N727, N726 } : 1'b0;
  assign { lce_data_resp_o[41:41], lce_data_resp_o[39:0] } = (N16)? { N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57 } : 
                                                             (N17)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                             (N18)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                             (N19)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign lce_data_resp_v_o = (N16)? N98 : 
                             (N17)? 1'b0 : 
                             (N18)? 1'b0 : 
                             (N19)? 1'b0 : 1'b0;
  assign lce_cmd_yumi_lo = (N16)? N99 : 
                           (N17)? lce_data_cmd_ready_i : 
                           (N18)? N722 : 
                           (N19)? 1'b0 : 1'b0;
  assign tag_mem_pkt_o = (N16)? { N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N843 } : 
                         (N17)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                         (N18)? { N713, N712, N711, N710, N709, N708, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                         (N19)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign tag_mem_pkt_v_o = (N16)? N140 : 
                           (N17)? 1'b0 : 
                           (N18)? N714 : 
                           (N19)? 1'b0 : 1'b0;
  assign set_tag_received_o = (N16)? N142 : 
                              (N17)? 1'b0 : 
                              (N18)? 1'b0 : 
                              (N19)? 1'b0 : 1'b0;
  assign set_tag_wakeup_received_o = (N16)? N143 : 
                                     (N17)? 1'b0 : 
                                     (N18)? 1'b0 : 
                                     (N19)? 1'b0 : 1'b0;
  assign { lce_resp_o[42:42], lce_resp_o[39:0] } = (N16)? { N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145 } : 
                                                   (N17)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                   (N18)? { N723, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                   (N19)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { lce_data_cmd_o[517:5], lce_data_cmd_o[2:0] } = (N16)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                          (N17)? { N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, lce_cmd_li_target__0_, lce_cmd_li_target_way_id__2_, lce_cmd_li_target_way_id__1_, lce_cmd_li_target_way_id__0_ } : 
                                                          (N18)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                          (N19)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign lce_data_cmd_v_o = (N16)? 1'b0 : 
                            (N17)? 1'b1 : 
                            (N18)? 1'b0 : 
                            (N19)? 1'b0 : 1'b0;
  assign stat_mem_pkt_o[9:4] = (N16)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                               (N17)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                               (N18)? { N720, N719, N718, N717, N716, N715 } : 
                               (N19)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign stat_mem_pkt_v_o = (N16)? 1'b0 : 
                            (N17)? 1'b0 : 
                            (N18)? N721 : 
                            (N19)? 1'b0 : 1'b0;
  assign { N733, N732 } = (N20)? { 1'b0, 1'b0 } : 
                          (N21)? state_n : 1'b0;
  assign N20 = N731;
  assign N21 = N730;
  assign N734 = (N20)? 1'b0 : 
                (N21)? N725 : 1'b0;
  assign N735 = (N20)? 1'b0 : 
                (N21)? N187 : 1'b0;
  assign N736 = (N20)? 1'b0 : 
                (N21)? N144 : 1'b0;
  assign N22 = ~state_r[0];
  assign N24 = ~N23;
  assign N25 = ~state_r[1];
  assign N27 = ~N26;
  assign N30 = N856 | N859;
  assign N31 = N853 | N30;
  assign N32 = N847 | N31;
  assign N33 = N843 | N32;
  assign N34 = ~N33;
  assign N35 = ~data_mem_pkt_yumi_i;
  assign N36 = lce_data_resp_ready_i & lce_cmd_v_li;
  assign N37 = ~flag_invalidate_r;
  assign N39 = flag_invalidate_r | lce_resp_yumi_i;
  assign N40 = ~N39;
  assign N42 = flag_invalidate_r | tag_mem_pkt_yumi_i;
  assign N56 = ~N30;
  assign N100 = ~N32;
  assign N141 = ~N31;
  assign N187 = ~lce_data_cmd_ready_i;
  assign N188 = ~flag_data_buffered_r;
  assign N701 = N850 | N838;
  assign N702 = ~N701;
  assign N703 = tag_mem_pkt_yumi_i & stat_mem_pkt_yumi_i;
  assign N704 = ~lce_resp_yumi_i;
  assign N707 = N844 & lce_resp_yumi_i;
  assign N728 = ~lce_resp_yumi_i;
  assign N729 = flag_invalidate_r & N728;
  assign N730 = ~reset_i;
  assign N731 = reset_i;
  assign N737 = N24 & N730;
  assign N738 = N27 & N730;
  assign N739 = flag_data_buffered_r & N738;
  assign N740 = N737 | N739;
  assign N741 = N28 & N730;
  assign N742 = N740 | N741;
  assign N743 = N29 & N730;
  assign N744 = N742 | N743;
  assign N745 = ~N744;
  assign N746 = N730 & N745;
  assign N747 = N24 & N730;
  assign N748 = N27 & N730;
  assign N749 = flag_data_buffered_r & N748;
  assign N750 = N747 | N749;
  assign N751 = N28 & N730;
  assign N752 = N750 | N751;
  assign N753 = N29 & N730;
  assign N754 = N752 | N753;
  assign N755 = ~N754;
  assign N756 = N730 & N755;
  assign N757 = N24 & N730;
  assign N758 = N27 & N730;
  assign N759 = flag_data_buffered_r & N758;
  assign N760 = N757 | N759;
  assign N761 = N28 & N730;
  assign N762 = N760 | N761;
  assign N763 = N29 & N730;
  assign N764 = N762 | N763;
  assign N765 = ~N764;
  assign N766 = N730 & N765;
  assign N767 = N24 & N730;
  assign N768 = N27 & N730;
  assign N769 = flag_data_buffered_r & N768;
  assign N770 = N767 | N769;
  assign N771 = N28 & N730;
  assign N772 = N770 | N771;
  assign N773 = N29 & N730;
  assign N774 = N772 | N773;
  assign N775 = ~N774;
  assign N776 = N730 & N775;
  assign N777 = N24 & N730;
  assign N778 = N27 & N730;
  assign N779 = flag_data_buffered_r & N778;
  assign N780 = N777 | N779;
  assign N781 = N28 & N730;
  assign N782 = N780 | N781;
  assign N783 = N29 & N730;
  assign N784 = N782 | N783;
  assign N785 = ~N784;
  assign N786 = N730 & N785;
  assign N787 = N24 & N730;
  assign N788 = N27 & N730;
  assign N789 = flag_data_buffered_r & N788;
  assign N790 = N787 | N789;
  assign N791 = N28 & N730;
  assign N792 = N790 | N791;
  assign N793 = N29 & N730;
  assign N794 = N792 | N793;
  assign N795 = ~N794;
  assign N796 = N730 & N795;
  assign N797 = N782 | N793;
  assign N798 = ~N797;
  assign N799 = N730 & N798;
  assign N800 = N730 & N785;
  assign N801 = N772 | N783;
  assign N802 = ~N801;
  assign N803 = N730 & N802;
  assign N804 = N730 & N775;
  assign N805 = N730 & N775;
  assign N806 = N762 | N773;
  assign N807 = ~N806;
  assign N808 = N730 & N807;
  assign N809 = N730 & N765;
  assign N810 = N730 & N765;
  assign N811 = N752 | N763;
  assign N812 = ~N811;
  assign N813 = N730 & N812;
  assign N814 = N730 & N755;
  assign N815 = N730 & N755;
  assign N816 = N742 | N753;
  assign N817 = ~N816;
  assign N818 = N730 & N817;
  assign N819 = N730 & N745;
  assign N820 = N730 & N745;
  assign N821 = N730 & N745;
  assign N822 = N730 & N745;
  assign N823 = N730 & N745;
  assign N824 = ~N743;
  assign N825 = N737 | N738;
  assign N826 = N825 | N743;
  assign N827 = ~N826;
  assign N828 = N737 | N741;
  assign N829 = N828 | N743;
  assign N830 = ~N829;
  assign N831 = N738 | N741;
  assign N832 = N831 | N743;
  assign N833 = ~N832;

  always @(posedge clk_i) begin
    if(N746) begin
      { data_r[511:511], data_r[0:0] } <= { data_mem_data_i[511:511], data_mem_data_i[0:0] };
    end 
    if(N756) begin
      { data_r[510:510] } <= { data_mem_data_i[510:510] };
    end 
    if(N766) begin
      { data_r[509:509] } <= { data_mem_data_i[509:509] };
    end 
    if(N776) begin
      { data_r[508:508] } <= { data_mem_data_i[508:508] };
    end 
    if(N786) begin
      { data_r[507:507], data_r[489:413] } <= { data_mem_data_i[507:507], data_mem_data_i[489:413] };
    end 
    if(N796) begin
      { data_r[506:493] } <= { data_mem_data_i[506:493] };
    end 
    if(N799) begin
      { data_r[492:490] } <= { data_mem_data_i[492:490] };
    end 
    if(N800) begin
      { data_r[412:394] } <= { data_mem_data_i[412:394] };
    end 
    if(N803) begin
      { data_r[393:391] } <= { data_mem_data_i[393:391] };
    end 
    if(N804) begin
      { data_r[390:314] } <= { data_mem_data_i[390:314] };
    end 
    if(N805) begin
      { data_r[313:295] } <= { data_mem_data_i[313:295] };
    end 
    if(N808) begin
      { data_r[294:292] } <= { data_mem_data_i[294:292] };
    end 
    if(N809) begin
      { data_r[291:215] } <= { data_mem_data_i[291:215] };
    end 
    if(N810) begin
      { data_r[214:196] } <= { data_mem_data_i[214:196] };
    end 
    if(N813) begin
      { data_r[195:193] } <= { data_mem_data_i[195:193] };
    end 
    if(N814) begin
      { data_r[192:116] } <= { data_mem_data_i[192:116] };
    end 
    if(N815) begin
      { data_r[115:97] } <= { data_mem_data_i[115:97] };
    end 
    if(N818) begin
      { data_r[96:94] } <= { data_mem_data_i[96:94] };
    end 
    if(N819) begin
      { data_r[93:17], data_r[4:4] } <= { data_mem_data_i[93:17], data_mem_data_i[4:4] };
    end 
    if(N820) begin
      { data_r[16:5] } <= { data_mem_data_i[16:5] };
    end 
    if(N821) begin
      { data_r[3:3] } <= { data_mem_data_i[3:3] };
    end 
    if(N822) begin
      { data_r[2:2] } <= { data_mem_data_i[2:2] };
    end 
    if(N823) begin
      { data_r[1:1] } <= { data_mem_data_i[1:1] };
    end 
    if(N824) begin
      { state_r[1:0] } <= { N733, N732 };
    end 
    if(N827) begin
      { syn_ack_cnt_r[0:0] } <= { N734 };
    end 
    if(N830) begin
      flag_data_buffered_r <= N735;
    end 
    if(N833) begin
      flag_invalidate_r <= N736;
    end 
  end


endmodule



module bsg_mem_1r1w_synth_width_p518_els_p2_read_write_same_addr_p0_harden_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [517:0] w_data_i;
  input [0:0] r_addr_i;
  output [517:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [517:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18;
  reg [1035:0] mem;
  assign r_data_o[517] = (N3)? mem[517] : 
                         (N0)? mem[1035] : 1'b0;
  assign N0 = r_addr_i[0];
  assign r_data_o[516] = (N3)? mem[516] : 
                         (N0)? mem[1034] : 1'b0;
  assign r_data_o[515] = (N3)? mem[515] : 
                         (N0)? mem[1033] : 1'b0;
  assign r_data_o[514] = (N3)? mem[514] : 
                         (N0)? mem[1032] : 1'b0;
  assign r_data_o[513] = (N3)? mem[513] : 
                         (N0)? mem[1031] : 1'b0;
  assign r_data_o[512] = (N3)? mem[512] : 
                         (N0)? mem[1030] : 1'b0;
  assign r_data_o[511] = (N3)? mem[511] : 
                         (N0)? mem[1029] : 1'b0;
  assign r_data_o[510] = (N3)? mem[510] : 
                         (N0)? mem[1028] : 1'b0;
  assign r_data_o[509] = (N3)? mem[509] : 
                         (N0)? mem[1027] : 1'b0;
  assign r_data_o[508] = (N3)? mem[508] : 
                         (N0)? mem[1026] : 1'b0;
  assign r_data_o[507] = (N3)? mem[507] : 
                         (N0)? mem[1025] : 1'b0;
  assign r_data_o[506] = (N3)? mem[506] : 
                         (N0)? mem[1024] : 1'b0;
  assign r_data_o[505] = (N3)? mem[505] : 
                         (N0)? mem[1023] : 1'b0;
  assign r_data_o[504] = (N3)? mem[504] : 
                         (N0)? mem[1022] : 1'b0;
  assign r_data_o[503] = (N3)? mem[503] : 
                         (N0)? mem[1021] : 1'b0;
  assign r_data_o[502] = (N3)? mem[502] : 
                         (N0)? mem[1020] : 1'b0;
  assign r_data_o[501] = (N3)? mem[501] : 
                         (N0)? mem[1019] : 1'b0;
  assign r_data_o[500] = (N3)? mem[500] : 
                         (N0)? mem[1018] : 1'b0;
  assign r_data_o[499] = (N3)? mem[499] : 
                         (N0)? mem[1017] : 1'b0;
  assign r_data_o[498] = (N3)? mem[498] : 
                         (N0)? mem[1016] : 1'b0;
  assign r_data_o[497] = (N3)? mem[497] : 
                         (N0)? mem[1015] : 1'b0;
  assign r_data_o[496] = (N3)? mem[496] : 
                         (N0)? mem[1014] : 1'b0;
  assign r_data_o[495] = (N3)? mem[495] : 
                         (N0)? mem[1013] : 1'b0;
  assign r_data_o[494] = (N3)? mem[494] : 
                         (N0)? mem[1012] : 1'b0;
  assign r_data_o[493] = (N3)? mem[493] : 
                         (N0)? mem[1011] : 1'b0;
  assign r_data_o[492] = (N3)? mem[492] : 
                         (N0)? mem[1010] : 1'b0;
  assign r_data_o[491] = (N3)? mem[491] : 
                         (N0)? mem[1009] : 1'b0;
  assign r_data_o[490] = (N3)? mem[490] : 
                         (N0)? mem[1008] : 1'b0;
  assign r_data_o[489] = (N3)? mem[489] : 
                         (N0)? mem[1007] : 1'b0;
  assign r_data_o[488] = (N3)? mem[488] : 
                         (N0)? mem[1006] : 1'b0;
  assign r_data_o[487] = (N3)? mem[487] : 
                         (N0)? mem[1005] : 1'b0;
  assign r_data_o[486] = (N3)? mem[486] : 
                         (N0)? mem[1004] : 1'b0;
  assign r_data_o[485] = (N3)? mem[485] : 
                         (N0)? mem[1003] : 1'b0;
  assign r_data_o[484] = (N3)? mem[484] : 
                         (N0)? mem[1002] : 1'b0;
  assign r_data_o[483] = (N3)? mem[483] : 
                         (N0)? mem[1001] : 1'b0;
  assign r_data_o[482] = (N3)? mem[482] : 
                         (N0)? mem[1000] : 1'b0;
  assign r_data_o[481] = (N3)? mem[481] : 
                         (N0)? mem[999] : 1'b0;
  assign r_data_o[480] = (N3)? mem[480] : 
                         (N0)? mem[998] : 1'b0;
  assign r_data_o[479] = (N3)? mem[479] : 
                         (N0)? mem[997] : 1'b0;
  assign r_data_o[478] = (N3)? mem[478] : 
                         (N0)? mem[996] : 1'b0;
  assign r_data_o[477] = (N3)? mem[477] : 
                         (N0)? mem[995] : 1'b0;
  assign r_data_o[476] = (N3)? mem[476] : 
                         (N0)? mem[994] : 1'b0;
  assign r_data_o[475] = (N3)? mem[475] : 
                         (N0)? mem[993] : 1'b0;
  assign r_data_o[474] = (N3)? mem[474] : 
                         (N0)? mem[992] : 1'b0;
  assign r_data_o[473] = (N3)? mem[473] : 
                         (N0)? mem[991] : 1'b0;
  assign r_data_o[472] = (N3)? mem[472] : 
                         (N0)? mem[990] : 1'b0;
  assign r_data_o[471] = (N3)? mem[471] : 
                         (N0)? mem[989] : 1'b0;
  assign r_data_o[470] = (N3)? mem[470] : 
                         (N0)? mem[988] : 1'b0;
  assign r_data_o[469] = (N3)? mem[469] : 
                         (N0)? mem[987] : 1'b0;
  assign r_data_o[468] = (N3)? mem[468] : 
                         (N0)? mem[986] : 1'b0;
  assign r_data_o[467] = (N3)? mem[467] : 
                         (N0)? mem[985] : 1'b0;
  assign r_data_o[466] = (N3)? mem[466] : 
                         (N0)? mem[984] : 1'b0;
  assign r_data_o[465] = (N3)? mem[465] : 
                         (N0)? mem[983] : 1'b0;
  assign r_data_o[464] = (N3)? mem[464] : 
                         (N0)? mem[982] : 1'b0;
  assign r_data_o[463] = (N3)? mem[463] : 
                         (N0)? mem[981] : 1'b0;
  assign r_data_o[462] = (N3)? mem[462] : 
                         (N0)? mem[980] : 1'b0;
  assign r_data_o[461] = (N3)? mem[461] : 
                         (N0)? mem[979] : 1'b0;
  assign r_data_o[460] = (N3)? mem[460] : 
                         (N0)? mem[978] : 1'b0;
  assign r_data_o[459] = (N3)? mem[459] : 
                         (N0)? mem[977] : 1'b0;
  assign r_data_o[458] = (N3)? mem[458] : 
                         (N0)? mem[976] : 1'b0;
  assign r_data_o[457] = (N3)? mem[457] : 
                         (N0)? mem[975] : 1'b0;
  assign r_data_o[456] = (N3)? mem[456] : 
                         (N0)? mem[974] : 1'b0;
  assign r_data_o[455] = (N3)? mem[455] : 
                         (N0)? mem[973] : 1'b0;
  assign r_data_o[454] = (N3)? mem[454] : 
                         (N0)? mem[972] : 1'b0;
  assign r_data_o[453] = (N3)? mem[453] : 
                         (N0)? mem[971] : 1'b0;
  assign r_data_o[452] = (N3)? mem[452] : 
                         (N0)? mem[970] : 1'b0;
  assign r_data_o[451] = (N3)? mem[451] : 
                         (N0)? mem[969] : 1'b0;
  assign r_data_o[450] = (N3)? mem[450] : 
                         (N0)? mem[968] : 1'b0;
  assign r_data_o[449] = (N3)? mem[449] : 
                         (N0)? mem[967] : 1'b0;
  assign r_data_o[448] = (N3)? mem[448] : 
                         (N0)? mem[966] : 1'b0;
  assign r_data_o[447] = (N3)? mem[447] : 
                         (N0)? mem[965] : 1'b0;
  assign r_data_o[446] = (N3)? mem[446] : 
                         (N0)? mem[964] : 1'b0;
  assign r_data_o[445] = (N3)? mem[445] : 
                         (N0)? mem[963] : 1'b0;
  assign r_data_o[444] = (N3)? mem[444] : 
                         (N0)? mem[962] : 1'b0;
  assign r_data_o[443] = (N3)? mem[443] : 
                         (N0)? mem[961] : 1'b0;
  assign r_data_o[442] = (N3)? mem[442] : 
                         (N0)? mem[960] : 1'b0;
  assign r_data_o[441] = (N3)? mem[441] : 
                         (N0)? mem[959] : 1'b0;
  assign r_data_o[440] = (N3)? mem[440] : 
                         (N0)? mem[958] : 1'b0;
  assign r_data_o[439] = (N3)? mem[439] : 
                         (N0)? mem[957] : 1'b0;
  assign r_data_o[438] = (N3)? mem[438] : 
                         (N0)? mem[956] : 1'b0;
  assign r_data_o[437] = (N3)? mem[437] : 
                         (N0)? mem[955] : 1'b0;
  assign r_data_o[436] = (N3)? mem[436] : 
                         (N0)? mem[954] : 1'b0;
  assign r_data_o[435] = (N3)? mem[435] : 
                         (N0)? mem[953] : 1'b0;
  assign r_data_o[434] = (N3)? mem[434] : 
                         (N0)? mem[952] : 1'b0;
  assign r_data_o[433] = (N3)? mem[433] : 
                         (N0)? mem[951] : 1'b0;
  assign r_data_o[432] = (N3)? mem[432] : 
                         (N0)? mem[950] : 1'b0;
  assign r_data_o[431] = (N3)? mem[431] : 
                         (N0)? mem[949] : 1'b0;
  assign r_data_o[430] = (N3)? mem[430] : 
                         (N0)? mem[948] : 1'b0;
  assign r_data_o[429] = (N3)? mem[429] : 
                         (N0)? mem[947] : 1'b0;
  assign r_data_o[428] = (N3)? mem[428] : 
                         (N0)? mem[946] : 1'b0;
  assign r_data_o[427] = (N3)? mem[427] : 
                         (N0)? mem[945] : 1'b0;
  assign r_data_o[426] = (N3)? mem[426] : 
                         (N0)? mem[944] : 1'b0;
  assign r_data_o[425] = (N3)? mem[425] : 
                         (N0)? mem[943] : 1'b0;
  assign r_data_o[424] = (N3)? mem[424] : 
                         (N0)? mem[942] : 1'b0;
  assign r_data_o[423] = (N3)? mem[423] : 
                         (N0)? mem[941] : 1'b0;
  assign r_data_o[422] = (N3)? mem[422] : 
                         (N0)? mem[940] : 1'b0;
  assign r_data_o[421] = (N3)? mem[421] : 
                         (N0)? mem[939] : 1'b0;
  assign r_data_o[420] = (N3)? mem[420] : 
                         (N0)? mem[938] : 1'b0;
  assign r_data_o[419] = (N3)? mem[419] : 
                         (N0)? mem[937] : 1'b0;
  assign r_data_o[418] = (N3)? mem[418] : 
                         (N0)? mem[936] : 1'b0;
  assign r_data_o[417] = (N3)? mem[417] : 
                         (N0)? mem[935] : 1'b0;
  assign r_data_o[416] = (N3)? mem[416] : 
                         (N0)? mem[934] : 1'b0;
  assign r_data_o[415] = (N3)? mem[415] : 
                         (N0)? mem[933] : 1'b0;
  assign r_data_o[414] = (N3)? mem[414] : 
                         (N0)? mem[932] : 1'b0;
  assign r_data_o[413] = (N3)? mem[413] : 
                         (N0)? mem[931] : 1'b0;
  assign r_data_o[412] = (N3)? mem[412] : 
                         (N0)? mem[930] : 1'b0;
  assign r_data_o[411] = (N3)? mem[411] : 
                         (N0)? mem[929] : 1'b0;
  assign r_data_o[410] = (N3)? mem[410] : 
                         (N0)? mem[928] : 1'b0;
  assign r_data_o[409] = (N3)? mem[409] : 
                         (N0)? mem[927] : 1'b0;
  assign r_data_o[408] = (N3)? mem[408] : 
                         (N0)? mem[926] : 1'b0;
  assign r_data_o[407] = (N3)? mem[407] : 
                         (N0)? mem[925] : 1'b0;
  assign r_data_o[406] = (N3)? mem[406] : 
                         (N0)? mem[924] : 1'b0;
  assign r_data_o[405] = (N3)? mem[405] : 
                         (N0)? mem[923] : 1'b0;
  assign r_data_o[404] = (N3)? mem[404] : 
                         (N0)? mem[922] : 1'b0;
  assign r_data_o[403] = (N3)? mem[403] : 
                         (N0)? mem[921] : 1'b0;
  assign r_data_o[402] = (N3)? mem[402] : 
                         (N0)? mem[920] : 1'b0;
  assign r_data_o[401] = (N3)? mem[401] : 
                         (N0)? mem[919] : 1'b0;
  assign r_data_o[400] = (N3)? mem[400] : 
                         (N0)? mem[918] : 1'b0;
  assign r_data_o[399] = (N3)? mem[399] : 
                         (N0)? mem[917] : 1'b0;
  assign r_data_o[398] = (N3)? mem[398] : 
                         (N0)? mem[916] : 1'b0;
  assign r_data_o[397] = (N3)? mem[397] : 
                         (N0)? mem[915] : 1'b0;
  assign r_data_o[396] = (N3)? mem[396] : 
                         (N0)? mem[914] : 1'b0;
  assign r_data_o[395] = (N3)? mem[395] : 
                         (N0)? mem[913] : 1'b0;
  assign r_data_o[394] = (N3)? mem[394] : 
                         (N0)? mem[912] : 1'b0;
  assign r_data_o[393] = (N3)? mem[393] : 
                         (N0)? mem[911] : 1'b0;
  assign r_data_o[392] = (N3)? mem[392] : 
                         (N0)? mem[910] : 1'b0;
  assign r_data_o[391] = (N3)? mem[391] : 
                         (N0)? mem[909] : 1'b0;
  assign r_data_o[390] = (N3)? mem[390] : 
                         (N0)? mem[908] : 1'b0;
  assign r_data_o[389] = (N3)? mem[389] : 
                         (N0)? mem[907] : 1'b0;
  assign r_data_o[388] = (N3)? mem[388] : 
                         (N0)? mem[906] : 1'b0;
  assign r_data_o[387] = (N3)? mem[387] : 
                         (N0)? mem[905] : 1'b0;
  assign r_data_o[386] = (N3)? mem[386] : 
                         (N0)? mem[904] : 1'b0;
  assign r_data_o[385] = (N3)? mem[385] : 
                         (N0)? mem[903] : 1'b0;
  assign r_data_o[384] = (N3)? mem[384] : 
                         (N0)? mem[902] : 1'b0;
  assign r_data_o[383] = (N3)? mem[383] : 
                         (N0)? mem[901] : 1'b0;
  assign r_data_o[382] = (N3)? mem[382] : 
                         (N0)? mem[900] : 1'b0;
  assign r_data_o[381] = (N3)? mem[381] : 
                         (N0)? mem[899] : 1'b0;
  assign r_data_o[380] = (N3)? mem[380] : 
                         (N0)? mem[898] : 1'b0;
  assign r_data_o[379] = (N3)? mem[379] : 
                         (N0)? mem[897] : 1'b0;
  assign r_data_o[378] = (N3)? mem[378] : 
                         (N0)? mem[896] : 1'b0;
  assign r_data_o[377] = (N3)? mem[377] : 
                         (N0)? mem[895] : 1'b0;
  assign r_data_o[376] = (N3)? mem[376] : 
                         (N0)? mem[894] : 1'b0;
  assign r_data_o[375] = (N3)? mem[375] : 
                         (N0)? mem[893] : 1'b0;
  assign r_data_o[374] = (N3)? mem[374] : 
                         (N0)? mem[892] : 1'b0;
  assign r_data_o[373] = (N3)? mem[373] : 
                         (N0)? mem[891] : 1'b0;
  assign r_data_o[372] = (N3)? mem[372] : 
                         (N0)? mem[890] : 1'b0;
  assign r_data_o[371] = (N3)? mem[371] : 
                         (N0)? mem[889] : 1'b0;
  assign r_data_o[370] = (N3)? mem[370] : 
                         (N0)? mem[888] : 1'b0;
  assign r_data_o[369] = (N3)? mem[369] : 
                         (N0)? mem[887] : 1'b0;
  assign r_data_o[368] = (N3)? mem[368] : 
                         (N0)? mem[886] : 1'b0;
  assign r_data_o[367] = (N3)? mem[367] : 
                         (N0)? mem[885] : 1'b0;
  assign r_data_o[366] = (N3)? mem[366] : 
                         (N0)? mem[884] : 1'b0;
  assign r_data_o[365] = (N3)? mem[365] : 
                         (N0)? mem[883] : 1'b0;
  assign r_data_o[364] = (N3)? mem[364] : 
                         (N0)? mem[882] : 1'b0;
  assign r_data_o[363] = (N3)? mem[363] : 
                         (N0)? mem[881] : 1'b0;
  assign r_data_o[362] = (N3)? mem[362] : 
                         (N0)? mem[880] : 1'b0;
  assign r_data_o[361] = (N3)? mem[361] : 
                         (N0)? mem[879] : 1'b0;
  assign r_data_o[360] = (N3)? mem[360] : 
                         (N0)? mem[878] : 1'b0;
  assign r_data_o[359] = (N3)? mem[359] : 
                         (N0)? mem[877] : 1'b0;
  assign r_data_o[358] = (N3)? mem[358] : 
                         (N0)? mem[876] : 1'b0;
  assign r_data_o[357] = (N3)? mem[357] : 
                         (N0)? mem[875] : 1'b0;
  assign r_data_o[356] = (N3)? mem[356] : 
                         (N0)? mem[874] : 1'b0;
  assign r_data_o[355] = (N3)? mem[355] : 
                         (N0)? mem[873] : 1'b0;
  assign r_data_o[354] = (N3)? mem[354] : 
                         (N0)? mem[872] : 1'b0;
  assign r_data_o[353] = (N3)? mem[353] : 
                         (N0)? mem[871] : 1'b0;
  assign r_data_o[352] = (N3)? mem[352] : 
                         (N0)? mem[870] : 1'b0;
  assign r_data_o[351] = (N3)? mem[351] : 
                         (N0)? mem[869] : 1'b0;
  assign r_data_o[350] = (N3)? mem[350] : 
                         (N0)? mem[868] : 1'b0;
  assign r_data_o[349] = (N3)? mem[349] : 
                         (N0)? mem[867] : 1'b0;
  assign r_data_o[348] = (N3)? mem[348] : 
                         (N0)? mem[866] : 1'b0;
  assign r_data_o[347] = (N3)? mem[347] : 
                         (N0)? mem[865] : 1'b0;
  assign r_data_o[346] = (N3)? mem[346] : 
                         (N0)? mem[864] : 1'b0;
  assign r_data_o[345] = (N3)? mem[345] : 
                         (N0)? mem[863] : 1'b0;
  assign r_data_o[344] = (N3)? mem[344] : 
                         (N0)? mem[862] : 1'b0;
  assign r_data_o[343] = (N3)? mem[343] : 
                         (N0)? mem[861] : 1'b0;
  assign r_data_o[342] = (N3)? mem[342] : 
                         (N0)? mem[860] : 1'b0;
  assign r_data_o[341] = (N3)? mem[341] : 
                         (N0)? mem[859] : 1'b0;
  assign r_data_o[340] = (N3)? mem[340] : 
                         (N0)? mem[858] : 1'b0;
  assign r_data_o[339] = (N3)? mem[339] : 
                         (N0)? mem[857] : 1'b0;
  assign r_data_o[338] = (N3)? mem[338] : 
                         (N0)? mem[856] : 1'b0;
  assign r_data_o[337] = (N3)? mem[337] : 
                         (N0)? mem[855] : 1'b0;
  assign r_data_o[336] = (N3)? mem[336] : 
                         (N0)? mem[854] : 1'b0;
  assign r_data_o[335] = (N3)? mem[335] : 
                         (N0)? mem[853] : 1'b0;
  assign r_data_o[334] = (N3)? mem[334] : 
                         (N0)? mem[852] : 1'b0;
  assign r_data_o[333] = (N3)? mem[333] : 
                         (N0)? mem[851] : 1'b0;
  assign r_data_o[332] = (N3)? mem[332] : 
                         (N0)? mem[850] : 1'b0;
  assign r_data_o[331] = (N3)? mem[331] : 
                         (N0)? mem[849] : 1'b0;
  assign r_data_o[330] = (N3)? mem[330] : 
                         (N0)? mem[848] : 1'b0;
  assign r_data_o[329] = (N3)? mem[329] : 
                         (N0)? mem[847] : 1'b0;
  assign r_data_o[328] = (N3)? mem[328] : 
                         (N0)? mem[846] : 1'b0;
  assign r_data_o[327] = (N3)? mem[327] : 
                         (N0)? mem[845] : 1'b0;
  assign r_data_o[326] = (N3)? mem[326] : 
                         (N0)? mem[844] : 1'b0;
  assign r_data_o[325] = (N3)? mem[325] : 
                         (N0)? mem[843] : 1'b0;
  assign r_data_o[324] = (N3)? mem[324] : 
                         (N0)? mem[842] : 1'b0;
  assign r_data_o[323] = (N3)? mem[323] : 
                         (N0)? mem[841] : 1'b0;
  assign r_data_o[322] = (N3)? mem[322] : 
                         (N0)? mem[840] : 1'b0;
  assign r_data_o[321] = (N3)? mem[321] : 
                         (N0)? mem[839] : 1'b0;
  assign r_data_o[320] = (N3)? mem[320] : 
                         (N0)? mem[838] : 1'b0;
  assign r_data_o[319] = (N3)? mem[319] : 
                         (N0)? mem[837] : 1'b0;
  assign r_data_o[318] = (N3)? mem[318] : 
                         (N0)? mem[836] : 1'b0;
  assign r_data_o[317] = (N3)? mem[317] : 
                         (N0)? mem[835] : 1'b0;
  assign r_data_o[316] = (N3)? mem[316] : 
                         (N0)? mem[834] : 1'b0;
  assign r_data_o[315] = (N3)? mem[315] : 
                         (N0)? mem[833] : 1'b0;
  assign r_data_o[314] = (N3)? mem[314] : 
                         (N0)? mem[832] : 1'b0;
  assign r_data_o[313] = (N3)? mem[313] : 
                         (N0)? mem[831] : 1'b0;
  assign r_data_o[312] = (N3)? mem[312] : 
                         (N0)? mem[830] : 1'b0;
  assign r_data_o[311] = (N3)? mem[311] : 
                         (N0)? mem[829] : 1'b0;
  assign r_data_o[310] = (N3)? mem[310] : 
                         (N0)? mem[828] : 1'b0;
  assign r_data_o[309] = (N3)? mem[309] : 
                         (N0)? mem[827] : 1'b0;
  assign r_data_o[308] = (N3)? mem[308] : 
                         (N0)? mem[826] : 1'b0;
  assign r_data_o[307] = (N3)? mem[307] : 
                         (N0)? mem[825] : 1'b0;
  assign r_data_o[306] = (N3)? mem[306] : 
                         (N0)? mem[824] : 1'b0;
  assign r_data_o[305] = (N3)? mem[305] : 
                         (N0)? mem[823] : 1'b0;
  assign r_data_o[304] = (N3)? mem[304] : 
                         (N0)? mem[822] : 1'b0;
  assign r_data_o[303] = (N3)? mem[303] : 
                         (N0)? mem[821] : 1'b0;
  assign r_data_o[302] = (N3)? mem[302] : 
                         (N0)? mem[820] : 1'b0;
  assign r_data_o[301] = (N3)? mem[301] : 
                         (N0)? mem[819] : 1'b0;
  assign r_data_o[300] = (N3)? mem[300] : 
                         (N0)? mem[818] : 1'b0;
  assign r_data_o[299] = (N3)? mem[299] : 
                         (N0)? mem[817] : 1'b0;
  assign r_data_o[298] = (N3)? mem[298] : 
                         (N0)? mem[816] : 1'b0;
  assign r_data_o[297] = (N3)? mem[297] : 
                         (N0)? mem[815] : 1'b0;
  assign r_data_o[296] = (N3)? mem[296] : 
                         (N0)? mem[814] : 1'b0;
  assign r_data_o[295] = (N3)? mem[295] : 
                         (N0)? mem[813] : 1'b0;
  assign r_data_o[294] = (N3)? mem[294] : 
                         (N0)? mem[812] : 1'b0;
  assign r_data_o[293] = (N3)? mem[293] : 
                         (N0)? mem[811] : 1'b0;
  assign r_data_o[292] = (N3)? mem[292] : 
                         (N0)? mem[810] : 1'b0;
  assign r_data_o[291] = (N3)? mem[291] : 
                         (N0)? mem[809] : 1'b0;
  assign r_data_o[290] = (N3)? mem[290] : 
                         (N0)? mem[808] : 1'b0;
  assign r_data_o[289] = (N3)? mem[289] : 
                         (N0)? mem[807] : 1'b0;
  assign r_data_o[288] = (N3)? mem[288] : 
                         (N0)? mem[806] : 1'b0;
  assign r_data_o[287] = (N3)? mem[287] : 
                         (N0)? mem[805] : 1'b0;
  assign r_data_o[286] = (N3)? mem[286] : 
                         (N0)? mem[804] : 1'b0;
  assign r_data_o[285] = (N3)? mem[285] : 
                         (N0)? mem[803] : 1'b0;
  assign r_data_o[284] = (N3)? mem[284] : 
                         (N0)? mem[802] : 1'b0;
  assign r_data_o[283] = (N3)? mem[283] : 
                         (N0)? mem[801] : 1'b0;
  assign r_data_o[282] = (N3)? mem[282] : 
                         (N0)? mem[800] : 1'b0;
  assign r_data_o[281] = (N3)? mem[281] : 
                         (N0)? mem[799] : 1'b0;
  assign r_data_o[280] = (N3)? mem[280] : 
                         (N0)? mem[798] : 1'b0;
  assign r_data_o[279] = (N3)? mem[279] : 
                         (N0)? mem[797] : 1'b0;
  assign r_data_o[278] = (N3)? mem[278] : 
                         (N0)? mem[796] : 1'b0;
  assign r_data_o[277] = (N3)? mem[277] : 
                         (N0)? mem[795] : 1'b0;
  assign r_data_o[276] = (N3)? mem[276] : 
                         (N0)? mem[794] : 1'b0;
  assign r_data_o[275] = (N3)? mem[275] : 
                         (N0)? mem[793] : 1'b0;
  assign r_data_o[274] = (N3)? mem[274] : 
                         (N0)? mem[792] : 1'b0;
  assign r_data_o[273] = (N3)? mem[273] : 
                         (N0)? mem[791] : 1'b0;
  assign r_data_o[272] = (N3)? mem[272] : 
                         (N0)? mem[790] : 1'b0;
  assign r_data_o[271] = (N3)? mem[271] : 
                         (N0)? mem[789] : 1'b0;
  assign r_data_o[270] = (N3)? mem[270] : 
                         (N0)? mem[788] : 1'b0;
  assign r_data_o[269] = (N3)? mem[269] : 
                         (N0)? mem[787] : 1'b0;
  assign r_data_o[268] = (N3)? mem[268] : 
                         (N0)? mem[786] : 1'b0;
  assign r_data_o[267] = (N3)? mem[267] : 
                         (N0)? mem[785] : 1'b0;
  assign r_data_o[266] = (N3)? mem[266] : 
                         (N0)? mem[784] : 1'b0;
  assign r_data_o[265] = (N3)? mem[265] : 
                         (N0)? mem[783] : 1'b0;
  assign r_data_o[264] = (N3)? mem[264] : 
                         (N0)? mem[782] : 1'b0;
  assign r_data_o[263] = (N3)? mem[263] : 
                         (N0)? mem[781] : 1'b0;
  assign r_data_o[262] = (N3)? mem[262] : 
                         (N0)? mem[780] : 1'b0;
  assign r_data_o[261] = (N3)? mem[261] : 
                         (N0)? mem[779] : 1'b0;
  assign r_data_o[260] = (N3)? mem[260] : 
                         (N0)? mem[778] : 1'b0;
  assign r_data_o[259] = (N3)? mem[259] : 
                         (N0)? mem[777] : 1'b0;
  assign r_data_o[258] = (N3)? mem[258] : 
                         (N0)? mem[776] : 1'b0;
  assign r_data_o[257] = (N3)? mem[257] : 
                         (N0)? mem[775] : 1'b0;
  assign r_data_o[256] = (N3)? mem[256] : 
                         (N0)? mem[774] : 1'b0;
  assign r_data_o[255] = (N3)? mem[255] : 
                         (N0)? mem[773] : 1'b0;
  assign r_data_o[254] = (N3)? mem[254] : 
                         (N0)? mem[772] : 1'b0;
  assign r_data_o[253] = (N3)? mem[253] : 
                         (N0)? mem[771] : 1'b0;
  assign r_data_o[252] = (N3)? mem[252] : 
                         (N0)? mem[770] : 1'b0;
  assign r_data_o[251] = (N3)? mem[251] : 
                         (N0)? mem[769] : 1'b0;
  assign r_data_o[250] = (N3)? mem[250] : 
                         (N0)? mem[768] : 1'b0;
  assign r_data_o[249] = (N3)? mem[249] : 
                         (N0)? mem[767] : 1'b0;
  assign r_data_o[248] = (N3)? mem[248] : 
                         (N0)? mem[766] : 1'b0;
  assign r_data_o[247] = (N3)? mem[247] : 
                         (N0)? mem[765] : 1'b0;
  assign r_data_o[246] = (N3)? mem[246] : 
                         (N0)? mem[764] : 1'b0;
  assign r_data_o[245] = (N3)? mem[245] : 
                         (N0)? mem[763] : 1'b0;
  assign r_data_o[244] = (N3)? mem[244] : 
                         (N0)? mem[762] : 1'b0;
  assign r_data_o[243] = (N3)? mem[243] : 
                         (N0)? mem[761] : 1'b0;
  assign r_data_o[242] = (N3)? mem[242] : 
                         (N0)? mem[760] : 1'b0;
  assign r_data_o[241] = (N3)? mem[241] : 
                         (N0)? mem[759] : 1'b0;
  assign r_data_o[240] = (N3)? mem[240] : 
                         (N0)? mem[758] : 1'b0;
  assign r_data_o[239] = (N3)? mem[239] : 
                         (N0)? mem[757] : 1'b0;
  assign r_data_o[238] = (N3)? mem[238] : 
                         (N0)? mem[756] : 1'b0;
  assign r_data_o[237] = (N3)? mem[237] : 
                         (N0)? mem[755] : 1'b0;
  assign r_data_o[236] = (N3)? mem[236] : 
                         (N0)? mem[754] : 1'b0;
  assign r_data_o[235] = (N3)? mem[235] : 
                         (N0)? mem[753] : 1'b0;
  assign r_data_o[234] = (N3)? mem[234] : 
                         (N0)? mem[752] : 1'b0;
  assign r_data_o[233] = (N3)? mem[233] : 
                         (N0)? mem[751] : 1'b0;
  assign r_data_o[232] = (N3)? mem[232] : 
                         (N0)? mem[750] : 1'b0;
  assign r_data_o[231] = (N3)? mem[231] : 
                         (N0)? mem[749] : 1'b0;
  assign r_data_o[230] = (N3)? mem[230] : 
                         (N0)? mem[748] : 1'b0;
  assign r_data_o[229] = (N3)? mem[229] : 
                         (N0)? mem[747] : 1'b0;
  assign r_data_o[228] = (N3)? mem[228] : 
                         (N0)? mem[746] : 1'b0;
  assign r_data_o[227] = (N3)? mem[227] : 
                         (N0)? mem[745] : 1'b0;
  assign r_data_o[226] = (N3)? mem[226] : 
                         (N0)? mem[744] : 1'b0;
  assign r_data_o[225] = (N3)? mem[225] : 
                         (N0)? mem[743] : 1'b0;
  assign r_data_o[224] = (N3)? mem[224] : 
                         (N0)? mem[742] : 1'b0;
  assign r_data_o[223] = (N3)? mem[223] : 
                         (N0)? mem[741] : 1'b0;
  assign r_data_o[222] = (N3)? mem[222] : 
                         (N0)? mem[740] : 1'b0;
  assign r_data_o[221] = (N3)? mem[221] : 
                         (N0)? mem[739] : 1'b0;
  assign r_data_o[220] = (N3)? mem[220] : 
                         (N0)? mem[738] : 1'b0;
  assign r_data_o[219] = (N3)? mem[219] : 
                         (N0)? mem[737] : 1'b0;
  assign r_data_o[218] = (N3)? mem[218] : 
                         (N0)? mem[736] : 1'b0;
  assign r_data_o[217] = (N3)? mem[217] : 
                         (N0)? mem[735] : 1'b0;
  assign r_data_o[216] = (N3)? mem[216] : 
                         (N0)? mem[734] : 1'b0;
  assign r_data_o[215] = (N3)? mem[215] : 
                         (N0)? mem[733] : 1'b0;
  assign r_data_o[214] = (N3)? mem[214] : 
                         (N0)? mem[732] : 1'b0;
  assign r_data_o[213] = (N3)? mem[213] : 
                         (N0)? mem[731] : 1'b0;
  assign r_data_o[212] = (N3)? mem[212] : 
                         (N0)? mem[730] : 1'b0;
  assign r_data_o[211] = (N3)? mem[211] : 
                         (N0)? mem[729] : 1'b0;
  assign r_data_o[210] = (N3)? mem[210] : 
                         (N0)? mem[728] : 1'b0;
  assign r_data_o[209] = (N3)? mem[209] : 
                         (N0)? mem[727] : 1'b0;
  assign r_data_o[208] = (N3)? mem[208] : 
                         (N0)? mem[726] : 1'b0;
  assign r_data_o[207] = (N3)? mem[207] : 
                         (N0)? mem[725] : 1'b0;
  assign r_data_o[206] = (N3)? mem[206] : 
                         (N0)? mem[724] : 1'b0;
  assign r_data_o[205] = (N3)? mem[205] : 
                         (N0)? mem[723] : 1'b0;
  assign r_data_o[204] = (N3)? mem[204] : 
                         (N0)? mem[722] : 1'b0;
  assign r_data_o[203] = (N3)? mem[203] : 
                         (N0)? mem[721] : 1'b0;
  assign r_data_o[202] = (N3)? mem[202] : 
                         (N0)? mem[720] : 1'b0;
  assign r_data_o[201] = (N3)? mem[201] : 
                         (N0)? mem[719] : 1'b0;
  assign r_data_o[200] = (N3)? mem[200] : 
                         (N0)? mem[718] : 1'b0;
  assign r_data_o[199] = (N3)? mem[199] : 
                         (N0)? mem[717] : 1'b0;
  assign r_data_o[198] = (N3)? mem[198] : 
                         (N0)? mem[716] : 1'b0;
  assign r_data_o[197] = (N3)? mem[197] : 
                         (N0)? mem[715] : 1'b0;
  assign r_data_o[196] = (N3)? mem[196] : 
                         (N0)? mem[714] : 1'b0;
  assign r_data_o[195] = (N3)? mem[195] : 
                         (N0)? mem[713] : 1'b0;
  assign r_data_o[194] = (N3)? mem[194] : 
                         (N0)? mem[712] : 1'b0;
  assign r_data_o[193] = (N3)? mem[193] : 
                         (N0)? mem[711] : 1'b0;
  assign r_data_o[192] = (N3)? mem[192] : 
                         (N0)? mem[710] : 1'b0;
  assign r_data_o[191] = (N3)? mem[191] : 
                         (N0)? mem[709] : 1'b0;
  assign r_data_o[190] = (N3)? mem[190] : 
                         (N0)? mem[708] : 1'b0;
  assign r_data_o[189] = (N3)? mem[189] : 
                         (N0)? mem[707] : 1'b0;
  assign r_data_o[188] = (N3)? mem[188] : 
                         (N0)? mem[706] : 1'b0;
  assign r_data_o[187] = (N3)? mem[187] : 
                         (N0)? mem[705] : 1'b0;
  assign r_data_o[186] = (N3)? mem[186] : 
                         (N0)? mem[704] : 1'b0;
  assign r_data_o[185] = (N3)? mem[185] : 
                         (N0)? mem[703] : 1'b0;
  assign r_data_o[184] = (N3)? mem[184] : 
                         (N0)? mem[702] : 1'b0;
  assign r_data_o[183] = (N3)? mem[183] : 
                         (N0)? mem[701] : 1'b0;
  assign r_data_o[182] = (N3)? mem[182] : 
                         (N0)? mem[700] : 1'b0;
  assign r_data_o[181] = (N3)? mem[181] : 
                         (N0)? mem[699] : 1'b0;
  assign r_data_o[180] = (N3)? mem[180] : 
                         (N0)? mem[698] : 1'b0;
  assign r_data_o[179] = (N3)? mem[179] : 
                         (N0)? mem[697] : 1'b0;
  assign r_data_o[178] = (N3)? mem[178] : 
                         (N0)? mem[696] : 1'b0;
  assign r_data_o[177] = (N3)? mem[177] : 
                         (N0)? mem[695] : 1'b0;
  assign r_data_o[176] = (N3)? mem[176] : 
                         (N0)? mem[694] : 1'b0;
  assign r_data_o[175] = (N3)? mem[175] : 
                         (N0)? mem[693] : 1'b0;
  assign r_data_o[174] = (N3)? mem[174] : 
                         (N0)? mem[692] : 1'b0;
  assign r_data_o[173] = (N3)? mem[173] : 
                         (N0)? mem[691] : 1'b0;
  assign r_data_o[172] = (N3)? mem[172] : 
                         (N0)? mem[690] : 1'b0;
  assign r_data_o[171] = (N3)? mem[171] : 
                         (N0)? mem[689] : 1'b0;
  assign r_data_o[170] = (N3)? mem[170] : 
                         (N0)? mem[688] : 1'b0;
  assign r_data_o[169] = (N3)? mem[169] : 
                         (N0)? mem[687] : 1'b0;
  assign r_data_o[168] = (N3)? mem[168] : 
                         (N0)? mem[686] : 1'b0;
  assign r_data_o[167] = (N3)? mem[167] : 
                         (N0)? mem[685] : 1'b0;
  assign r_data_o[166] = (N3)? mem[166] : 
                         (N0)? mem[684] : 1'b0;
  assign r_data_o[165] = (N3)? mem[165] : 
                         (N0)? mem[683] : 1'b0;
  assign r_data_o[164] = (N3)? mem[164] : 
                         (N0)? mem[682] : 1'b0;
  assign r_data_o[163] = (N3)? mem[163] : 
                         (N0)? mem[681] : 1'b0;
  assign r_data_o[162] = (N3)? mem[162] : 
                         (N0)? mem[680] : 1'b0;
  assign r_data_o[161] = (N3)? mem[161] : 
                         (N0)? mem[679] : 1'b0;
  assign r_data_o[160] = (N3)? mem[160] : 
                         (N0)? mem[678] : 1'b0;
  assign r_data_o[159] = (N3)? mem[159] : 
                         (N0)? mem[677] : 1'b0;
  assign r_data_o[158] = (N3)? mem[158] : 
                         (N0)? mem[676] : 1'b0;
  assign r_data_o[157] = (N3)? mem[157] : 
                         (N0)? mem[675] : 1'b0;
  assign r_data_o[156] = (N3)? mem[156] : 
                         (N0)? mem[674] : 1'b0;
  assign r_data_o[155] = (N3)? mem[155] : 
                         (N0)? mem[673] : 1'b0;
  assign r_data_o[154] = (N3)? mem[154] : 
                         (N0)? mem[672] : 1'b0;
  assign r_data_o[153] = (N3)? mem[153] : 
                         (N0)? mem[671] : 1'b0;
  assign r_data_o[152] = (N3)? mem[152] : 
                         (N0)? mem[670] : 1'b0;
  assign r_data_o[151] = (N3)? mem[151] : 
                         (N0)? mem[669] : 1'b0;
  assign r_data_o[150] = (N3)? mem[150] : 
                         (N0)? mem[668] : 1'b0;
  assign r_data_o[149] = (N3)? mem[149] : 
                         (N0)? mem[667] : 1'b0;
  assign r_data_o[148] = (N3)? mem[148] : 
                         (N0)? mem[666] : 1'b0;
  assign r_data_o[147] = (N3)? mem[147] : 
                         (N0)? mem[665] : 1'b0;
  assign r_data_o[146] = (N3)? mem[146] : 
                         (N0)? mem[664] : 1'b0;
  assign r_data_o[145] = (N3)? mem[145] : 
                         (N0)? mem[663] : 1'b0;
  assign r_data_o[144] = (N3)? mem[144] : 
                         (N0)? mem[662] : 1'b0;
  assign r_data_o[143] = (N3)? mem[143] : 
                         (N0)? mem[661] : 1'b0;
  assign r_data_o[142] = (N3)? mem[142] : 
                         (N0)? mem[660] : 1'b0;
  assign r_data_o[141] = (N3)? mem[141] : 
                         (N0)? mem[659] : 1'b0;
  assign r_data_o[140] = (N3)? mem[140] : 
                         (N0)? mem[658] : 1'b0;
  assign r_data_o[139] = (N3)? mem[139] : 
                         (N0)? mem[657] : 1'b0;
  assign r_data_o[138] = (N3)? mem[138] : 
                         (N0)? mem[656] : 1'b0;
  assign r_data_o[137] = (N3)? mem[137] : 
                         (N0)? mem[655] : 1'b0;
  assign r_data_o[136] = (N3)? mem[136] : 
                         (N0)? mem[654] : 1'b0;
  assign r_data_o[135] = (N3)? mem[135] : 
                         (N0)? mem[653] : 1'b0;
  assign r_data_o[134] = (N3)? mem[134] : 
                         (N0)? mem[652] : 1'b0;
  assign r_data_o[133] = (N3)? mem[133] : 
                         (N0)? mem[651] : 1'b0;
  assign r_data_o[132] = (N3)? mem[132] : 
                         (N0)? mem[650] : 1'b0;
  assign r_data_o[131] = (N3)? mem[131] : 
                         (N0)? mem[649] : 1'b0;
  assign r_data_o[130] = (N3)? mem[130] : 
                         (N0)? mem[648] : 1'b0;
  assign r_data_o[129] = (N3)? mem[129] : 
                         (N0)? mem[647] : 1'b0;
  assign r_data_o[128] = (N3)? mem[128] : 
                         (N0)? mem[646] : 1'b0;
  assign r_data_o[127] = (N3)? mem[127] : 
                         (N0)? mem[645] : 1'b0;
  assign r_data_o[126] = (N3)? mem[126] : 
                         (N0)? mem[644] : 1'b0;
  assign r_data_o[125] = (N3)? mem[125] : 
                         (N0)? mem[643] : 1'b0;
  assign r_data_o[124] = (N3)? mem[124] : 
                         (N0)? mem[642] : 1'b0;
  assign r_data_o[123] = (N3)? mem[123] : 
                         (N0)? mem[641] : 1'b0;
  assign r_data_o[122] = (N3)? mem[122] : 
                         (N0)? mem[640] : 1'b0;
  assign r_data_o[121] = (N3)? mem[121] : 
                         (N0)? mem[639] : 1'b0;
  assign r_data_o[120] = (N3)? mem[120] : 
                         (N0)? mem[638] : 1'b0;
  assign r_data_o[119] = (N3)? mem[119] : 
                         (N0)? mem[637] : 1'b0;
  assign r_data_o[118] = (N3)? mem[118] : 
                         (N0)? mem[636] : 1'b0;
  assign r_data_o[117] = (N3)? mem[117] : 
                         (N0)? mem[635] : 1'b0;
  assign r_data_o[116] = (N3)? mem[116] : 
                         (N0)? mem[634] : 1'b0;
  assign r_data_o[115] = (N3)? mem[115] : 
                         (N0)? mem[633] : 1'b0;
  assign r_data_o[114] = (N3)? mem[114] : 
                         (N0)? mem[632] : 1'b0;
  assign r_data_o[113] = (N3)? mem[113] : 
                         (N0)? mem[631] : 1'b0;
  assign r_data_o[112] = (N3)? mem[112] : 
                         (N0)? mem[630] : 1'b0;
  assign r_data_o[111] = (N3)? mem[111] : 
                         (N0)? mem[629] : 1'b0;
  assign r_data_o[110] = (N3)? mem[110] : 
                         (N0)? mem[628] : 1'b0;
  assign r_data_o[109] = (N3)? mem[109] : 
                         (N0)? mem[627] : 1'b0;
  assign r_data_o[108] = (N3)? mem[108] : 
                         (N0)? mem[626] : 1'b0;
  assign r_data_o[107] = (N3)? mem[107] : 
                         (N0)? mem[625] : 1'b0;
  assign r_data_o[106] = (N3)? mem[106] : 
                         (N0)? mem[624] : 1'b0;
  assign r_data_o[105] = (N3)? mem[105] : 
                         (N0)? mem[623] : 1'b0;
  assign r_data_o[104] = (N3)? mem[104] : 
                         (N0)? mem[622] : 1'b0;
  assign r_data_o[103] = (N3)? mem[103] : 
                         (N0)? mem[621] : 1'b0;
  assign r_data_o[102] = (N3)? mem[102] : 
                         (N0)? mem[620] : 1'b0;
  assign r_data_o[101] = (N3)? mem[101] : 
                         (N0)? mem[619] : 1'b0;
  assign r_data_o[100] = (N3)? mem[100] : 
                         (N0)? mem[618] : 1'b0;
  assign r_data_o[99] = (N3)? mem[99] : 
                        (N0)? mem[617] : 1'b0;
  assign r_data_o[98] = (N3)? mem[98] : 
                        (N0)? mem[616] : 1'b0;
  assign r_data_o[97] = (N3)? mem[97] : 
                        (N0)? mem[615] : 1'b0;
  assign r_data_o[96] = (N3)? mem[96] : 
                        (N0)? mem[614] : 1'b0;
  assign r_data_o[95] = (N3)? mem[95] : 
                        (N0)? mem[613] : 1'b0;
  assign r_data_o[94] = (N3)? mem[94] : 
                        (N0)? mem[612] : 1'b0;
  assign r_data_o[93] = (N3)? mem[93] : 
                        (N0)? mem[611] : 1'b0;
  assign r_data_o[92] = (N3)? mem[92] : 
                        (N0)? mem[610] : 1'b0;
  assign r_data_o[91] = (N3)? mem[91] : 
                        (N0)? mem[609] : 1'b0;
  assign r_data_o[90] = (N3)? mem[90] : 
                        (N0)? mem[608] : 1'b0;
  assign r_data_o[89] = (N3)? mem[89] : 
                        (N0)? mem[607] : 1'b0;
  assign r_data_o[88] = (N3)? mem[88] : 
                        (N0)? mem[606] : 1'b0;
  assign r_data_o[87] = (N3)? mem[87] : 
                        (N0)? mem[605] : 1'b0;
  assign r_data_o[86] = (N3)? mem[86] : 
                        (N0)? mem[604] : 1'b0;
  assign r_data_o[85] = (N3)? mem[85] : 
                        (N0)? mem[603] : 1'b0;
  assign r_data_o[84] = (N3)? mem[84] : 
                        (N0)? mem[602] : 1'b0;
  assign r_data_o[83] = (N3)? mem[83] : 
                        (N0)? mem[601] : 1'b0;
  assign r_data_o[82] = (N3)? mem[82] : 
                        (N0)? mem[600] : 1'b0;
  assign r_data_o[81] = (N3)? mem[81] : 
                        (N0)? mem[599] : 1'b0;
  assign r_data_o[80] = (N3)? mem[80] : 
                        (N0)? mem[598] : 1'b0;
  assign r_data_o[79] = (N3)? mem[79] : 
                        (N0)? mem[597] : 1'b0;
  assign r_data_o[78] = (N3)? mem[78] : 
                        (N0)? mem[596] : 1'b0;
  assign r_data_o[77] = (N3)? mem[77] : 
                        (N0)? mem[595] : 1'b0;
  assign r_data_o[76] = (N3)? mem[76] : 
                        (N0)? mem[594] : 1'b0;
  assign r_data_o[75] = (N3)? mem[75] : 
                        (N0)? mem[593] : 1'b0;
  assign r_data_o[74] = (N3)? mem[74] : 
                        (N0)? mem[592] : 1'b0;
  assign r_data_o[73] = (N3)? mem[73] : 
                        (N0)? mem[591] : 1'b0;
  assign r_data_o[72] = (N3)? mem[72] : 
                        (N0)? mem[590] : 1'b0;
  assign r_data_o[71] = (N3)? mem[71] : 
                        (N0)? mem[589] : 1'b0;
  assign r_data_o[70] = (N3)? mem[70] : 
                        (N0)? mem[588] : 1'b0;
  assign r_data_o[69] = (N3)? mem[69] : 
                        (N0)? mem[587] : 1'b0;
  assign r_data_o[68] = (N3)? mem[68] : 
                        (N0)? mem[586] : 1'b0;
  assign r_data_o[67] = (N3)? mem[67] : 
                        (N0)? mem[585] : 1'b0;
  assign r_data_o[66] = (N3)? mem[66] : 
                        (N0)? mem[584] : 1'b0;
  assign r_data_o[65] = (N3)? mem[65] : 
                        (N0)? mem[583] : 1'b0;
  assign r_data_o[64] = (N3)? mem[64] : 
                        (N0)? mem[582] : 1'b0;
  assign r_data_o[63] = (N3)? mem[63] : 
                        (N0)? mem[581] : 1'b0;
  assign r_data_o[62] = (N3)? mem[62] : 
                        (N0)? mem[580] : 1'b0;
  assign r_data_o[61] = (N3)? mem[61] : 
                        (N0)? mem[579] : 1'b0;
  assign r_data_o[60] = (N3)? mem[60] : 
                        (N0)? mem[578] : 1'b0;
  assign r_data_o[59] = (N3)? mem[59] : 
                        (N0)? mem[577] : 1'b0;
  assign r_data_o[58] = (N3)? mem[58] : 
                        (N0)? mem[576] : 1'b0;
  assign r_data_o[57] = (N3)? mem[57] : 
                        (N0)? mem[575] : 1'b0;
  assign r_data_o[56] = (N3)? mem[56] : 
                        (N0)? mem[574] : 1'b0;
  assign r_data_o[55] = (N3)? mem[55] : 
                        (N0)? mem[573] : 1'b0;
  assign r_data_o[54] = (N3)? mem[54] : 
                        (N0)? mem[572] : 1'b0;
  assign r_data_o[53] = (N3)? mem[53] : 
                        (N0)? mem[571] : 1'b0;
  assign r_data_o[52] = (N3)? mem[52] : 
                        (N0)? mem[570] : 1'b0;
  assign r_data_o[51] = (N3)? mem[51] : 
                        (N0)? mem[569] : 1'b0;
  assign r_data_o[50] = (N3)? mem[50] : 
                        (N0)? mem[568] : 1'b0;
  assign r_data_o[49] = (N3)? mem[49] : 
                        (N0)? mem[567] : 1'b0;
  assign r_data_o[48] = (N3)? mem[48] : 
                        (N0)? mem[566] : 1'b0;
  assign r_data_o[47] = (N3)? mem[47] : 
                        (N0)? mem[565] : 1'b0;
  assign r_data_o[46] = (N3)? mem[46] : 
                        (N0)? mem[564] : 1'b0;
  assign r_data_o[45] = (N3)? mem[45] : 
                        (N0)? mem[563] : 1'b0;
  assign r_data_o[44] = (N3)? mem[44] : 
                        (N0)? mem[562] : 1'b0;
  assign r_data_o[43] = (N3)? mem[43] : 
                        (N0)? mem[561] : 1'b0;
  assign r_data_o[42] = (N3)? mem[42] : 
                        (N0)? mem[560] : 1'b0;
  assign r_data_o[41] = (N3)? mem[41] : 
                        (N0)? mem[559] : 1'b0;
  assign r_data_o[40] = (N3)? mem[40] : 
                        (N0)? mem[558] : 1'b0;
  assign r_data_o[39] = (N3)? mem[39] : 
                        (N0)? mem[557] : 1'b0;
  assign r_data_o[38] = (N3)? mem[38] : 
                        (N0)? mem[556] : 1'b0;
  assign r_data_o[37] = (N3)? mem[37] : 
                        (N0)? mem[555] : 1'b0;
  assign r_data_o[36] = (N3)? mem[36] : 
                        (N0)? mem[554] : 1'b0;
  assign r_data_o[35] = (N3)? mem[35] : 
                        (N0)? mem[553] : 1'b0;
  assign r_data_o[34] = (N3)? mem[34] : 
                        (N0)? mem[552] : 1'b0;
  assign r_data_o[33] = (N3)? mem[33] : 
                        (N0)? mem[551] : 1'b0;
  assign r_data_o[32] = (N3)? mem[32] : 
                        (N0)? mem[550] : 1'b0;
  assign r_data_o[31] = (N3)? mem[31] : 
                        (N0)? mem[549] : 1'b0;
  assign r_data_o[30] = (N3)? mem[30] : 
                        (N0)? mem[548] : 1'b0;
  assign r_data_o[29] = (N3)? mem[29] : 
                        (N0)? mem[547] : 1'b0;
  assign r_data_o[28] = (N3)? mem[28] : 
                        (N0)? mem[546] : 1'b0;
  assign r_data_o[27] = (N3)? mem[27] : 
                        (N0)? mem[545] : 1'b0;
  assign r_data_o[26] = (N3)? mem[26] : 
                        (N0)? mem[544] : 1'b0;
  assign r_data_o[25] = (N3)? mem[25] : 
                        (N0)? mem[543] : 1'b0;
  assign r_data_o[24] = (N3)? mem[24] : 
                        (N0)? mem[542] : 1'b0;
  assign r_data_o[23] = (N3)? mem[23] : 
                        (N0)? mem[541] : 1'b0;
  assign r_data_o[22] = (N3)? mem[22] : 
                        (N0)? mem[540] : 1'b0;
  assign r_data_o[21] = (N3)? mem[21] : 
                        (N0)? mem[539] : 1'b0;
  assign r_data_o[20] = (N3)? mem[20] : 
                        (N0)? mem[538] : 1'b0;
  assign r_data_o[19] = (N3)? mem[19] : 
                        (N0)? mem[537] : 1'b0;
  assign r_data_o[18] = (N3)? mem[18] : 
                        (N0)? mem[536] : 1'b0;
  assign r_data_o[17] = (N3)? mem[17] : 
                        (N0)? mem[535] : 1'b0;
  assign r_data_o[16] = (N3)? mem[16] : 
                        (N0)? mem[534] : 1'b0;
  assign r_data_o[15] = (N3)? mem[15] : 
                        (N0)? mem[533] : 1'b0;
  assign r_data_o[14] = (N3)? mem[14] : 
                        (N0)? mem[532] : 1'b0;
  assign r_data_o[13] = (N3)? mem[13] : 
                        (N0)? mem[531] : 1'b0;
  assign r_data_o[12] = (N3)? mem[12] : 
                        (N0)? mem[530] : 1'b0;
  assign r_data_o[11] = (N3)? mem[11] : 
                        (N0)? mem[529] : 1'b0;
  assign r_data_o[10] = (N3)? mem[10] : 
                        (N0)? mem[528] : 1'b0;
  assign r_data_o[9] = (N3)? mem[9] : 
                       (N0)? mem[527] : 1'b0;
  assign r_data_o[8] = (N3)? mem[8] : 
                       (N0)? mem[526] : 1'b0;
  assign r_data_o[7] = (N3)? mem[7] : 
                       (N0)? mem[525] : 1'b0;
  assign r_data_o[6] = (N3)? mem[6] : 
                       (N0)? mem[524] : 1'b0;
  assign r_data_o[5] = (N3)? mem[5] : 
                       (N0)? mem[523] : 1'b0;
  assign r_data_o[4] = (N3)? mem[4] : 
                       (N0)? mem[522] : 1'b0;
  assign r_data_o[3] = (N3)? mem[3] : 
                       (N0)? mem[521] : 1'b0;
  assign r_data_o[2] = (N3)? mem[2] : 
                       (N0)? mem[520] : 1'b0;
  assign r_data_o[1] = (N3)? mem[1] : 
                       (N0)? mem[519] : 1'b0;
  assign r_data_o[0] = (N3)? mem[0] : 
                       (N0)? mem[518] : 1'b0;
  assign N5 = ~w_addr_i[0];
  assign { N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7 } = (N1)? { w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], N5, N5, N5, N5, N5, N5 } : 
                                                                       (N2)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N1 = w_v_i;
  assign N2 = N4;
  assign N3 = ~r_addr_i[0];
  assign N4 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N13) begin
      { mem[1035:937], mem[518:518] } <= { w_data_i[517:419], w_data_i[0:0] };
    end 
    if(N14) begin
      { mem[936:838], mem[519:519] } <= { w_data_i[418:320], w_data_i[1:1] };
    end 
    if(N15) begin
      { mem[837:739], mem[520:520] } <= { w_data_i[319:221], w_data_i[2:2] };
    end 
    if(N16) begin
      { mem[738:640], mem[521:521] } <= { w_data_i[220:122], w_data_i[3:3] };
    end 
    if(N17) begin
      { mem[639:541], mem[522:522] } <= { w_data_i[121:23], w_data_i[4:4] };
    end 
    if(N18) begin
      { mem[540:523] } <= { w_data_i[22:5] };
    end 
    if(N7) begin
      { mem[517:419], mem[0:0] } <= { w_data_i[517:419], w_data_i[0:0] };
    end 
    if(N8) begin
      { mem[418:320], mem[1:1] } <= { w_data_i[418:320], w_data_i[1:1] };
    end 
    if(N9) begin
      { mem[319:221], mem[2:2] } <= { w_data_i[319:221], w_data_i[2:2] };
    end 
    if(N10) begin
      { mem[220:122], mem[3:3] } <= { w_data_i[220:122], w_data_i[3:3] };
    end 
    if(N11) begin
      { mem[121:23], mem[4:4] } <= { w_data_i[121:23], w_data_i[4:4] };
    end 
    if(N12) begin
      { mem[22:5] } <= { w_data_i[22:5] };
    end 
  end


endmodule



module bsg_mem_1r1w_width_p518_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [517:0] w_data_i;
  input [0:0] r_addr_i;
  output [517:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [517:0] r_data_o;

  bsg_mem_1r1w_synth_width_p518_els_p2_read_write_same_addr_p0_harden_p0
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i[0]),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i[0]),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_two_fifo_width_p518
(
  clk_i,
  reset_i,
  ready_o,
  data_i,
  v_i,
  v_o,
  data_o,
  yumi_i
);

  input [517:0] data_i;
  output [517:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [517:0] data_o;
  wire ready_o,v_o,N0,N1,enq_i,n_0_net_,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,
  N15,N16,N17,N18,N19,N20,N21,N22,N23,N24;
  reg full_r,tail_r,head_r,empty_r;

  bsg_mem_1r1w_width_p518_els_p2_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enq_i),
    .w_addr_i(tail_r),
    .w_data_i(data_i),
    .r_v_i(n_0_net_),
    .r_addr_i(head_r),
    .r_data_o(data_o)
  );

  assign N9 = (N0)? 1'b1 : 
              (N1)? N5 : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign N10 = (N0)? 1'b0 : 
               (N1)? N4 : 1'b0;
  assign N11 = (N0)? 1'b1 : 
               (N1)? yumi_i : 1'b0;
  assign N12 = (N0)? 1'b0 : 
               (N1)? N6 : 1'b0;
  assign N13 = (N0)? 1'b1 : 
               (N1)? N7 : 1'b0;
  assign N14 = (N0)? 1'b0 : 
               (N1)? N8 : 1'b0;
  assign n_0_net_ = ~empty_r;
  assign v_o = ~empty_r;
  assign ready_o = ~full_r;
  assign enq_i = v_i & N15;
  assign N15 = ~full_r;
  assign N2 = ~reset_i;
  assign N3 = reset_i;
  assign N5 = enq_i;
  assign N4 = ~tail_r;
  assign N6 = ~head_r;
  assign N7 = N17 | N19;
  assign N17 = empty_r & N16;
  assign N16 = ~enq_i;
  assign N19 = N18 & N16;
  assign N18 = N15 & yumi_i;
  assign N8 = N23 | N24;
  assign N23 = N21 & N22;
  assign N21 = N20 & enq_i;
  assign N20 = ~empty_r;
  assign N22 = ~yumi_i;
  assign N24 = full_r & N22;

  always @(posedge clk_i) begin
    if(1'b1) begin
      full_r <= N14;
      empty_r <= N13;
    end 
    if(N9) begin
      tail_r <= N10;
    end 
    if(N11) begin
      head_r <= N12;
    end 
  end


endmodule



module bp_fe_lce_data_cmd_02
(
  clk_i,
  reset_i,
  cce_data_received_o,
  tr_data_received_o,
  uncached_data_received_o,
  miss_addr_i,
  lce_data_cmd_i,
  lce_data_cmd_v_i,
  lce_data_cmd_ready_o,
  data_mem_pkt_v_o,
  data_mem_pkt_o,
  data_mem_pkt_yumi_i
);

  input [38:0] miss_addr_i;
  input [517:0] lce_data_cmd_i;
  output [522:0] data_mem_pkt_o;
  input clk_i;
  input reset_i;
  input lce_data_cmd_v_i;
  input data_mem_pkt_yumi_i;
  output cce_data_received_o;
  output tr_data_received_o;
  output uncached_data_received_o;
  output lce_data_cmd_ready_o;
  output data_mem_pkt_v_o;
  wire [522:0] data_mem_pkt_o;
  wire cce_data_received_o,tr_data_received_o,uncached_data_received_o,
  lce_data_cmd_ready_o,data_mem_pkt_v_o,lce_data_cmd_li_dst_id__0_,lce_data_cmd_li_msg_type__1_,
  lce_data_cmd_li_msg_type__0_,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9;
  assign data_mem_pkt_o[0] = 1'b0;
  assign data_mem_pkt_o[522] = miss_addr_i[11];
  assign data_mem_pkt_o[521] = miss_addr_i[10];
  assign data_mem_pkt_o[520] = miss_addr_i[9];
  assign data_mem_pkt_o[519] = miss_addr_i[8];
  assign data_mem_pkt_o[518] = miss_addr_i[7];
  assign data_mem_pkt_o[517] = miss_addr_i[6];

  bsg_two_fifo_width_p518
  rv_adapter
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(lce_data_cmd_ready_o),
    .data_i(lce_data_cmd_i),
    .v_i(lce_data_cmd_v_i),
    .v_o(data_mem_pkt_v_o),
    .data_o({ data_mem_pkt_o[513:2], lce_data_cmd_li_dst_id__0_, lce_data_cmd_li_msg_type__1_, lce_data_cmd_li_msg_type__0_, data_mem_pkt_o[516:514] }),
    .yumi_i(data_mem_pkt_yumi_i)
  );

  assign N0 = ~lce_data_cmd_li_msg_type__0_;
  assign N1 = N0 | lce_data_cmd_li_msg_type__1_;
  assign N2 = ~N1;
  assign N3 = lce_data_cmd_li_msg_type__0_ | lce_data_cmd_li_msg_type__1_;
  assign N4 = ~N3;
  assign N5 = ~lce_data_cmd_li_msg_type__1_;
  assign N6 = lce_data_cmd_li_msg_type__0_ | N5;
  assign N7 = ~N6;
  assign N8 = lce_data_cmd_li_msg_type__0_ | N5;
  assign N9 = ~N8;
  assign data_mem_pkt_o[1] = N9;
  assign cce_data_received_o = data_mem_pkt_yumi_i & N2;
  assign tr_data_received_o = data_mem_pkt_yumi_i & N4;
  assign uncached_data_received_o = data_mem_pkt_yumi_i & N7;

endmodule



module bp_fe_lce_02
(
  clk_i,
  reset_i,
  freeze_i,
  cfg_w_v_i,
  cfg_addr_i,
  cfg_data_i,
  id_i,
  ready_o,
  cache_miss_o,
  miss_i,
  miss_addr_i,
  uncached_req_i,
  data_mem_data_i,
  data_mem_pkt_o,
  data_mem_pkt_v_o,
  data_mem_pkt_yumi_i,
  tag_mem_pkt_o,
  tag_mem_pkt_v_o,
  tag_mem_pkt_yumi_i,
  stat_mem_pkt_v_o,
  stat_mem_pkt_o,
  lru_way_i,
  stat_mem_pkt_yumi_i,
  lce_req_o,
  lce_req_v_o,
  lce_req_ready_i,
  lce_resp_o,
  lce_resp_v_o,
  lce_resp_ready_i,
  lce_data_resp_o,
  lce_data_resp_v_o,
  lce_data_resp_ready_i,
  lce_cmd_i,
  lce_cmd_v_i,
  lce_cmd_ready_o,
  lce_data_cmd_i,
  lce_data_cmd_v_i,
  lce_data_cmd_ready_o,
  lce_data_cmd_o,
  lce_data_cmd_v_o,
  lce_data_cmd_ready_i,
  lce_mode_o
);

  input [15:0] cfg_addr_i;
  input [31:0] cfg_data_i;
  input [0:0] id_i;
  input [38:0] miss_addr_i;
  input [511:0] data_mem_data_i;
  output [522:0] data_mem_pkt_o;
  output [39:0] tag_mem_pkt_o;
  output [9:0] stat_mem_pkt_o;
  input [2:0] lru_way_i;
  output [113:0] lce_req_o;
  output [42:0] lce_resp_o;
  output [553:0] lce_data_resp_o;
  input [52:0] lce_cmd_i;
  input [517:0] lce_data_cmd_i;
  output [517:0] lce_data_cmd_o;
  input clk_i;
  input reset_i;
  input freeze_i;
  input cfg_w_v_i;
  input miss_i;
  input uncached_req_i;
  input data_mem_pkt_yumi_i;
  input tag_mem_pkt_yumi_i;
  input stat_mem_pkt_yumi_i;
  input lce_req_ready_i;
  input lce_resp_ready_i;
  input lce_data_resp_ready_i;
  input lce_cmd_v_i;
  input lce_data_cmd_v_i;
  input lce_data_cmd_ready_i;
  output ready_o;
  output cache_miss_o;
  output data_mem_pkt_v_o;
  output tag_mem_pkt_v_o;
  output stat_mem_pkt_v_o;
  output lce_req_v_o;
  output lce_resp_v_o;
  output lce_data_resp_v_o;
  output lce_cmd_ready_o;
  output lce_data_cmd_ready_o;
  output lce_data_cmd_v_o;
  output lce_mode_o;
  wire [522:0] data_mem_pkt_o,lce_cmd_data_mem_pkt_lo,lce_data_cmd_data_mem_pkt_lo;
  wire [39:0] tag_mem_pkt_o;
  wire [9:0] stat_mem_pkt_o;
  wire [113:0] lce_req_o;
  wire [42:0] lce_resp_o,lce_req_lce_resp_lo,lce_cmd_lce_resp_lo;
  wire [553:0] lce_data_resp_o;
  wire [517:0] lce_data_cmd_o;
  wire ready_o,cache_miss_o,data_mem_pkt_v_o,tag_mem_pkt_v_o,stat_mem_pkt_v_o,
  lce_req_v_o,lce_resp_v_o,lce_data_resp_v_o,lce_cmd_ready_o,lce_data_cmd_ready_o,
  lce_data_cmd_v_o,N0,N1,N2,N3,N4,N5,N6,lce_mode_w_v,N7,N8,N9,N10,N11,N12,N13,
  tr_data_received,cce_data_received,uncached_data_received,set_tag_received,
  set_tag_wakeup_received,lce_req_lce_resp_v_lo,lce_req_lce_resp_yumi_li,lce_ready_lo,
  lce_cmd_data_mem_pkt_v_lo,lce_cmd_data_mem_pkt_yumi_li,lce_cmd_lce_resp_v_lo,
  lce_cmd_lce_resp_yumi_li,lce_data_cmd_data_mem_pkt_v_lo,lce_data_cmd_data_mem_pkt_yumi_li,N14,
  N15,N16,N17,lce_ready,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,
  N33,N34,N35,N36,N37,N38,N39,N40;
  wire [38:0] miss_addr_lo;
  reg lce_mode_o;

  bp_fe_lce_req_02
  lce_req_inst
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .id_i(id_i[0]),
    .miss_i(miss_i),
    .miss_addr_i(miss_addr_i),
    .lru_way_i(lru_way_i),
    .uncached_req_i(uncached_req_i),
    .cache_miss_o(cache_miss_o),
    .miss_addr_o(miss_addr_lo),
    .tr_data_received_i(tr_data_received),
    .cce_data_received_i(cce_data_received),
    .uncached_data_received_i(uncached_data_received),
    .set_tag_received_i(set_tag_received),
    .set_tag_wakeup_received_i(set_tag_wakeup_received),
    .lce_req_o(lce_req_o),
    .lce_req_v_o(lce_req_v_o),
    .lce_req_ready_i(lce_req_ready_i),
    .lce_resp_o(lce_req_lce_resp_lo),
    .lce_resp_v_o(lce_req_lce_resp_v_lo),
    .lce_resp_yumi_i(lce_req_lce_resp_yumi_li)
  );


  bp_fe_lce_cmd_02
  lce_cmd_inst
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .id_i(id_i[0]),
    .lce_ready_o(lce_ready_lo),
    .set_tag_received_o(set_tag_received),
    .set_tag_wakeup_received_o(set_tag_wakeup_received),
    .data_mem_data_i(data_mem_data_i),
    .data_mem_pkt_o(lce_cmd_data_mem_pkt_lo),
    .data_mem_pkt_v_o(lce_cmd_data_mem_pkt_v_lo),
    .data_mem_pkt_yumi_i(lce_cmd_data_mem_pkt_yumi_li),
    .tag_mem_pkt_o(tag_mem_pkt_o),
    .tag_mem_pkt_v_o(tag_mem_pkt_v_o),
    .tag_mem_pkt_yumi_i(tag_mem_pkt_yumi_i),
    .stat_mem_pkt_v_o(stat_mem_pkt_v_o),
    .stat_mem_pkt_o(stat_mem_pkt_o),
    .stat_mem_pkt_yumi_i(stat_mem_pkt_yumi_i),
    .lce_resp_o(lce_cmd_lce_resp_lo),
    .lce_resp_v_o(lce_cmd_lce_resp_v_lo),
    .lce_resp_yumi_i(lce_cmd_lce_resp_yumi_li),
    .lce_data_resp_o(lce_data_resp_o),
    .lce_data_resp_v_o(lce_data_resp_v_o),
    .lce_data_resp_ready_i(lce_data_resp_ready_i),
    .lce_cmd_i(lce_cmd_i),
    .lce_cmd_v_i(lce_cmd_v_i),
    .lce_cmd_ready_o(lce_cmd_ready_o),
    .lce_data_cmd_o(lce_data_cmd_o),
    .lce_data_cmd_v_o(lce_data_cmd_v_o),
    .lce_data_cmd_ready_i(lce_data_cmd_ready_i)
  );


  bp_fe_lce_data_cmd_02
  lce_data_cmd
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .cce_data_received_o(cce_data_received),
    .tr_data_received_o(tr_data_received),
    .uncached_data_received_o(uncached_data_received),
    .miss_addr_i(miss_addr_lo),
    .lce_data_cmd_i(lce_data_cmd_i),
    .lce_data_cmd_v_i(lce_data_cmd_v_i),
    .lce_data_cmd_ready_o(lce_data_cmd_ready_o),
    .data_mem_pkt_v_o(lce_data_cmd_data_mem_pkt_v_lo),
    .data_mem_pkt_o(lce_data_cmd_data_mem_pkt_lo),
    .data_mem_pkt_yumi_i(lce_data_cmd_data_mem_pkt_yumi_li)
  );

  assign N18 = ~lce_mode_o;
  assign N19 = ~cfg_addr_i[5];
  assign N20 = ~cfg_addr_i[1];
  assign N21 = cfg_addr_i[14] | cfg_addr_i[15];
  assign N22 = cfg_addr_i[13] | N21;
  assign N23 = cfg_addr_i[12] | N22;
  assign N24 = cfg_addr_i[11] | N23;
  assign N25 = cfg_addr_i[10] | N24;
  assign N26 = cfg_addr_i[9] | N25;
  assign N27 = cfg_addr_i[8] | N26;
  assign N28 = cfg_addr_i[7] | N27;
  assign N29 = cfg_addr_i[6] | N28;
  assign N30 = N19 | N29;
  assign N31 = cfg_addr_i[4] | N30;
  assign N32 = cfg_addr_i[3] | N31;
  assign N33 = cfg_addr_i[2] | N32;
  assign N34 = N20 | N33;
  assign N35 = cfg_addr_i[0] | N34;
  assign N36 = ~N35;
  assign N10 = (N0)? 1'b1 : 
               (N13)? 1'b1 : 
               (N9)? 1'b0 : 1'b0;
  assign N0 = N7;
  assign N11 = (N0)? 1'b0 : 
               (N13)? cfg_data_i[0] : 1'b0;
  assign data_mem_pkt_v_o = (N1)? 1'b1 : 
                            (N2)? lce_cmd_data_mem_pkt_v_lo : 1'b0;
  assign N1 = lce_data_cmd_data_mem_pkt_v_lo;
  assign N2 = N14;
  assign data_mem_pkt_o = (N1)? lce_data_cmd_data_mem_pkt_lo : 
                          (N2)? lce_cmd_data_mem_pkt_lo : 1'b0;
  assign lce_data_cmd_data_mem_pkt_yumi_li = (N1)? data_mem_pkt_yumi_i : 
                                             (N2)? 1'b0 : 1'b0;
  assign lce_cmd_data_mem_pkt_yumi_li = (N1)? 1'b0 : 
                                        (N2)? data_mem_pkt_yumi_i : 1'b0;
  assign lce_resp_v_o = (N3)? 1'b1 : 
                        (N4)? lce_cmd_lce_resp_v_lo : 1'b0;
  assign N3 = lce_req_lce_resp_v_lo;
  assign N4 = N15;
  assign lce_resp_o = (N3)? lce_req_lce_resp_lo : 
                      (N4)? lce_cmd_lce_resp_lo : 1'b0;
  assign lce_req_lce_resp_yumi_li = (N3)? lce_resp_ready_i : 
                                    (N4)? 1'b0 : 1'b0;
  assign lce_cmd_lce_resp_yumi_li = (N3)? 1'b0 : 
                                    (N4)? N16 : 1'b0;
  assign lce_ready = (N5)? N17 : 
                     (N6)? lce_ready_lo : 1'b0;
  assign N5 = N18;
  assign N6 = lce_mode_o;
  assign lce_mode_w_v = N37 & N36;
  assign N37 = freeze_i & cfg_w_v_i;
  assign N7 = reset_i;
  assign N8 = lce_mode_w_v | N7;
  assign N9 = ~N8;
  assign N12 = ~N7;
  assign N13 = lce_mode_w_v & N12;
  assign N14 = ~lce_data_cmd_data_mem_pkt_v_lo;
  assign N15 = ~lce_req_lce_resp_v_lo;
  assign N16 = lce_cmd_lce_resp_v_lo & lce_resp_ready_i;
  assign N17 = ~freeze_i;
  assign ready_o = N39 & N40;
  assign N39 = lce_ready & N38;
  assign N38 = ~1'b0;
  assign N40 = ~cache_miss_o;

  always @(posedge clk_i) begin
    if(N10) begin
      lce_mode_o <= N11;
    end 
  end


endmodule



module bsg_mux_width_p64_els_p8
(
  data_i,
  sel_i,
  data_o
);

  input [511:0] data_i;
  input [2:0] sel_i;
  output [63:0] data_o;
  wire [63:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14;
  assign data_o[63] = (N7)? data_i[63] : 
                      (N9)? data_i[127] : 
                      (N11)? data_i[191] : 
                      (N13)? data_i[255] : 
                      (N8)? data_i[319] : 
                      (N10)? data_i[383] : 
                      (N12)? data_i[447] : 
                      (N14)? data_i[511] : 1'b0;
  assign data_o[62] = (N7)? data_i[62] : 
                      (N9)? data_i[126] : 
                      (N11)? data_i[190] : 
                      (N13)? data_i[254] : 
                      (N8)? data_i[318] : 
                      (N10)? data_i[382] : 
                      (N12)? data_i[446] : 
                      (N14)? data_i[510] : 1'b0;
  assign data_o[61] = (N7)? data_i[61] : 
                      (N9)? data_i[125] : 
                      (N11)? data_i[189] : 
                      (N13)? data_i[253] : 
                      (N8)? data_i[317] : 
                      (N10)? data_i[381] : 
                      (N12)? data_i[445] : 
                      (N14)? data_i[509] : 1'b0;
  assign data_o[60] = (N7)? data_i[60] : 
                      (N9)? data_i[124] : 
                      (N11)? data_i[188] : 
                      (N13)? data_i[252] : 
                      (N8)? data_i[316] : 
                      (N10)? data_i[380] : 
                      (N12)? data_i[444] : 
                      (N14)? data_i[508] : 1'b0;
  assign data_o[59] = (N7)? data_i[59] : 
                      (N9)? data_i[123] : 
                      (N11)? data_i[187] : 
                      (N13)? data_i[251] : 
                      (N8)? data_i[315] : 
                      (N10)? data_i[379] : 
                      (N12)? data_i[443] : 
                      (N14)? data_i[507] : 1'b0;
  assign data_o[58] = (N7)? data_i[58] : 
                      (N9)? data_i[122] : 
                      (N11)? data_i[186] : 
                      (N13)? data_i[250] : 
                      (N8)? data_i[314] : 
                      (N10)? data_i[378] : 
                      (N12)? data_i[442] : 
                      (N14)? data_i[506] : 1'b0;
  assign data_o[57] = (N7)? data_i[57] : 
                      (N9)? data_i[121] : 
                      (N11)? data_i[185] : 
                      (N13)? data_i[249] : 
                      (N8)? data_i[313] : 
                      (N10)? data_i[377] : 
                      (N12)? data_i[441] : 
                      (N14)? data_i[505] : 1'b0;
  assign data_o[56] = (N7)? data_i[56] : 
                      (N9)? data_i[120] : 
                      (N11)? data_i[184] : 
                      (N13)? data_i[248] : 
                      (N8)? data_i[312] : 
                      (N10)? data_i[376] : 
                      (N12)? data_i[440] : 
                      (N14)? data_i[504] : 1'b0;
  assign data_o[55] = (N7)? data_i[55] : 
                      (N9)? data_i[119] : 
                      (N11)? data_i[183] : 
                      (N13)? data_i[247] : 
                      (N8)? data_i[311] : 
                      (N10)? data_i[375] : 
                      (N12)? data_i[439] : 
                      (N14)? data_i[503] : 1'b0;
  assign data_o[54] = (N7)? data_i[54] : 
                      (N9)? data_i[118] : 
                      (N11)? data_i[182] : 
                      (N13)? data_i[246] : 
                      (N8)? data_i[310] : 
                      (N10)? data_i[374] : 
                      (N12)? data_i[438] : 
                      (N14)? data_i[502] : 1'b0;
  assign data_o[53] = (N7)? data_i[53] : 
                      (N9)? data_i[117] : 
                      (N11)? data_i[181] : 
                      (N13)? data_i[245] : 
                      (N8)? data_i[309] : 
                      (N10)? data_i[373] : 
                      (N12)? data_i[437] : 
                      (N14)? data_i[501] : 1'b0;
  assign data_o[52] = (N7)? data_i[52] : 
                      (N9)? data_i[116] : 
                      (N11)? data_i[180] : 
                      (N13)? data_i[244] : 
                      (N8)? data_i[308] : 
                      (N10)? data_i[372] : 
                      (N12)? data_i[436] : 
                      (N14)? data_i[500] : 1'b0;
  assign data_o[51] = (N7)? data_i[51] : 
                      (N9)? data_i[115] : 
                      (N11)? data_i[179] : 
                      (N13)? data_i[243] : 
                      (N8)? data_i[307] : 
                      (N10)? data_i[371] : 
                      (N12)? data_i[435] : 
                      (N14)? data_i[499] : 1'b0;
  assign data_o[50] = (N7)? data_i[50] : 
                      (N9)? data_i[114] : 
                      (N11)? data_i[178] : 
                      (N13)? data_i[242] : 
                      (N8)? data_i[306] : 
                      (N10)? data_i[370] : 
                      (N12)? data_i[434] : 
                      (N14)? data_i[498] : 1'b0;
  assign data_o[49] = (N7)? data_i[49] : 
                      (N9)? data_i[113] : 
                      (N11)? data_i[177] : 
                      (N13)? data_i[241] : 
                      (N8)? data_i[305] : 
                      (N10)? data_i[369] : 
                      (N12)? data_i[433] : 
                      (N14)? data_i[497] : 1'b0;
  assign data_o[48] = (N7)? data_i[48] : 
                      (N9)? data_i[112] : 
                      (N11)? data_i[176] : 
                      (N13)? data_i[240] : 
                      (N8)? data_i[304] : 
                      (N10)? data_i[368] : 
                      (N12)? data_i[432] : 
                      (N14)? data_i[496] : 1'b0;
  assign data_o[47] = (N7)? data_i[47] : 
                      (N9)? data_i[111] : 
                      (N11)? data_i[175] : 
                      (N13)? data_i[239] : 
                      (N8)? data_i[303] : 
                      (N10)? data_i[367] : 
                      (N12)? data_i[431] : 
                      (N14)? data_i[495] : 1'b0;
  assign data_o[46] = (N7)? data_i[46] : 
                      (N9)? data_i[110] : 
                      (N11)? data_i[174] : 
                      (N13)? data_i[238] : 
                      (N8)? data_i[302] : 
                      (N10)? data_i[366] : 
                      (N12)? data_i[430] : 
                      (N14)? data_i[494] : 1'b0;
  assign data_o[45] = (N7)? data_i[45] : 
                      (N9)? data_i[109] : 
                      (N11)? data_i[173] : 
                      (N13)? data_i[237] : 
                      (N8)? data_i[301] : 
                      (N10)? data_i[365] : 
                      (N12)? data_i[429] : 
                      (N14)? data_i[493] : 1'b0;
  assign data_o[44] = (N7)? data_i[44] : 
                      (N9)? data_i[108] : 
                      (N11)? data_i[172] : 
                      (N13)? data_i[236] : 
                      (N8)? data_i[300] : 
                      (N10)? data_i[364] : 
                      (N12)? data_i[428] : 
                      (N14)? data_i[492] : 1'b0;
  assign data_o[43] = (N7)? data_i[43] : 
                      (N9)? data_i[107] : 
                      (N11)? data_i[171] : 
                      (N13)? data_i[235] : 
                      (N8)? data_i[299] : 
                      (N10)? data_i[363] : 
                      (N12)? data_i[427] : 
                      (N14)? data_i[491] : 1'b0;
  assign data_o[42] = (N7)? data_i[42] : 
                      (N9)? data_i[106] : 
                      (N11)? data_i[170] : 
                      (N13)? data_i[234] : 
                      (N8)? data_i[298] : 
                      (N10)? data_i[362] : 
                      (N12)? data_i[426] : 
                      (N14)? data_i[490] : 1'b0;
  assign data_o[41] = (N7)? data_i[41] : 
                      (N9)? data_i[105] : 
                      (N11)? data_i[169] : 
                      (N13)? data_i[233] : 
                      (N8)? data_i[297] : 
                      (N10)? data_i[361] : 
                      (N12)? data_i[425] : 
                      (N14)? data_i[489] : 1'b0;
  assign data_o[40] = (N7)? data_i[40] : 
                      (N9)? data_i[104] : 
                      (N11)? data_i[168] : 
                      (N13)? data_i[232] : 
                      (N8)? data_i[296] : 
                      (N10)? data_i[360] : 
                      (N12)? data_i[424] : 
                      (N14)? data_i[488] : 1'b0;
  assign data_o[39] = (N7)? data_i[39] : 
                      (N9)? data_i[103] : 
                      (N11)? data_i[167] : 
                      (N13)? data_i[231] : 
                      (N8)? data_i[295] : 
                      (N10)? data_i[359] : 
                      (N12)? data_i[423] : 
                      (N14)? data_i[487] : 1'b0;
  assign data_o[38] = (N7)? data_i[38] : 
                      (N9)? data_i[102] : 
                      (N11)? data_i[166] : 
                      (N13)? data_i[230] : 
                      (N8)? data_i[294] : 
                      (N10)? data_i[358] : 
                      (N12)? data_i[422] : 
                      (N14)? data_i[486] : 1'b0;
  assign data_o[37] = (N7)? data_i[37] : 
                      (N9)? data_i[101] : 
                      (N11)? data_i[165] : 
                      (N13)? data_i[229] : 
                      (N8)? data_i[293] : 
                      (N10)? data_i[357] : 
                      (N12)? data_i[421] : 
                      (N14)? data_i[485] : 1'b0;
  assign data_o[36] = (N7)? data_i[36] : 
                      (N9)? data_i[100] : 
                      (N11)? data_i[164] : 
                      (N13)? data_i[228] : 
                      (N8)? data_i[292] : 
                      (N10)? data_i[356] : 
                      (N12)? data_i[420] : 
                      (N14)? data_i[484] : 1'b0;
  assign data_o[35] = (N7)? data_i[35] : 
                      (N9)? data_i[99] : 
                      (N11)? data_i[163] : 
                      (N13)? data_i[227] : 
                      (N8)? data_i[291] : 
                      (N10)? data_i[355] : 
                      (N12)? data_i[419] : 
                      (N14)? data_i[483] : 1'b0;
  assign data_o[34] = (N7)? data_i[34] : 
                      (N9)? data_i[98] : 
                      (N11)? data_i[162] : 
                      (N13)? data_i[226] : 
                      (N8)? data_i[290] : 
                      (N10)? data_i[354] : 
                      (N12)? data_i[418] : 
                      (N14)? data_i[482] : 1'b0;
  assign data_o[33] = (N7)? data_i[33] : 
                      (N9)? data_i[97] : 
                      (N11)? data_i[161] : 
                      (N13)? data_i[225] : 
                      (N8)? data_i[289] : 
                      (N10)? data_i[353] : 
                      (N12)? data_i[417] : 
                      (N14)? data_i[481] : 1'b0;
  assign data_o[32] = (N7)? data_i[32] : 
                      (N9)? data_i[96] : 
                      (N11)? data_i[160] : 
                      (N13)? data_i[224] : 
                      (N8)? data_i[288] : 
                      (N10)? data_i[352] : 
                      (N12)? data_i[416] : 
                      (N14)? data_i[480] : 1'b0;
  assign data_o[31] = (N7)? data_i[31] : 
                      (N9)? data_i[95] : 
                      (N11)? data_i[159] : 
                      (N13)? data_i[223] : 
                      (N8)? data_i[287] : 
                      (N10)? data_i[351] : 
                      (N12)? data_i[415] : 
                      (N14)? data_i[479] : 1'b0;
  assign data_o[30] = (N7)? data_i[30] : 
                      (N9)? data_i[94] : 
                      (N11)? data_i[158] : 
                      (N13)? data_i[222] : 
                      (N8)? data_i[286] : 
                      (N10)? data_i[350] : 
                      (N12)? data_i[414] : 
                      (N14)? data_i[478] : 1'b0;
  assign data_o[29] = (N7)? data_i[29] : 
                      (N9)? data_i[93] : 
                      (N11)? data_i[157] : 
                      (N13)? data_i[221] : 
                      (N8)? data_i[285] : 
                      (N10)? data_i[349] : 
                      (N12)? data_i[413] : 
                      (N14)? data_i[477] : 1'b0;
  assign data_o[28] = (N7)? data_i[28] : 
                      (N9)? data_i[92] : 
                      (N11)? data_i[156] : 
                      (N13)? data_i[220] : 
                      (N8)? data_i[284] : 
                      (N10)? data_i[348] : 
                      (N12)? data_i[412] : 
                      (N14)? data_i[476] : 1'b0;
  assign data_o[27] = (N7)? data_i[27] : 
                      (N9)? data_i[91] : 
                      (N11)? data_i[155] : 
                      (N13)? data_i[219] : 
                      (N8)? data_i[283] : 
                      (N10)? data_i[347] : 
                      (N12)? data_i[411] : 
                      (N14)? data_i[475] : 1'b0;
  assign data_o[26] = (N7)? data_i[26] : 
                      (N9)? data_i[90] : 
                      (N11)? data_i[154] : 
                      (N13)? data_i[218] : 
                      (N8)? data_i[282] : 
                      (N10)? data_i[346] : 
                      (N12)? data_i[410] : 
                      (N14)? data_i[474] : 1'b0;
  assign data_o[25] = (N7)? data_i[25] : 
                      (N9)? data_i[89] : 
                      (N11)? data_i[153] : 
                      (N13)? data_i[217] : 
                      (N8)? data_i[281] : 
                      (N10)? data_i[345] : 
                      (N12)? data_i[409] : 
                      (N14)? data_i[473] : 1'b0;
  assign data_o[24] = (N7)? data_i[24] : 
                      (N9)? data_i[88] : 
                      (N11)? data_i[152] : 
                      (N13)? data_i[216] : 
                      (N8)? data_i[280] : 
                      (N10)? data_i[344] : 
                      (N12)? data_i[408] : 
                      (N14)? data_i[472] : 1'b0;
  assign data_o[23] = (N7)? data_i[23] : 
                      (N9)? data_i[87] : 
                      (N11)? data_i[151] : 
                      (N13)? data_i[215] : 
                      (N8)? data_i[279] : 
                      (N10)? data_i[343] : 
                      (N12)? data_i[407] : 
                      (N14)? data_i[471] : 1'b0;
  assign data_o[22] = (N7)? data_i[22] : 
                      (N9)? data_i[86] : 
                      (N11)? data_i[150] : 
                      (N13)? data_i[214] : 
                      (N8)? data_i[278] : 
                      (N10)? data_i[342] : 
                      (N12)? data_i[406] : 
                      (N14)? data_i[470] : 1'b0;
  assign data_o[21] = (N7)? data_i[21] : 
                      (N9)? data_i[85] : 
                      (N11)? data_i[149] : 
                      (N13)? data_i[213] : 
                      (N8)? data_i[277] : 
                      (N10)? data_i[341] : 
                      (N12)? data_i[405] : 
                      (N14)? data_i[469] : 1'b0;
  assign data_o[20] = (N7)? data_i[20] : 
                      (N9)? data_i[84] : 
                      (N11)? data_i[148] : 
                      (N13)? data_i[212] : 
                      (N8)? data_i[276] : 
                      (N10)? data_i[340] : 
                      (N12)? data_i[404] : 
                      (N14)? data_i[468] : 1'b0;
  assign data_o[19] = (N7)? data_i[19] : 
                      (N9)? data_i[83] : 
                      (N11)? data_i[147] : 
                      (N13)? data_i[211] : 
                      (N8)? data_i[275] : 
                      (N10)? data_i[339] : 
                      (N12)? data_i[403] : 
                      (N14)? data_i[467] : 1'b0;
  assign data_o[18] = (N7)? data_i[18] : 
                      (N9)? data_i[82] : 
                      (N11)? data_i[146] : 
                      (N13)? data_i[210] : 
                      (N8)? data_i[274] : 
                      (N10)? data_i[338] : 
                      (N12)? data_i[402] : 
                      (N14)? data_i[466] : 1'b0;
  assign data_o[17] = (N7)? data_i[17] : 
                      (N9)? data_i[81] : 
                      (N11)? data_i[145] : 
                      (N13)? data_i[209] : 
                      (N8)? data_i[273] : 
                      (N10)? data_i[337] : 
                      (N12)? data_i[401] : 
                      (N14)? data_i[465] : 1'b0;
  assign data_o[16] = (N7)? data_i[16] : 
                      (N9)? data_i[80] : 
                      (N11)? data_i[144] : 
                      (N13)? data_i[208] : 
                      (N8)? data_i[272] : 
                      (N10)? data_i[336] : 
                      (N12)? data_i[400] : 
                      (N14)? data_i[464] : 1'b0;
  assign data_o[15] = (N7)? data_i[15] : 
                      (N9)? data_i[79] : 
                      (N11)? data_i[143] : 
                      (N13)? data_i[207] : 
                      (N8)? data_i[271] : 
                      (N10)? data_i[335] : 
                      (N12)? data_i[399] : 
                      (N14)? data_i[463] : 1'b0;
  assign data_o[14] = (N7)? data_i[14] : 
                      (N9)? data_i[78] : 
                      (N11)? data_i[142] : 
                      (N13)? data_i[206] : 
                      (N8)? data_i[270] : 
                      (N10)? data_i[334] : 
                      (N12)? data_i[398] : 
                      (N14)? data_i[462] : 1'b0;
  assign data_o[13] = (N7)? data_i[13] : 
                      (N9)? data_i[77] : 
                      (N11)? data_i[141] : 
                      (N13)? data_i[205] : 
                      (N8)? data_i[269] : 
                      (N10)? data_i[333] : 
                      (N12)? data_i[397] : 
                      (N14)? data_i[461] : 1'b0;
  assign data_o[12] = (N7)? data_i[12] : 
                      (N9)? data_i[76] : 
                      (N11)? data_i[140] : 
                      (N13)? data_i[204] : 
                      (N8)? data_i[268] : 
                      (N10)? data_i[332] : 
                      (N12)? data_i[396] : 
                      (N14)? data_i[460] : 1'b0;
  assign data_o[11] = (N7)? data_i[11] : 
                      (N9)? data_i[75] : 
                      (N11)? data_i[139] : 
                      (N13)? data_i[203] : 
                      (N8)? data_i[267] : 
                      (N10)? data_i[331] : 
                      (N12)? data_i[395] : 
                      (N14)? data_i[459] : 1'b0;
  assign data_o[10] = (N7)? data_i[10] : 
                      (N9)? data_i[74] : 
                      (N11)? data_i[138] : 
                      (N13)? data_i[202] : 
                      (N8)? data_i[266] : 
                      (N10)? data_i[330] : 
                      (N12)? data_i[394] : 
                      (N14)? data_i[458] : 1'b0;
  assign data_o[9] = (N7)? data_i[9] : 
                     (N9)? data_i[73] : 
                     (N11)? data_i[137] : 
                     (N13)? data_i[201] : 
                     (N8)? data_i[265] : 
                     (N10)? data_i[329] : 
                     (N12)? data_i[393] : 
                     (N14)? data_i[457] : 1'b0;
  assign data_o[8] = (N7)? data_i[8] : 
                     (N9)? data_i[72] : 
                     (N11)? data_i[136] : 
                     (N13)? data_i[200] : 
                     (N8)? data_i[264] : 
                     (N10)? data_i[328] : 
                     (N12)? data_i[392] : 
                     (N14)? data_i[456] : 1'b0;
  assign data_o[7] = (N7)? data_i[7] : 
                     (N9)? data_i[71] : 
                     (N11)? data_i[135] : 
                     (N13)? data_i[199] : 
                     (N8)? data_i[263] : 
                     (N10)? data_i[327] : 
                     (N12)? data_i[391] : 
                     (N14)? data_i[455] : 1'b0;
  assign data_o[6] = (N7)? data_i[6] : 
                     (N9)? data_i[70] : 
                     (N11)? data_i[134] : 
                     (N13)? data_i[198] : 
                     (N8)? data_i[262] : 
                     (N10)? data_i[326] : 
                     (N12)? data_i[390] : 
                     (N14)? data_i[454] : 1'b0;
  assign data_o[5] = (N7)? data_i[5] : 
                     (N9)? data_i[69] : 
                     (N11)? data_i[133] : 
                     (N13)? data_i[197] : 
                     (N8)? data_i[261] : 
                     (N10)? data_i[325] : 
                     (N12)? data_i[389] : 
                     (N14)? data_i[453] : 1'b0;
  assign data_o[4] = (N7)? data_i[4] : 
                     (N9)? data_i[68] : 
                     (N11)? data_i[132] : 
                     (N13)? data_i[196] : 
                     (N8)? data_i[260] : 
                     (N10)? data_i[324] : 
                     (N12)? data_i[388] : 
                     (N14)? data_i[452] : 1'b0;
  assign data_o[3] = (N7)? data_i[3] : 
                     (N9)? data_i[67] : 
                     (N11)? data_i[131] : 
                     (N13)? data_i[195] : 
                     (N8)? data_i[259] : 
                     (N10)? data_i[323] : 
                     (N12)? data_i[387] : 
                     (N14)? data_i[451] : 1'b0;
  assign data_o[2] = (N7)? data_i[2] : 
                     (N9)? data_i[66] : 
                     (N11)? data_i[130] : 
                     (N13)? data_i[194] : 
                     (N8)? data_i[258] : 
                     (N10)? data_i[322] : 
                     (N12)? data_i[386] : 
                     (N14)? data_i[450] : 1'b0;
  assign data_o[1] = (N7)? data_i[1] : 
                     (N9)? data_i[65] : 
                     (N11)? data_i[129] : 
                     (N13)? data_i[193] : 
                     (N8)? data_i[257] : 
                     (N10)? data_i[321] : 
                     (N12)? data_i[385] : 
                     (N14)? data_i[449] : 1'b0;
  assign data_o[0] = (N7)? data_i[0] : 
                     (N9)? data_i[64] : 
                     (N11)? data_i[128] : 
                     (N13)? data_i[192] : 
                     (N8)? data_i[256] : 
                     (N10)? data_i[320] : 
                     (N12)? data_i[384] : 
                     (N14)? data_i[448] : 1'b0;
  assign N0 = ~sel_i[0];
  assign N1 = ~sel_i[1];
  assign N2 = N0 & N1;
  assign N3 = N0 & sel_i[1];
  assign N4 = sel_i[0] & N1;
  assign N5 = sel_i[0] & sel_i[1];
  assign N6 = ~sel_i[2];
  assign N7 = N2 & N6;
  assign N8 = N2 & sel_i[2];
  assign N9 = N4 & N6;
  assign N10 = N4 & sel_i[2];
  assign N11 = N3 & N6;
  assign N12 = N3 & sel_i[2];
  assign N13 = N5 & N6;
  assign N14 = N5 & sel_i[2];

endmodule



module bsg_mux_width_p64_els_p2
(
  data_i,
  sel_i,
  data_o
);

  input [127:0] data_i;
  input [0:0] sel_i;
  output [63:0] data_o;
  wire [63:0] data_o;
  wire N0,N1;
  assign data_o[63] = (N1)? data_i[63] : 
                      (N0)? data_i[127] : 1'b0;
  assign N0 = sel_i[0];
  assign data_o[62] = (N1)? data_i[62] : 
                      (N0)? data_i[126] : 1'b0;
  assign data_o[61] = (N1)? data_i[61] : 
                      (N0)? data_i[125] : 1'b0;
  assign data_o[60] = (N1)? data_i[60] : 
                      (N0)? data_i[124] : 1'b0;
  assign data_o[59] = (N1)? data_i[59] : 
                      (N0)? data_i[123] : 1'b0;
  assign data_o[58] = (N1)? data_i[58] : 
                      (N0)? data_i[122] : 1'b0;
  assign data_o[57] = (N1)? data_i[57] : 
                      (N0)? data_i[121] : 1'b0;
  assign data_o[56] = (N1)? data_i[56] : 
                      (N0)? data_i[120] : 1'b0;
  assign data_o[55] = (N1)? data_i[55] : 
                      (N0)? data_i[119] : 1'b0;
  assign data_o[54] = (N1)? data_i[54] : 
                      (N0)? data_i[118] : 1'b0;
  assign data_o[53] = (N1)? data_i[53] : 
                      (N0)? data_i[117] : 1'b0;
  assign data_o[52] = (N1)? data_i[52] : 
                      (N0)? data_i[116] : 1'b0;
  assign data_o[51] = (N1)? data_i[51] : 
                      (N0)? data_i[115] : 1'b0;
  assign data_o[50] = (N1)? data_i[50] : 
                      (N0)? data_i[114] : 1'b0;
  assign data_o[49] = (N1)? data_i[49] : 
                      (N0)? data_i[113] : 1'b0;
  assign data_o[48] = (N1)? data_i[48] : 
                      (N0)? data_i[112] : 1'b0;
  assign data_o[47] = (N1)? data_i[47] : 
                      (N0)? data_i[111] : 1'b0;
  assign data_o[46] = (N1)? data_i[46] : 
                      (N0)? data_i[110] : 1'b0;
  assign data_o[45] = (N1)? data_i[45] : 
                      (N0)? data_i[109] : 1'b0;
  assign data_o[44] = (N1)? data_i[44] : 
                      (N0)? data_i[108] : 1'b0;
  assign data_o[43] = (N1)? data_i[43] : 
                      (N0)? data_i[107] : 1'b0;
  assign data_o[42] = (N1)? data_i[42] : 
                      (N0)? data_i[106] : 1'b0;
  assign data_o[41] = (N1)? data_i[41] : 
                      (N0)? data_i[105] : 1'b0;
  assign data_o[40] = (N1)? data_i[40] : 
                      (N0)? data_i[104] : 1'b0;
  assign data_o[39] = (N1)? data_i[39] : 
                      (N0)? data_i[103] : 1'b0;
  assign data_o[38] = (N1)? data_i[38] : 
                      (N0)? data_i[102] : 1'b0;
  assign data_o[37] = (N1)? data_i[37] : 
                      (N0)? data_i[101] : 1'b0;
  assign data_o[36] = (N1)? data_i[36] : 
                      (N0)? data_i[100] : 1'b0;
  assign data_o[35] = (N1)? data_i[35] : 
                      (N0)? data_i[99] : 1'b0;
  assign data_o[34] = (N1)? data_i[34] : 
                      (N0)? data_i[98] : 1'b0;
  assign data_o[33] = (N1)? data_i[33] : 
                      (N0)? data_i[97] : 1'b0;
  assign data_o[32] = (N1)? data_i[32] : 
                      (N0)? data_i[96] : 1'b0;
  assign data_o[31] = (N1)? data_i[31] : 
                      (N0)? data_i[95] : 1'b0;
  assign data_o[30] = (N1)? data_i[30] : 
                      (N0)? data_i[94] : 1'b0;
  assign data_o[29] = (N1)? data_i[29] : 
                      (N0)? data_i[93] : 1'b0;
  assign data_o[28] = (N1)? data_i[28] : 
                      (N0)? data_i[92] : 1'b0;
  assign data_o[27] = (N1)? data_i[27] : 
                      (N0)? data_i[91] : 1'b0;
  assign data_o[26] = (N1)? data_i[26] : 
                      (N0)? data_i[90] : 1'b0;
  assign data_o[25] = (N1)? data_i[25] : 
                      (N0)? data_i[89] : 1'b0;
  assign data_o[24] = (N1)? data_i[24] : 
                      (N0)? data_i[88] : 1'b0;
  assign data_o[23] = (N1)? data_i[23] : 
                      (N0)? data_i[87] : 1'b0;
  assign data_o[22] = (N1)? data_i[22] : 
                      (N0)? data_i[86] : 1'b0;
  assign data_o[21] = (N1)? data_i[21] : 
                      (N0)? data_i[85] : 1'b0;
  assign data_o[20] = (N1)? data_i[20] : 
                      (N0)? data_i[84] : 1'b0;
  assign data_o[19] = (N1)? data_i[19] : 
                      (N0)? data_i[83] : 1'b0;
  assign data_o[18] = (N1)? data_i[18] : 
                      (N0)? data_i[82] : 1'b0;
  assign data_o[17] = (N1)? data_i[17] : 
                      (N0)? data_i[81] : 1'b0;
  assign data_o[16] = (N1)? data_i[16] : 
                      (N0)? data_i[80] : 1'b0;
  assign data_o[15] = (N1)? data_i[15] : 
                      (N0)? data_i[79] : 1'b0;
  assign data_o[14] = (N1)? data_i[14] : 
                      (N0)? data_i[78] : 1'b0;
  assign data_o[13] = (N1)? data_i[13] : 
                      (N0)? data_i[77] : 1'b0;
  assign data_o[12] = (N1)? data_i[12] : 
                      (N0)? data_i[76] : 1'b0;
  assign data_o[11] = (N1)? data_i[11] : 
                      (N0)? data_i[75] : 1'b0;
  assign data_o[10] = (N1)? data_i[10] : 
                      (N0)? data_i[74] : 1'b0;
  assign data_o[9] = (N1)? data_i[9] : 
                     (N0)? data_i[73] : 1'b0;
  assign data_o[8] = (N1)? data_i[8] : 
                     (N0)? data_i[72] : 1'b0;
  assign data_o[7] = (N1)? data_i[7] : 
                     (N0)? data_i[71] : 1'b0;
  assign data_o[6] = (N1)? data_i[6] : 
                     (N0)? data_i[70] : 1'b0;
  assign data_o[5] = (N1)? data_i[5] : 
                     (N0)? data_i[69] : 1'b0;
  assign data_o[4] = (N1)? data_i[4] : 
                     (N0)? data_i[68] : 1'b0;
  assign data_o[3] = (N1)? data_i[3] : 
                     (N0)? data_i[67] : 1'b0;
  assign data_o[2] = (N1)? data_i[2] : 
                     (N0)? data_i[66] : 1'b0;
  assign data_o[1] = (N1)? data_i[1] : 
                     (N0)? data_i[65] : 1'b0;
  assign data_o[0] = (N1)? data_i[0] : 
                     (N0)? data_i[64] : 1'b0;
  assign N1 = ~sel_i[0];

endmodule



module bsg_swap_width_p64
(
  data_i,
  swap_i,
  data_o
);

  input [127:0] data_i;
  output [127:0] data_o;
  input swap_i;
  wire [127:0] data_o;
  wire N0,N1,N2;
  assign data_o = (N0)? { data_i[63:0], data_i[127:64] } : 
                  (N1)? data_i : 1'b0;
  assign N0 = swap_i;
  assign N1 = N2;
  assign N2 = ~swap_i;

endmodule



module bsg_swap_width_p128
(
  data_i,
  swap_i,
  data_o
);

  input [255:0] data_i;
  output [255:0] data_o;
  input swap_i;
  wire [255:0] data_o;
  wire N0,N1,N2;
  assign data_o = (N0)? { data_i[127:0], data_i[255:128] } : 
                  (N1)? data_i : 1'b0;
  assign N0 = swap_i;
  assign N1 = N2;
  assign N2 = ~swap_i;

endmodule



module bsg_swap_width_p256
(
  data_i,
  swap_i,
  data_o
);

  input [511:0] data_i;
  output [511:0] data_o;
  input swap_i;
  wire [511:0] data_o;
  wire N0,N1,N2;
  assign data_o = (N0)? { data_i[255:0], data_i[511:256] } : 
                  (N1)? data_i : 1'b0;
  assign N0 = swap_i;
  assign N1 = N2;
  assign N2 = ~swap_i;

endmodule



module bsg_mux_butterfly_width_p64_els_p8
(
  data_i,
  sel_i,
  data_o
);

  input [511:0] data_i;
  input [2:0] sel_i;
  output [511:0] data_o;
  wire [511:0] data_o;
  wire data_stage_1__511_,data_stage_1__510_,data_stage_1__509_,data_stage_1__508_,
  data_stage_1__507_,data_stage_1__506_,data_stage_1__505_,data_stage_1__504_,
  data_stage_1__503_,data_stage_1__502_,data_stage_1__501_,data_stage_1__500_,
  data_stage_1__499_,data_stage_1__498_,data_stage_1__497_,data_stage_1__496_,
  data_stage_1__495_,data_stage_1__494_,data_stage_1__493_,data_stage_1__492_,data_stage_1__491_,
  data_stage_1__490_,data_stage_1__489_,data_stage_1__488_,data_stage_1__487_,
  data_stage_1__486_,data_stage_1__485_,data_stage_1__484_,data_stage_1__483_,
  data_stage_1__482_,data_stage_1__481_,data_stage_1__480_,data_stage_1__479_,
  data_stage_1__478_,data_stage_1__477_,data_stage_1__476_,data_stage_1__475_,
  data_stage_1__474_,data_stage_1__473_,data_stage_1__472_,data_stage_1__471_,data_stage_1__470_,
  data_stage_1__469_,data_stage_1__468_,data_stage_1__467_,data_stage_1__466_,
  data_stage_1__465_,data_stage_1__464_,data_stage_1__463_,data_stage_1__462_,
  data_stage_1__461_,data_stage_1__460_,data_stage_1__459_,data_stage_1__458_,
  data_stage_1__457_,data_stage_1__456_,data_stage_1__455_,data_stage_1__454_,
  data_stage_1__453_,data_stage_1__452_,data_stage_1__451_,data_stage_1__450_,data_stage_1__449_,
  data_stage_1__448_,data_stage_1__447_,data_stage_1__446_,data_stage_1__445_,
  data_stage_1__444_,data_stage_1__443_,data_stage_1__442_,data_stage_1__441_,
  data_stage_1__440_,data_stage_1__439_,data_stage_1__438_,data_stage_1__437_,
  data_stage_1__436_,data_stage_1__435_,data_stage_1__434_,data_stage_1__433_,data_stage_1__432_,
  data_stage_1__431_,data_stage_1__430_,data_stage_1__429_,data_stage_1__428_,
  data_stage_1__427_,data_stage_1__426_,data_stage_1__425_,data_stage_1__424_,
  data_stage_1__423_,data_stage_1__422_,data_stage_1__421_,data_stage_1__420_,
  data_stage_1__419_,data_stage_1__418_,data_stage_1__417_,data_stage_1__416_,
  data_stage_1__415_,data_stage_1__414_,data_stage_1__413_,data_stage_1__412_,data_stage_1__411_,
  data_stage_1__410_,data_stage_1__409_,data_stage_1__408_,data_stage_1__407_,
  data_stage_1__406_,data_stage_1__405_,data_stage_1__404_,data_stage_1__403_,
  data_stage_1__402_,data_stage_1__401_,data_stage_1__400_,data_stage_1__399_,
  data_stage_1__398_,data_stage_1__397_,data_stage_1__396_,data_stage_1__395_,
  data_stage_1__394_,data_stage_1__393_,data_stage_1__392_,data_stage_1__391_,data_stage_1__390_,
  data_stage_1__389_,data_stage_1__388_,data_stage_1__387_,data_stage_1__386_,
  data_stage_1__385_,data_stage_1__384_,data_stage_1__383_,data_stage_1__382_,
  data_stage_1__381_,data_stage_1__380_,data_stage_1__379_,data_stage_1__378_,
  data_stage_1__377_,data_stage_1__376_,data_stage_1__375_,data_stage_1__374_,
  data_stage_1__373_,data_stage_1__372_,data_stage_1__371_,data_stage_1__370_,data_stage_1__369_,
  data_stage_1__368_,data_stage_1__367_,data_stage_1__366_,data_stage_1__365_,
  data_stage_1__364_,data_stage_1__363_,data_stage_1__362_,data_stage_1__361_,
  data_stage_1__360_,data_stage_1__359_,data_stage_1__358_,data_stage_1__357_,
  data_stage_1__356_,data_stage_1__355_,data_stage_1__354_,data_stage_1__353_,data_stage_1__352_,
  data_stage_1__351_,data_stage_1__350_,data_stage_1__349_,data_stage_1__348_,
  data_stage_1__347_,data_stage_1__346_,data_stage_1__345_,data_stage_1__344_,
  data_stage_1__343_,data_stage_1__342_,data_stage_1__341_,data_stage_1__340_,
  data_stage_1__339_,data_stage_1__338_,data_stage_1__337_,data_stage_1__336_,
  data_stage_1__335_,data_stage_1__334_,data_stage_1__333_,data_stage_1__332_,data_stage_1__331_,
  data_stage_1__330_,data_stage_1__329_,data_stage_1__328_,data_stage_1__327_,
  data_stage_1__326_,data_stage_1__325_,data_stage_1__324_,data_stage_1__323_,
  data_stage_1__322_,data_stage_1__321_,data_stage_1__320_,data_stage_1__319_,
  data_stage_1__318_,data_stage_1__317_,data_stage_1__316_,data_stage_1__315_,
  data_stage_1__314_,data_stage_1__313_,data_stage_1__312_,data_stage_1__311_,data_stage_1__310_,
  data_stage_1__309_,data_stage_1__308_,data_stage_1__307_,data_stage_1__306_,
  data_stage_1__305_,data_stage_1__304_,data_stage_1__303_,data_stage_1__302_,
  data_stage_1__301_,data_stage_1__300_,data_stage_1__299_,data_stage_1__298_,
  data_stage_1__297_,data_stage_1__296_,data_stage_1__295_,data_stage_1__294_,
  data_stage_1__293_,data_stage_1__292_,data_stage_1__291_,data_stage_1__290_,data_stage_1__289_,
  data_stage_1__288_,data_stage_1__287_,data_stage_1__286_,data_stage_1__285_,
  data_stage_1__284_,data_stage_1__283_,data_stage_1__282_,data_stage_1__281_,
  data_stage_1__280_,data_stage_1__279_,data_stage_1__278_,data_stage_1__277_,
  data_stage_1__276_,data_stage_1__275_,data_stage_1__274_,data_stage_1__273_,data_stage_1__272_,
  data_stage_1__271_,data_stage_1__270_,data_stage_1__269_,data_stage_1__268_,
  data_stage_1__267_,data_stage_1__266_,data_stage_1__265_,data_stage_1__264_,
  data_stage_1__263_,data_stage_1__262_,data_stage_1__261_,data_stage_1__260_,
  data_stage_1__259_,data_stage_1__258_,data_stage_1__257_,data_stage_1__256_,
  data_stage_1__255_,data_stage_1__254_,data_stage_1__253_,data_stage_1__252_,data_stage_1__251_,
  data_stage_1__250_,data_stage_1__249_,data_stage_1__248_,data_stage_1__247_,
  data_stage_1__246_,data_stage_1__245_,data_stage_1__244_,data_stage_1__243_,
  data_stage_1__242_,data_stage_1__241_,data_stage_1__240_,data_stage_1__239_,
  data_stage_1__238_,data_stage_1__237_,data_stage_1__236_,data_stage_1__235_,
  data_stage_1__234_,data_stage_1__233_,data_stage_1__232_,data_stage_1__231_,data_stage_1__230_,
  data_stage_1__229_,data_stage_1__228_,data_stage_1__227_,data_stage_1__226_,
  data_stage_1__225_,data_stage_1__224_,data_stage_1__223_,data_stage_1__222_,
  data_stage_1__221_,data_stage_1__220_,data_stage_1__219_,data_stage_1__218_,
  data_stage_1__217_,data_stage_1__216_,data_stage_1__215_,data_stage_1__214_,
  data_stage_1__213_,data_stage_1__212_,data_stage_1__211_,data_stage_1__210_,data_stage_1__209_,
  data_stage_1__208_,data_stage_1__207_,data_stage_1__206_,data_stage_1__205_,
  data_stage_1__204_,data_stage_1__203_,data_stage_1__202_,data_stage_1__201_,
  data_stage_1__200_,data_stage_1__199_,data_stage_1__198_,data_stage_1__197_,
  data_stage_1__196_,data_stage_1__195_,data_stage_1__194_,data_stage_1__193_,data_stage_1__192_,
  data_stage_1__191_,data_stage_1__190_,data_stage_1__189_,data_stage_1__188_,
  data_stage_1__187_,data_stage_1__186_,data_stage_1__185_,data_stage_1__184_,
  data_stage_1__183_,data_stage_1__182_,data_stage_1__181_,data_stage_1__180_,
  data_stage_1__179_,data_stage_1__178_,data_stage_1__177_,data_stage_1__176_,
  data_stage_1__175_,data_stage_1__174_,data_stage_1__173_,data_stage_1__172_,data_stage_1__171_,
  data_stage_1__170_,data_stage_1__169_,data_stage_1__168_,data_stage_1__167_,
  data_stage_1__166_,data_stage_1__165_,data_stage_1__164_,data_stage_1__163_,
  data_stage_1__162_,data_stage_1__161_,data_stage_1__160_,data_stage_1__159_,
  data_stage_1__158_,data_stage_1__157_,data_stage_1__156_,data_stage_1__155_,
  data_stage_1__154_,data_stage_1__153_,data_stage_1__152_,data_stage_1__151_,data_stage_1__150_,
  data_stage_1__149_,data_stage_1__148_,data_stage_1__147_,data_stage_1__146_,
  data_stage_1__145_,data_stage_1__144_,data_stage_1__143_,data_stage_1__142_,
  data_stage_1__141_,data_stage_1__140_,data_stage_1__139_,data_stage_1__138_,
  data_stage_1__137_,data_stage_1__136_,data_stage_1__135_,data_stage_1__134_,
  data_stage_1__133_,data_stage_1__132_,data_stage_1__131_,data_stage_1__130_,data_stage_1__129_,
  data_stage_1__128_,data_stage_1__127_,data_stage_1__126_,data_stage_1__125_,
  data_stage_1__124_,data_stage_1__123_,data_stage_1__122_,data_stage_1__121_,
  data_stage_1__120_,data_stage_1__119_,data_stage_1__118_,data_stage_1__117_,
  data_stage_1__116_,data_stage_1__115_,data_stage_1__114_,data_stage_1__113_,data_stage_1__112_,
  data_stage_1__111_,data_stage_1__110_,data_stage_1__109_,data_stage_1__108_,
  data_stage_1__107_,data_stage_1__106_,data_stage_1__105_,data_stage_1__104_,
  data_stage_1__103_,data_stage_1__102_,data_stage_1__101_,data_stage_1__100_,
  data_stage_1__99_,data_stage_1__98_,data_stage_1__97_,data_stage_1__96_,data_stage_1__95_,
  data_stage_1__94_,data_stage_1__93_,data_stage_1__92_,data_stage_1__91_,
  data_stage_1__90_,data_stage_1__89_,data_stage_1__88_,data_stage_1__87_,data_stage_1__86_,
  data_stage_1__85_,data_stage_1__84_,data_stage_1__83_,data_stage_1__82_,
  data_stage_1__81_,data_stage_1__80_,data_stage_1__79_,data_stage_1__78_,
  data_stage_1__77_,data_stage_1__76_,data_stage_1__75_,data_stage_1__74_,data_stage_1__73_,
  data_stage_1__72_,data_stage_1__71_,data_stage_1__70_,data_stage_1__69_,
  data_stage_1__68_,data_stage_1__67_,data_stage_1__66_,data_stage_1__65_,data_stage_1__64_,
  data_stage_1__63_,data_stage_1__62_,data_stage_1__61_,data_stage_1__60_,
  data_stage_1__59_,data_stage_1__58_,data_stage_1__57_,data_stage_1__56_,data_stage_1__55_,
  data_stage_1__54_,data_stage_1__53_,data_stage_1__52_,data_stage_1__51_,
  data_stage_1__50_,data_stage_1__49_,data_stage_1__48_,data_stage_1__47_,data_stage_1__46_,
  data_stage_1__45_,data_stage_1__44_,data_stage_1__43_,data_stage_1__42_,
  data_stage_1__41_,data_stage_1__40_,data_stage_1__39_,data_stage_1__38_,
  data_stage_1__37_,data_stage_1__36_,data_stage_1__35_,data_stage_1__34_,data_stage_1__33_,
  data_stage_1__32_,data_stage_1__31_,data_stage_1__30_,data_stage_1__29_,
  data_stage_1__28_,data_stage_1__27_,data_stage_1__26_,data_stage_1__25_,data_stage_1__24_,
  data_stage_1__23_,data_stage_1__22_,data_stage_1__21_,data_stage_1__20_,
  data_stage_1__19_,data_stage_1__18_,data_stage_1__17_,data_stage_1__16_,data_stage_1__15_,
  data_stage_1__14_,data_stage_1__13_,data_stage_1__12_,data_stage_1__11_,
  data_stage_1__10_,data_stage_1__9_,data_stage_1__8_,data_stage_1__7_,data_stage_1__6_,
  data_stage_1__5_,data_stage_1__4_,data_stage_1__3_,data_stage_1__2_,
  data_stage_1__1_,data_stage_1__0_,data_stage_2__511_,data_stage_2__510_,data_stage_2__509_,
  data_stage_2__508_,data_stage_2__507_,data_stage_2__506_,data_stage_2__505_,
  data_stage_2__504_,data_stage_2__503_,data_stage_2__502_,data_stage_2__501_,
  data_stage_2__500_,data_stage_2__499_,data_stage_2__498_,data_stage_2__497_,
  data_stage_2__496_,data_stage_2__495_,data_stage_2__494_,data_stage_2__493_,data_stage_2__492_,
  data_stage_2__491_,data_stage_2__490_,data_stage_2__489_,data_stage_2__488_,
  data_stage_2__487_,data_stage_2__486_,data_stage_2__485_,data_stage_2__484_,
  data_stage_2__483_,data_stage_2__482_,data_stage_2__481_,data_stage_2__480_,
  data_stage_2__479_,data_stage_2__478_,data_stage_2__477_,data_stage_2__476_,
  data_stage_2__475_,data_stage_2__474_,data_stage_2__473_,data_stage_2__472_,data_stage_2__471_,
  data_stage_2__470_,data_stage_2__469_,data_stage_2__468_,data_stage_2__467_,
  data_stage_2__466_,data_stage_2__465_,data_stage_2__464_,data_stage_2__463_,
  data_stage_2__462_,data_stage_2__461_,data_stage_2__460_,data_stage_2__459_,
  data_stage_2__458_,data_stage_2__457_,data_stage_2__456_,data_stage_2__455_,data_stage_2__454_,
  data_stage_2__453_,data_stage_2__452_,data_stage_2__451_,data_stage_2__450_,
  data_stage_2__449_,data_stage_2__448_,data_stage_2__447_,data_stage_2__446_,
  data_stage_2__445_,data_stage_2__444_,data_stage_2__443_,data_stage_2__442_,
  data_stage_2__441_,data_stage_2__440_,data_stage_2__439_,data_stage_2__438_,
  data_stage_2__437_,data_stage_2__436_,data_stage_2__435_,data_stage_2__434_,data_stage_2__433_,
  data_stage_2__432_,data_stage_2__431_,data_stage_2__430_,data_stage_2__429_,
  data_stage_2__428_,data_stage_2__427_,data_stage_2__426_,data_stage_2__425_,
  data_stage_2__424_,data_stage_2__423_,data_stage_2__422_,data_stage_2__421_,
  data_stage_2__420_,data_stage_2__419_,data_stage_2__418_,data_stage_2__417_,
  data_stage_2__416_,data_stage_2__415_,data_stage_2__414_,data_stage_2__413_,data_stage_2__412_,
  data_stage_2__411_,data_stage_2__410_,data_stage_2__409_,data_stage_2__408_,
  data_stage_2__407_,data_stage_2__406_,data_stage_2__405_,data_stage_2__404_,
  data_stage_2__403_,data_stage_2__402_,data_stage_2__401_,data_stage_2__400_,
  data_stage_2__399_,data_stage_2__398_,data_stage_2__397_,data_stage_2__396_,
  data_stage_2__395_,data_stage_2__394_,data_stage_2__393_,data_stage_2__392_,data_stage_2__391_,
  data_stage_2__390_,data_stage_2__389_,data_stage_2__388_,data_stage_2__387_,
  data_stage_2__386_,data_stage_2__385_,data_stage_2__384_,data_stage_2__383_,
  data_stage_2__382_,data_stage_2__381_,data_stage_2__380_,data_stage_2__379_,
  data_stage_2__378_,data_stage_2__377_,data_stage_2__376_,data_stage_2__375_,data_stage_2__374_,
  data_stage_2__373_,data_stage_2__372_,data_stage_2__371_,data_stage_2__370_,
  data_stage_2__369_,data_stage_2__368_,data_stage_2__367_,data_stage_2__366_,
  data_stage_2__365_,data_stage_2__364_,data_stage_2__363_,data_stage_2__362_,
  data_stage_2__361_,data_stage_2__360_,data_stage_2__359_,data_stage_2__358_,
  data_stage_2__357_,data_stage_2__356_,data_stage_2__355_,data_stage_2__354_,data_stage_2__353_,
  data_stage_2__352_,data_stage_2__351_,data_stage_2__350_,data_stage_2__349_,
  data_stage_2__348_,data_stage_2__347_,data_stage_2__346_,data_stage_2__345_,
  data_stage_2__344_,data_stage_2__343_,data_stage_2__342_,data_stage_2__341_,
  data_stage_2__340_,data_stage_2__339_,data_stage_2__338_,data_stage_2__337_,
  data_stage_2__336_,data_stage_2__335_,data_stage_2__334_,data_stage_2__333_,data_stage_2__332_,
  data_stage_2__331_,data_stage_2__330_,data_stage_2__329_,data_stage_2__328_,
  data_stage_2__327_,data_stage_2__326_,data_stage_2__325_,data_stage_2__324_,
  data_stage_2__323_,data_stage_2__322_,data_stage_2__321_,data_stage_2__320_,
  data_stage_2__319_,data_stage_2__318_,data_stage_2__317_,data_stage_2__316_,
  data_stage_2__315_,data_stage_2__314_,data_stage_2__313_,data_stage_2__312_,data_stage_2__311_,
  data_stage_2__310_,data_stage_2__309_,data_stage_2__308_,data_stage_2__307_,
  data_stage_2__306_,data_stage_2__305_,data_stage_2__304_,data_stage_2__303_,
  data_stage_2__302_,data_stage_2__301_,data_stage_2__300_,data_stage_2__299_,
  data_stage_2__298_,data_stage_2__297_,data_stage_2__296_,data_stage_2__295_,data_stage_2__294_,
  data_stage_2__293_,data_stage_2__292_,data_stage_2__291_,data_stage_2__290_,
  data_stage_2__289_,data_stage_2__288_,data_stage_2__287_,data_stage_2__286_,
  data_stage_2__285_,data_stage_2__284_,data_stage_2__283_,data_stage_2__282_,
  data_stage_2__281_,data_stage_2__280_,data_stage_2__279_,data_stage_2__278_,
  data_stage_2__277_,data_stage_2__276_,data_stage_2__275_,data_stage_2__274_,data_stage_2__273_,
  data_stage_2__272_,data_stage_2__271_,data_stage_2__270_,data_stage_2__269_,
  data_stage_2__268_,data_stage_2__267_,data_stage_2__266_,data_stage_2__265_,
  data_stage_2__264_,data_stage_2__263_,data_stage_2__262_,data_stage_2__261_,
  data_stage_2__260_,data_stage_2__259_,data_stage_2__258_,data_stage_2__257_,
  data_stage_2__256_,data_stage_2__255_,data_stage_2__254_,data_stage_2__253_,data_stage_2__252_,
  data_stage_2__251_,data_stage_2__250_,data_stage_2__249_,data_stage_2__248_,
  data_stage_2__247_,data_stage_2__246_,data_stage_2__245_,data_stage_2__244_,
  data_stage_2__243_,data_stage_2__242_,data_stage_2__241_,data_stage_2__240_,
  data_stage_2__239_,data_stage_2__238_,data_stage_2__237_,data_stage_2__236_,
  data_stage_2__235_,data_stage_2__234_,data_stage_2__233_,data_stage_2__232_,data_stage_2__231_,
  data_stage_2__230_,data_stage_2__229_,data_stage_2__228_,data_stage_2__227_,
  data_stage_2__226_,data_stage_2__225_,data_stage_2__224_,data_stage_2__223_,
  data_stage_2__222_,data_stage_2__221_,data_stage_2__220_,data_stage_2__219_,
  data_stage_2__218_,data_stage_2__217_,data_stage_2__216_,data_stage_2__215_,data_stage_2__214_,
  data_stage_2__213_,data_stage_2__212_,data_stage_2__211_,data_stage_2__210_,
  data_stage_2__209_,data_stage_2__208_,data_stage_2__207_,data_stage_2__206_,
  data_stage_2__205_,data_stage_2__204_,data_stage_2__203_,data_stage_2__202_,
  data_stage_2__201_,data_stage_2__200_,data_stage_2__199_,data_stage_2__198_,
  data_stage_2__197_,data_stage_2__196_,data_stage_2__195_,data_stage_2__194_,data_stage_2__193_,
  data_stage_2__192_,data_stage_2__191_,data_stage_2__190_,data_stage_2__189_,
  data_stage_2__188_,data_stage_2__187_,data_stage_2__186_,data_stage_2__185_,
  data_stage_2__184_,data_stage_2__183_,data_stage_2__182_,data_stage_2__181_,
  data_stage_2__180_,data_stage_2__179_,data_stage_2__178_,data_stage_2__177_,
  data_stage_2__176_,data_stage_2__175_,data_stage_2__174_,data_stage_2__173_,data_stage_2__172_,
  data_stage_2__171_,data_stage_2__170_,data_stage_2__169_,data_stage_2__168_,
  data_stage_2__167_,data_stage_2__166_,data_stage_2__165_,data_stage_2__164_,
  data_stage_2__163_,data_stage_2__162_,data_stage_2__161_,data_stage_2__160_,
  data_stage_2__159_,data_stage_2__158_,data_stage_2__157_,data_stage_2__156_,
  data_stage_2__155_,data_stage_2__154_,data_stage_2__153_,data_stage_2__152_,data_stage_2__151_,
  data_stage_2__150_,data_stage_2__149_,data_stage_2__148_,data_stage_2__147_,
  data_stage_2__146_,data_stage_2__145_,data_stage_2__144_,data_stage_2__143_,
  data_stage_2__142_,data_stage_2__141_,data_stage_2__140_,data_stage_2__139_,
  data_stage_2__138_,data_stage_2__137_,data_stage_2__136_,data_stage_2__135_,data_stage_2__134_,
  data_stage_2__133_,data_stage_2__132_,data_stage_2__131_,data_stage_2__130_,
  data_stage_2__129_,data_stage_2__128_,data_stage_2__127_,data_stage_2__126_,
  data_stage_2__125_,data_stage_2__124_,data_stage_2__123_,data_stage_2__122_,
  data_stage_2__121_,data_stage_2__120_,data_stage_2__119_,data_stage_2__118_,
  data_stage_2__117_,data_stage_2__116_,data_stage_2__115_,data_stage_2__114_,data_stage_2__113_,
  data_stage_2__112_,data_stage_2__111_,data_stage_2__110_,data_stage_2__109_,
  data_stage_2__108_,data_stage_2__107_,data_stage_2__106_,data_stage_2__105_,
  data_stage_2__104_,data_stage_2__103_,data_stage_2__102_,data_stage_2__101_,
  data_stage_2__100_,data_stage_2__99_,data_stage_2__98_,data_stage_2__97_,data_stage_2__96_,
  data_stage_2__95_,data_stage_2__94_,data_stage_2__93_,data_stage_2__92_,
  data_stage_2__91_,data_stage_2__90_,data_stage_2__89_,data_stage_2__88_,data_stage_2__87_,
  data_stage_2__86_,data_stage_2__85_,data_stage_2__84_,data_stage_2__83_,
  data_stage_2__82_,data_stage_2__81_,data_stage_2__80_,data_stage_2__79_,
  data_stage_2__78_,data_stage_2__77_,data_stage_2__76_,data_stage_2__75_,data_stage_2__74_,
  data_stage_2__73_,data_stage_2__72_,data_stage_2__71_,data_stage_2__70_,
  data_stage_2__69_,data_stage_2__68_,data_stage_2__67_,data_stage_2__66_,data_stage_2__65_,
  data_stage_2__64_,data_stage_2__63_,data_stage_2__62_,data_stage_2__61_,
  data_stage_2__60_,data_stage_2__59_,data_stage_2__58_,data_stage_2__57_,data_stage_2__56_,
  data_stage_2__55_,data_stage_2__54_,data_stage_2__53_,data_stage_2__52_,
  data_stage_2__51_,data_stage_2__50_,data_stage_2__49_,data_stage_2__48_,data_stage_2__47_,
  data_stage_2__46_,data_stage_2__45_,data_stage_2__44_,data_stage_2__43_,
  data_stage_2__42_,data_stage_2__41_,data_stage_2__40_,data_stage_2__39_,
  data_stage_2__38_,data_stage_2__37_,data_stage_2__36_,data_stage_2__35_,data_stage_2__34_,
  data_stage_2__33_,data_stage_2__32_,data_stage_2__31_,data_stage_2__30_,
  data_stage_2__29_,data_stage_2__28_,data_stage_2__27_,data_stage_2__26_,data_stage_2__25_,
  data_stage_2__24_,data_stage_2__23_,data_stage_2__22_,data_stage_2__21_,
  data_stage_2__20_,data_stage_2__19_,data_stage_2__18_,data_stage_2__17_,data_stage_2__16_,
  data_stage_2__15_,data_stage_2__14_,data_stage_2__13_,data_stage_2__12_,
  data_stage_2__11_,data_stage_2__10_,data_stage_2__9_,data_stage_2__8_,data_stage_2__7_,
  data_stage_2__6_,data_stage_2__5_,data_stage_2__4_,data_stage_2__3_,
  data_stage_2__2_,data_stage_2__1_,data_stage_2__0_;

  bsg_swap_width_p64
  mux_stage_0__mux_swap_0__swap_inst
  (
    .data_i(data_i[127:0]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__127_, data_stage_1__126_, data_stage_1__125_, data_stage_1__124_, data_stage_1__123_, data_stage_1__122_, data_stage_1__121_, data_stage_1__120_, data_stage_1__119_, data_stage_1__118_, data_stage_1__117_, data_stage_1__116_, data_stage_1__115_, data_stage_1__114_, data_stage_1__113_, data_stage_1__112_, data_stage_1__111_, data_stage_1__110_, data_stage_1__109_, data_stage_1__108_, data_stage_1__107_, data_stage_1__106_, data_stage_1__105_, data_stage_1__104_, data_stage_1__103_, data_stage_1__102_, data_stage_1__101_, data_stage_1__100_, data_stage_1__99_, data_stage_1__98_, data_stage_1__97_, data_stage_1__96_, data_stage_1__95_, data_stage_1__94_, data_stage_1__93_, data_stage_1__92_, data_stage_1__91_, data_stage_1__90_, data_stage_1__89_, data_stage_1__88_, data_stage_1__87_, data_stage_1__86_, data_stage_1__85_, data_stage_1__84_, data_stage_1__83_, data_stage_1__82_, data_stage_1__81_, data_stage_1__80_, data_stage_1__79_, data_stage_1__78_, data_stage_1__77_, data_stage_1__76_, data_stage_1__75_, data_stage_1__74_, data_stage_1__73_, data_stage_1__72_, data_stage_1__71_, data_stage_1__70_, data_stage_1__69_, data_stage_1__68_, data_stage_1__67_, data_stage_1__66_, data_stage_1__65_, data_stage_1__64_, data_stage_1__63_, data_stage_1__62_, data_stage_1__61_, data_stage_1__60_, data_stage_1__59_, data_stage_1__58_, data_stage_1__57_, data_stage_1__56_, data_stage_1__55_, data_stage_1__54_, data_stage_1__53_, data_stage_1__52_, data_stage_1__51_, data_stage_1__50_, data_stage_1__49_, data_stage_1__48_, data_stage_1__47_, data_stage_1__46_, data_stage_1__45_, data_stage_1__44_, data_stage_1__43_, data_stage_1__42_, data_stage_1__41_, data_stage_1__40_, data_stage_1__39_, data_stage_1__38_, data_stage_1__37_, data_stage_1__36_, data_stage_1__35_, data_stage_1__34_, data_stage_1__33_, data_stage_1__32_, data_stage_1__31_, data_stage_1__30_, data_stage_1__29_, data_stage_1__28_, data_stage_1__27_, data_stage_1__26_, data_stage_1__25_, data_stage_1__24_, data_stage_1__23_, data_stage_1__22_, data_stage_1__21_, data_stage_1__20_, data_stage_1__19_, data_stage_1__18_, data_stage_1__17_, data_stage_1__16_, data_stage_1__15_, data_stage_1__14_, data_stage_1__13_, data_stage_1__12_, data_stage_1__11_, data_stage_1__10_, data_stage_1__9_, data_stage_1__8_, data_stage_1__7_, data_stage_1__6_, data_stage_1__5_, data_stage_1__4_, data_stage_1__3_, data_stage_1__2_, data_stage_1__1_, data_stage_1__0_ })
  );


  bsg_swap_width_p64
  mux_stage_0__mux_swap_1__swap_inst
  (
    .data_i(data_i[255:128]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__255_, data_stage_1__254_, data_stage_1__253_, data_stage_1__252_, data_stage_1__251_, data_stage_1__250_, data_stage_1__249_, data_stage_1__248_, data_stage_1__247_, data_stage_1__246_, data_stage_1__245_, data_stage_1__244_, data_stage_1__243_, data_stage_1__242_, data_stage_1__241_, data_stage_1__240_, data_stage_1__239_, data_stage_1__238_, data_stage_1__237_, data_stage_1__236_, data_stage_1__235_, data_stage_1__234_, data_stage_1__233_, data_stage_1__232_, data_stage_1__231_, data_stage_1__230_, data_stage_1__229_, data_stage_1__228_, data_stage_1__227_, data_stage_1__226_, data_stage_1__225_, data_stage_1__224_, data_stage_1__223_, data_stage_1__222_, data_stage_1__221_, data_stage_1__220_, data_stage_1__219_, data_stage_1__218_, data_stage_1__217_, data_stage_1__216_, data_stage_1__215_, data_stage_1__214_, data_stage_1__213_, data_stage_1__212_, data_stage_1__211_, data_stage_1__210_, data_stage_1__209_, data_stage_1__208_, data_stage_1__207_, data_stage_1__206_, data_stage_1__205_, data_stage_1__204_, data_stage_1__203_, data_stage_1__202_, data_stage_1__201_, data_stage_1__200_, data_stage_1__199_, data_stage_1__198_, data_stage_1__197_, data_stage_1__196_, data_stage_1__195_, data_stage_1__194_, data_stage_1__193_, data_stage_1__192_, data_stage_1__191_, data_stage_1__190_, data_stage_1__189_, data_stage_1__188_, data_stage_1__187_, data_stage_1__186_, data_stage_1__185_, data_stage_1__184_, data_stage_1__183_, data_stage_1__182_, data_stage_1__181_, data_stage_1__180_, data_stage_1__179_, data_stage_1__178_, data_stage_1__177_, data_stage_1__176_, data_stage_1__175_, data_stage_1__174_, data_stage_1__173_, data_stage_1__172_, data_stage_1__171_, data_stage_1__170_, data_stage_1__169_, data_stage_1__168_, data_stage_1__167_, data_stage_1__166_, data_stage_1__165_, data_stage_1__164_, data_stage_1__163_, data_stage_1__162_, data_stage_1__161_, data_stage_1__160_, data_stage_1__159_, data_stage_1__158_, data_stage_1__157_, data_stage_1__156_, data_stage_1__155_, data_stage_1__154_, data_stage_1__153_, data_stage_1__152_, data_stage_1__151_, data_stage_1__150_, data_stage_1__149_, data_stage_1__148_, data_stage_1__147_, data_stage_1__146_, data_stage_1__145_, data_stage_1__144_, data_stage_1__143_, data_stage_1__142_, data_stage_1__141_, data_stage_1__140_, data_stage_1__139_, data_stage_1__138_, data_stage_1__137_, data_stage_1__136_, data_stage_1__135_, data_stage_1__134_, data_stage_1__133_, data_stage_1__132_, data_stage_1__131_, data_stage_1__130_, data_stage_1__129_, data_stage_1__128_ })
  );


  bsg_swap_width_p64
  mux_stage_0__mux_swap_2__swap_inst
  (
    .data_i(data_i[383:256]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__383_, data_stage_1__382_, data_stage_1__381_, data_stage_1__380_, data_stage_1__379_, data_stage_1__378_, data_stage_1__377_, data_stage_1__376_, data_stage_1__375_, data_stage_1__374_, data_stage_1__373_, data_stage_1__372_, data_stage_1__371_, data_stage_1__370_, data_stage_1__369_, data_stage_1__368_, data_stage_1__367_, data_stage_1__366_, data_stage_1__365_, data_stage_1__364_, data_stage_1__363_, data_stage_1__362_, data_stage_1__361_, data_stage_1__360_, data_stage_1__359_, data_stage_1__358_, data_stage_1__357_, data_stage_1__356_, data_stage_1__355_, data_stage_1__354_, data_stage_1__353_, data_stage_1__352_, data_stage_1__351_, data_stage_1__350_, data_stage_1__349_, data_stage_1__348_, data_stage_1__347_, data_stage_1__346_, data_stage_1__345_, data_stage_1__344_, data_stage_1__343_, data_stage_1__342_, data_stage_1__341_, data_stage_1__340_, data_stage_1__339_, data_stage_1__338_, data_stage_1__337_, data_stage_1__336_, data_stage_1__335_, data_stage_1__334_, data_stage_1__333_, data_stage_1__332_, data_stage_1__331_, data_stage_1__330_, data_stage_1__329_, data_stage_1__328_, data_stage_1__327_, data_stage_1__326_, data_stage_1__325_, data_stage_1__324_, data_stage_1__323_, data_stage_1__322_, data_stage_1__321_, data_stage_1__320_, data_stage_1__319_, data_stage_1__318_, data_stage_1__317_, data_stage_1__316_, data_stage_1__315_, data_stage_1__314_, data_stage_1__313_, data_stage_1__312_, data_stage_1__311_, data_stage_1__310_, data_stage_1__309_, data_stage_1__308_, data_stage_1__307_, data_stage_1__306_, data_stage_1__305_, data_stage_1__304_, data_stage_1__303_, data_stage_1__302_, data_stage_1__301_, data_stage_1__300_, data_stage_1__299_, data_stage_1__298_, data_stage_1__297_, data_stage_1__296_, data_stage_1__295_, data_stage_1__294_, data_stage_1__293_, data_stage_1__292_, data_stage_1__291_, data_stage_1__290_, data_stage_1__289_, data_stage_1__288_, data_stage_1__287_, data_stage_1__286_, data_stage_1__285_, data_stage_1__284_, data_stage_1__283_, data_stage_1__282_, data_stage_1__281_, data_stage_1__280_, data_stage_1__279_, data_stage_1__278_, data_stage_1__277_, data_stage_1__276_, data_stage_1__275_, data_stage_1__274_, data_stage_1__273_, data_stage_1__272_, data_stage_1__271_, data_stage_1__270_, data_stage_1__269_, data_stage_1__268_, data_stage_1__267_, data_stage_1__266_, data_stage_1__265_, data_stage_1__264_, data_stage_1__263_, data_stage_1__262_, data_stage_1__261_, data_stage_1__260_, data_stage_1__259_, data_stage_1__258_, data_stage_1__257_, data_stage_1__256_ })
  );


  bsg_swap_width_p64
  mux_stage_0__mux_swap_3__swap_inst
  (
    .data_i(data_i[511:384]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__511_, data_stage_1__510_, data_stage_1__509_, data_stage_1__508_, data_stage_1__507_, data_stage_1__506_, data_stage_1__505_, data_stage_1__504_, data_stage_1__503_, data_stage_1__502_, data_stage_1__501_, data_stage_1__500_, data_stage_1__499_, data_stage_1__498_, data_stage_1__497_, data_stage_1__496_, data_stage_1__495_, data_stage_1__494_, data_stage_1__493_, data_stage_1__492_, data_stage_1__491_, data_stage_1__490_, data_stage_1__489_, data_stage_1__488_, data_stage_1__487_, data_stage_1__486_, data_stage_1__485_, data_stage_1__484_, data_stage_1__483_, data_stage_1__482_, data_stage_1__481_, data_stage_1__480_, data_stage_1__479_, data_stage_1__478_, data_stage_1__477_, data_stage_1__476_, data_stage_1__475_, data_stage_1__474_, data_stage_1__473_, data_stage_1__472_, data_stage_1__471_, data_stage_1__470_, data_stage_1__469_, data_stage_1__468_, data_stage_1__467_, data_stage_1__466_, data_stage_1__465_, data_stage_1__464_, data_stage_1__463_, data_stage_1__462_, data_stage_1__461_, data_stage_1__460_, data_stage_1__459_, data_stage_1__458_, data_stage_1__457_, data_stage_1__456_, data_stage_1__455_, data_stage_1__454_, data_stage_1__453_, data_stage_1__452_, data_stage_1__451_, data_stage_1__450_, data_stage_1__449_, data_stage_1__448_, data_stage_1__447_, data_stage_1__446_, data_stage_1__445_, data_stage_1__444_, data_stage_1__443_, data_stage_1__442_, data_stage_1__441_, data_stage_1__440_, data_stage_1__439_, data_stage_1__438_, data_stage_1__437_, data_stage_1__436_, data_stage_1__435_, data_stage_1__434_, data_stage_1__433_, data_stage_1__432_, data_stage_1__431_, data_stage_1__430_, data_stage_1__429_, data_stage_1__428_, data_stage_1__427_, data_stage_1__426_, data_stage_1__425_, data_stage_1__424_, data_stage_1__423_, data_stage_1__422_, data_stage_1__421_, data_stage_1__420_, data_stage_1__419_, data_stage_1__418_, data_stage_1__417_, data_stage_1__416_, data_stage_1__415_, data_stage_1__414_, data_stage_1__413_, data_stage_1__412_, data_stage_1__411_, data_stage_1__410_, data_stage_1__409_, data_stage_1__408_, data_stage_1__407_, data_stage_1__406_, data_stage_1__405_, data_stage_1__404_, data_stage_1__403_, data_stage_1__402_, data_stage_1__401_, data_stage_1__400_, data_stage_1__399_, data_stage_1__398_, data_stage_1__397_, data_stage_1__396_, data_stage_1__395_, data_stage_1__394_, data_stage_1__393_, data_stage_1__392_, data_stage_1__391_, data_stage_1__390_, data_stage_1__389_, data_stage_1__388_, data_stage_1__387_, data_stage_1__386_, data_stage_1__385_, data_stage_1__384_ })
  );


  bsg_swap_width_p128
  mux_stage_1__mux_swap_0__swap_inst
  (
    .data_i({ data_stage_1__255_, data_stage_1__254_, data_stage_1__253_, data_stage_1__252_, data_stage_1__251_, data_stage_1__250_, data_stage_1__249_, data_stage_1__248_, data_stage_1__247_, data_stage_1__246_, data_stage_1__245_, data_stage_1__244_, data_stage_1__243_, data_stage_1__242_, data_stage_1__241_, data_stage_1__240_, data_stage_1__239_, data_stage_1__238_, data_stage_1__237_, data_stage_1__236_, data_stage_1__235_, data_stage_1__234_, data_stage_1__233_, data_stage_1__232_, data_stage_1__231_, data_stage_1__230_, data_stage_1__229_, data_stage_1__228_, data_stage_1__227_, data_stage_1__226_, data_stage_1__225_, data_stage_1__224_, data_stage_1__223_, data_stage_1__222_, data_stage_1__221_, data_stage_1__220_, data_stage_1__219_, data_stage_1__218_, data_stage_1__217_, data_stage_1__216_, data_stage_1__215_, data_stage_1__214_, data_stage_1__213_, data_stage_1__212_, data_stage_1__211_, data_stage_1__210_, data_stage_1__209_, data_stage_1__208_, data_stage_1__207_, data_stage_1__206_, data_stage_1__205_, data_stage_1__204_, data_stage_1__203_, data_stage_1__202_, data_stage_1__201_, data_stage_1__200_, data_stage_1__199_, data_stage_1__198_, data_stage_1__197_, data_stage_1__196_, data_stage_1__195_, data_stage_1__194_, data_stage_1__193_, data_stage_1__192_, data_stage_1__191_, data_stage_1__190_, data_stage_1__189_, data_stage_1__188_, data_stage_1__187_, data_stage_1__186_, data_stage_1__185_, data_stage_1__184_, data_stage_1__183_, data_stage_1__182_, data_stage_1__181_, data_stage_1__180_, data_stage_1__179_, data_stage_1__178_, data_stage_1__177_, data_stage_1__176_, data_stage_1__175_, data_stage_1__174_, data_stage_1__173_, data_stage_1__172_, data_stage_1__171_, data_stage_1__170_, data_stage_1__169_, data_stage_1__168_, data_stage_1__167_, data_stage_1__166_, data_stage_1__165_, data_stage_1__164_, data_stage_1__163_, data_stage_1__162_, data_stage_1__161_, data_stage_1__160_, data_stage_1__159_, data_stage_1__158_, data_stage_1__157_, data_stage_1__156_, data_stage_1__155_, data_stage_1__154_, data_stage_1__153_, data_stage_1__152_, data_stage_1__151_, data_stage_1__150_, data_stage_1__149_, data_stage_1__148_, data_stage_1__147_, data_stage_1__146_, data_stage_1__145_, data_stage_1__144_, data_stage_1__143_, data_stage_1__142_, data_stage_1__141_, data_stage_1__140_, data_stage_1__139_, data_stage_1__138_, data_stage_1__137_, data_stage_1__136_, data_stage_1__135_, data_stage_1__134_, data_stage_1__133_, data_stage_1__132_, data_stage_1__131_, data_stage_1__130_, data_stage_1__129_, data_stage_1__128_, data_stage_1__127_, data_stage_1__126_, data_stage_1__125_, data_stage_1__124_, data_stage_1__123_, data_stage_1__122_, data_stage_1__121_, data_stage_1__120_, data_stage_1__119_, data_stage_1__118_, data_stage_1__117_, data_stage_1__116_, data_stage_1__115_, data_stage_1__114_, data_stage_1__113_, data_stage_1__112_, data_stage_1__111_, data_stage_1__110_, data_stage_1__109_, data_stage_1__108_, data_stage_1__107_, data_stage_1__106_, data_stage_1__105_, data_stage_1__104_, data_stage_1__103_, data_stage_1__102_, data_stage_1__101_, data_stage_1__100_, data_stage_1__99_, data_stage_1__98_, data_stage_1__97_, data_stage_1__96_, data_stage_1__95_, data_stage_1__94_, data_stage_1__93_, data_stage_1__92_, data_stage_1__91_, data_stage_1__90_, data_stage_1__89_, data_stage_1__88_, data_stage_1__87_, data_stage_1__86_, data_stage_1__85_, data_stage_1__84_, data_stage_1__83_, data_stage_1__82_, data_stage_1__81_, data_stage_1__80_, data_stage_1__79_, data_stage_1__78_, data_stage_1__77_, data_stage_1__76_, data_stage_1__75_, data_stage_1__74_, data_stage_1__73_, data_stage_1__72_, data_stage_1__71_, data_stage_1__70_, data_stage_1__69_, data_stage_1__68_, data_stage_1__67_, data_stage_1__66_, data_stage_1__65_, data_stage_1__64_, data_stage_1__63_, data_stage_1__62_, data_stage_1__61_, data_stage_1__60_, data_stage_1__59_, data_stage_1__58_, data_stage_1__57_, data_stage_1__56_, data_stage_1__55_, data_stage_1__54_, data_stage_1__53_, data_stage_1__52_, data_stage_1__51_, data_stage_1__50_, data_stage_1__49_, data_stage_1__48_, data_stage_1__47_, data_stage_1__46_, data_stage_1__45_, data_stage_1__44_, data_stage_1__43_, data_stage_1__42_, data_stage_1__41_, data_stage_1__40_, data_stage_1__39_, data_stage_1__38_, data_stage_1__37_, data_stage_1__36_, data_stage_1__35_, data_stage_1__34_, data_stage_1__33_, data_stage_1__32_, data_stage_1__31_, data_stage_1__30_, data_stage_1__29_, data_stage_1__28_, data_stage_1__27_, data_stage_1__26_, data_stage_1__25_, data_stage_1__24_, data_stage_1__23_, data_stage_1__22_, data_stage_1__21_, data_stage_1__20_, data_stage_1__19_, data_stage_1__18_, data_stage_1__17_, data_stage_1__16_, data_stage_1__15_, data_stage_1__14_, data_stage_1__13_, data_stage_1__12_, data_stage_1__11_, data_stage_1__10_, data_stage_1__9_, data_stage_1__8_, data_stage_1__7_, data_stage_1__6_, data_stage_1__5_, data_stage_1__4_, data_stage_1__3_, data_stage_1__2_, data_stage_1__1_, data_stage_1__0_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__255_, data_stage_2__254_, data_stage_2__253_, data_stage_2__252_, data_stage_2__251_, data_stage_2__250_, data_stage_2__249_, data_stage_2__248_, data_stage_2__247_, data_stage_2__246_, data_stage_2__245_, data_stage_2__244_, data_stage_2__243_, data_stage_2__242_, data_stage_2__241_, data_stage_2__240_, data_stage_2__239_, data_stage_2__238_, data_stage_2__237_, data_stage_2__236_, data_stage_2__235_, data_stage_2__234_, data_stage_2__233_, data_stage_2__232_, data_stage_2__231_, data_stage_2__230_, data_stage_2__229_, data_stage_2__228_, data_stage_2__227_, data_stage_2__226_, data_stage_2__225_, data_stage_2__224_, data_stage_2__223_, data_stage_2__222_, data_stage_2__221_, data_stage_2__220_, data_stage_2__219_, data_stage_2__218_, data_stage_2__217_, data_stage_2__216_, data_stage_2__215_, data_stage_2__214_, data_stage_2__213_, data_stage_2__212_, data_stage_2__211_, data_stage_2__210_, data_stage_2__209_, data_stage_2__208_, data_stage_2__207_, data_stage_2__206_, data_stage_2__205_, data_stage_2__204_, data_stage_2__203_, data_stage_2__202_, data_stage_2__201_, data_stage_2__200_, data_stage_2__199_, data_stage_2__198_, data_stage_2__197_, data_stage_2__196_, data_stage_2__195_, data_stage_2__194_, data_stage_2__193_, data_stage_2__192_, data_stage_2__191_, data_stage_2__190_, data_stage_2__189_, data_stage_2__188_, data_stage_2__187_, data_stage_2__186_, data_stage_2__185_, data_stage_2__184_, data_stage_2__183_, data_stage_2__182_, data_stage_2__181_, data_stage_2__180_, data_stage_2__179_, data_stage_2__178_, data_stage_2__177_, data_stage_2__176_, data_stage_2__175_, data_stage_2__174_, data_stage_2__173_, data_stage_2__172_, data_stage_2__171_, data_stage_2__170_, data_stage_2__169_, data_stage_2__168_, data_stage_2__167_, data_stage_2__166_, data_stage_2__165_, data_stage_2__164_, data_stage_2__163_, data_stage_2__162_, data_stage_2__161_, data_stage_2__160_, data_stage_2__159_, data_stage_2__158_, data_stage_2__157_, data_stage_2__156_, data_stage_2__155_, data_stage_2__154_, data_stage_2__153_, data_stage_2__152_, data_stage_2__151_, data_stage_2__150_, data_stage_2__149_, data_stage_2__148_, data_stage_2__147_, data_stage_2__146_, data_stage_2__145_, data_stage_2__144_, data_stage_2__143_, data_stage_2__142_, data_stage_2__141_, data_stage_2__140_, data_stage_2__139_, data_stage_2__138_, data_stage_2__137_, data_stage_2__136_, data_stage_2__135_, data_stage_2__134_, data_stage_2__133_, data_stage_2__132_, data_stage_2__131_, data_stage_2__130_, data_stage_2__129_, data_stage_2__128_, data_stage_2__127_, data_stage_2__126_, data_stage_2__125_, data_stage_2__124_, data_stage_2__123_, data_stage_2__122_, data_stage_2__121_, data_stage_2__120_, data_stage_2__119_, data_stage_2__118_, data_stage_2__117_, data_stage_2__116_, data_stage_2__115_, data_stage_2__114_, data_stage_2__113_, data_stage_2__112_, data_stage_2__111_, data_stage_2__110_, data_stage_2__109_, data_stage_2__108_, data_stage_2__107_, data_stage_2__106_, data_stage_2__105_, data_stage_2__104_, data_stage_2__103_, data_stage_2__102_, data_stage_2__101_, data_stage_2__100_, data_stage_2__99_, data_stage_2__98_, data_stage_2__97_, data_stage_2__96_, data_stage_2__95_, data_stage_2__94_, data_stage_2__93_, data_stage_2__92_, data_stage_2__91_, data_stage_2__90_, data_stage_2__89_, data_stage_2__88_, data_stage_2__87_, data_stage_2__86_, data_stage_2__85_, data_stage_2__84_, data_stage_2__83_, data_stage_2__82_, data_stage_2__81_, data_stage_2__80_, data_stage_2__79_, data_stage_2__78_, data_stage_2__77_, data_stage_2__76_, data_stage_2__75_, data_stage_2__74_, data_stage_2__73_, data_stage_2__72_, data_stage_2__71_, data_stage_2__70_, data_stage_2__69_, data_stage_2__68_, data_stage_2__67_, data_stage_2__66_, data_stage_2__65_, data_stage_2__64_, data_stage_2__63_, data_stage_2__62_, data_stage_2__61_, data_stage_2__60_, data_stage_2__59_, data_stage_2__58_, data_stage_2__57_, data_stage_2__56_, data_stage_2__55_, data_stage_2__54_, data_stage_2__53_, data_stage_2__52_, data_stage_2__51_, data_stage_2__50_, data_stage_2__49_, data_stage_2__48_, data_stage_2__47_, data_stage_2__46_, data_stage_2__45_, data_stage_2__44_, data_stage_2__43_, data_stage_2__42_, data_stage_2__41_, data_stage_2__40_, data_stage_2__39_, data_stage_2__38_, data_stage_2__37_, data_stage_2__36_, data_stage_2__35_, data_stage_2__34_, data_stage_2__33_, data_stage_2__32_, data_stage_2__31_, data_stage_2__30_, data_stage_2__29_, data_stage_2__28_, data_stage_2__27_, data_stage_2__26_, data_stage_2__25_, data_stage_2__24_, data_stage_2__23_, data_stage_2__22_, data_stage_2__21_, data_stage_2__20_, data_stage_2__19_, data_stage_2__18_, data_stage_2__17_, data_stage_2__16_, data_stage_2__15_, data_stage_2__14_, data_stage_2__13_, data_stage_2__12_, data_stage_2__11_, data_stage_2__10_, data_stage_2__9_, data_stage_2__8_, data_stage_2__7_, data_stage_2__6_, data_stage_2__5_, data_stage_2__4_, data_stage_2__3_, data_stage_2__2_, data_stage_2__1_, data_stage_2__0_ })
  );


  bsg_swap_width_p128
  mux_stage_1__mux_swap_1__swap_inst
  (
    .data_i({ data_stage_1__511_, data_stage_1__510_, data_stage_1__509_, data_stage_1__508_, data_stage_1__507_, data_stage_1__506_, data_stage_1__505_, data_stage_1__504_, data_stage_1__503_, data_stage_1__502_, data_stage_1__501_, data_stage_1__500_, data_stage_1__499_, data_stage_1__498_, data_stage_1__497_, data_stage_1__496_, data_stage_1__495_, data_stage_1__494_, data_stage_1__493_, data_stage_1__492_, data_stage_1__491_, data_stage_1__490_, data_stage_1__489_, data_stage_1__488_, data_stage_1__487_, data_stage_1__486_, data_stage_1__485_, data_stage_1__484_, data_stage_1__483_, data_stage_1__482_, data_stage_1__481_, data_stage_1__480_, data_stage_1__479_, data_stage_1__478_, data_stage_1__477_, data_stage_1__476_, data_stage_1__475_, data_stage_1__474_, data_stage_1__473_, data_stage_1__472_, data_stage_1__471_, data_stage_1__470_, data_stage_1__469_, data_stage_1__468_, data_stage_1__467_, data_stage_1__466_, data_stage_1__465_, data_stage_1__464_, data_stage_1__463_, data_stage_1__462_, data_stage_1__461_, data_stage_1__460_, data_stage_1__459_, data_stage_1__458_, data_stage_1__457_, data_stage_1__456_, data_stage_1__455_, data_stage_1__454_, data_stage_1__453_, data_stage_1__452_, data_stage_1__451_, data_stage_1__450_, data_stage_1__449_, data_stage_1__448_, data_stage_1__447_, data_stage_1__446_, data_stage_1__445_, data_stage_1__444_, data_stage_1__443_, data_stage_1__442_, data_stage_1__441_, data_stage_1__440_, data_stage_1__439_, data_stage_1__438_, data_stage_1__437_, data_stage_1__436_, data_stage_1__435_, data_stage_1__434_, data_stage_1__433_, data_stage_1__432_, data_stage_1__431_, data_stage_1__430_, data_stage_1__429_, data_stage_1__428_, data_stage_1__427_, data_stage_1__426_, data_stage_1__425_, data_stage_1__424_, data_stage_1__423_, data_stage_1__422_, data_stage_1__421_, data_stage_1__420_, data_stage_1__419_, data_stage_1__418_, data_stage_1__417_, data_stage_1__416_, data_stage_1__415_, data_stage_1__414_, data_stage_1__413_, data_stage_1__412_, data_stage_1__411_, data_stage_1__410_, data_stage_1__409_, data_stage_1__408_, data_stage_1__407_, data_stage_1__406_, data_stage_1__405_, data_stage_1__404_, data_stage_1__403_, data_stage_1__402_, data_stage_1__401_, data_stage_1__400_, data_stage_1__399_, data_stage_1__398_, data_stage_1__397_, data_stage_1__396_, data_stage_1__395_, data_stage_1__394_, data_stage_1__393_, data_stage_1__392_, data_stage_1__391_, data_stage_1__390_, data_stage_1__389_, data_stage_1__388_, data_stage_1__387_, data_stage_1__386_, data_stage_1__385_, data_stage_1__384_, data_stage_1__383_, data_stage_1__382_, data_stage_1__381_, data_stage_1__380_, data_stage_1__379_, data_stage_1__378_, data_stage_1__377_, data_stage_1__376_, data_stage_1__375_, data_stage_1__374_, data_stage_1__373_, data_stage_1__372_, data_stage_1__371_, data_stage_1__370_, data_stage_1__369_, data_stage_1__368_, data_stage_1__367_, data_stage_1__366_, data_stage_1__365_, data_stage_1__364_, data_stage_1__363_, data_stage_1__362_, data_stage_1__361_, data_stage_1__360_, data_stage_1__359_, data_stage_1__358_, data_stage_1__357_, data_stage_1__356_, data_stage_1__355_, data_stage_1__354_, data_stage_1__353_, data_stage_1__352_, data_stage_1__351_, data_stage_1__350_, data_stage_1__349_, data_stage_1__348_, data_stage_1__347_, data_stage_1__346_, data_stage_1__345_, data_stage_1__344_, data_stage_1__343_, data_stage_1__342_, data_stage_1__341_, data_stage_1__340_, data_stage_1__339_, data_stage_1__338_, data_stage_1__337_, data_stage_1__336_, data_stage_1__335_, data_stage_1__334_, data_stage_1__333_, data_stage_1__332_, data_stage_1__331_, data_stage_1__330_, data_stage_1__329_, data_stage_1__328_, data_stage_1__327_, data_stage_1__326_, data_stage_1__325_, data_stage_1__324_, data_stage_1__323_, data_stage_1__322_, data_stage_1__321_, data_stage_1__320_, data_stage_1__319_, data_stage_1__318_, data_stage_1__317_, data_stage_1__316_, data_stage_1__315_, data_stage_1__314_, data_stage_1__313_, data_stage_1__312_, data_stage_1__311_, data_stage_1__310_, data_stage_1__309_, data_stage_1__308_, data_stage_1__307_, data_stage_1__306_, data_stage_1__305_, data_stage_1__304_, data_stage_1__303_, data_stage_1__302_, data_stage_1__301_, data_stage_1__300_, data_stage_1__299_, data_stage_1__298_, data_stage_1__297_, data_stage_1__296_, data_stage_1__295_, data_stage_1__294_, data_stage_1__293_, data_stage_1__292_, data_stage_1__291_, data_stage_1__290_, data_stage_1__289_, data_stage_1__288_, data_stage_1__287_, data_stage_1__286_, data_stage_1__285_, data_stage_1__284_, data_stage_1__283_, data_stage_1__282_, data_stage_1__281_, data_stage_1__280_, data_stage_1__279_, data_stage_1__278_, data_stage_1__277_, data_stage_1__276_, data_stage_1__275_, data_stage_1__274_, data_stage_1__273_, data_stage_1__272_, data_stage_1__271_, data_stage_1__270_, data_stage_1__269_, data_stage_1__268_, data_stage_1__267_, data_stage_1__266_, data_stage_1__265_, data_stage_1__264_, data_stage_1__263_, data_stage_1__262_, data_stage_1__261_, data_stage_1__260_, data_stage_1__259_, data_stage_1__258_, data_stage_1__257_, data_stage_1__256_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__511_, data_stage_2__510_, data_stage_2__509_, data_stage_2__508_, data_stage_2__507_, data_stage_2__506_, data_stage_2__505_, data_stage_2__504_, data_stage_2__503_, data_stage_2__502_, data_stage_2__501_, data_stage_2__500_, data_stage_2__499_, data_stage_2__498_, data_stage_2__497_, data_stage_2__496_, data_stage_2__495_, data_stage_2__494_, data_stage_2__493_, data_stage_2__492_, data_stage_2__491_, data_stage_2__490_, data_stage_2__489_, data_stage_2__488_, data_stage_2__487_, data_stage_2__486_, data_stage_2__485_, data_stage_2__484_, data_stage_2__483_, data_stage_2__482_, data_stage_2__481_, data_stage_2__480_, data_stage_2__479_, data_stage_2__478_, data_stage_2__477_, data_stage_2__476_, data_stage_2__475_, data_stage_2__474_, data_stage_2__473_, data_stage_2__472_, data_stage_2__471_, data_stage_2__470_, data_stage_2__469_, data_stage_2__468_, data_stage_2__467_, data_stage_2__466_, data_stage_2__465_, data_stage_2__464_, data_stage_2__463_, data_stage_2__462_, data_stage_2__461_, data_stage_2__460_, data_stage_2__459_, data_stage_2__458_, data_stage_2__457_, data_stage_2__456_, data_stage_2__455_, data_stage_2__454_, data_stage_2__453_, data_stage_2__452_, data_stage_2__451_, data_stage_2__450_, data_stage_2__449_, data_stage_2__448_, data_stage_2__447_, data_stage_2__446_, data_stage_2__445_, data_stage_2__444_, data_stage_2__443_, data_stage_2__442_, data_stage_2__441_, data_stage_2__440_, data_stage_2__439_, data_stage_2__438_, data_stage_2__437_, data_stage_2__436_, data_stage_2__435_, data_stage_2__434_, data_stage_2__433_, data_stage_2__432_, data_stage_2__431_, data_stage_2__430_, data_stage_2__429_, data_stage_2__428_, data_stage_2__427_, data_stage_2__426_, data_stage_2__425_, data_stage_2__424_, data_stage_2__423_, data_stage_2__422_, data_stage_2__421_, data_stage_2__420_, data_stage_2__419_, data_stage_2__418_, data_stage_2__417_, data_stage_2__416_, data_stage_2__415_, data_stage_2__414_, data_stage_2__413_, data_stage_2__412_, data_stage_2__411_, data_stage_2__410_, data_stage_2__409_, data_stage_2__408_, data_stage_2__407_, data_stage_2__406_, data_stage_2__405_, data_stage_2__404_, data_stage_2__403_, data_stage_2__402_, data_stage_2__401_, data_stage_2__400_, data_stage_2__399_, data_stage_2__398_, data_stage_2__397_, data_stage_2__396_, data_stage_2__395_, data_stage_2__394_, data_stage_2__393_, data_stage_2__392_, data_stage_2__391_, data_stage_2__390_, data_stage_2__389_, data_stage_2__388_, data_stage_2__387_, data_stage_2__386_, data_stage_2__385_, data_stage_2__384_, data_stage_2__383_, data_stage_2__382_, data_stage_2__381_, data_stage_2__380_, data_stage_2__379_, data_stage_2__378_, data_stage_2__377_, data_stage_2__376_, data_stage_2__375_, data_stage_2__374_, data_stage_2__373_, data_stage_2__372_, data_stage_2__371_, data_stage_2__370_, data_stage_2__369_, data_stage_2__368_, data_stage_2__367_, data_stage_2__366_, data_stage_2__365_, data_stage_2__364_, data_stage_2__363_, data_stage_2__362_, data_stage_2__361_, data_stage_2__360_, data_stage_2__359_, data_stage_2__358_, data_stage_2__357_, data_stage_2__356_, data_stage_2__355_, data_stage_2__354_, data_stage_2__353_, data_stage_2__352_, data_stage_2__351_, data_stage_2__350_, data_stage_2__349_, data_stage_2__348_, data_stage_2__347_, data_stage_2__346_, data_stage_2__345_, data_stage_2__344_, data_stage_2__343_, data_stage_2__342_, data_stage_2__341_, data_stage_2__340_, data_stage_2__339_, data_stage_2__338_, data_stage_2__337_, data_stage_2__336_, data_stage_2__335_, data_stage_2__334_, data_stage_2__333_, data_stage_2__332_, data_stage_2__331_, data_stage_2__330_, data_stage_2__329_, data_stage_2__328_, data_stage_2__327_, data_stage_2__326_, data_stage_2__325_, data_stage_2__324_, data_stage_2__323_, data_stage_2__322_, data_stage_2__321_, data_stage_2__320_, data_stage_2__319_, data_stage_2__318_, data_stage_2__317_, data_stage_2__316_, data_stage_2__315_, data_stage_2__314_, data_stage_2__313_, data_stage_2__312_, data_stage_2__311_, data_stage_2__310_, data_stage_2__309_, data_stage_2__308_, data_stage_2__307_, data_stage_2__306_, data_stage_2__305_, data_stage_2__304_, data_stage_2__303_, data_stage_2__302_, data_stage_2__301_, data_stage_2__300_, data_stage_2__299_, data_stage_2__298_, data_stage_2__297_, data_stage_2__296_, data_stage_2__295_, data_stage_2__294_, data_stage_2__293_, data_stage_2__292_, data_stage_2__291_, data_stage_2__290_, data_stage_2__289_, data_stage_2__288_, data_stage_2__287_, data_stage_2__286_, data_stage_2__285_, data_stage_2__284_, data_stage_2__283_, data_stage_2__282_, data_stage_2__281_, data_stage_2__280_, data_stage_2__279_, data_stage_2__278_, data_stage_2__277_, data_stage_2__276_, data_stage_2__275_, data_stage_2__274_, data_stage_2__273_, data_stage_2__272_, data_stage_2__271_, data_stage_2__270_, data_stage_2__269_, data_stage_2__268_, data_stage_2__267_, data_stage_2__266_, data_stage_2__265_, data_stage_2__264_, data_stage_2__263_, data_stage_2__262_, data_stage_2__261_, data_stage_2__260_, data_stage_2__259_, data_stage_2__258_, data_stage_2__257_, data_stage_2__256_ })
  );


  bsg_swap_width_p256
  mux_stage_2__mux_swap_0__swap_inst
  (
    .data_i({ data_stage_2__511_, data_stage_2__510_, data_stage_2__509_, data_stage_2__508_, data_stage_2__507_, data_stage_2__506_, data_stage_2__505_, data_stage_2__504_, data_stage_2__503_, data_stage_2__502_, data_stage_2__501_, data_stage_2__500_, data_stage_2__499_, data_stage_2__498_, data_stage_2__497_, data_stage_2__496_, data_stage_2__495_, data_stage_2__494_, data_stage_2__493_, data_stage_2__492_, data_stage_2__491_, data_stage_2__490_, data_stage_2__489_, data_stage_2__488_, data_stage_2__487_, data_stage_2__486_, data_stage_2__485_, data_stage_2__484_, data_stage_2__483_, data_stage_2__482_, data_stage_2__481_, data_stage_2__480_, data_stage_2__479_, data_stage_2__478_, data_stage_2__477_, data_stage_2__476_, data_stage_2__475_, data_stage_2__474_, data_stage_2__473_, data_stage_2__472_, data_stage_2__471_, data_stage_2__470_, data_stage_2__469_, data_stage_2__468_, data_stage_2__467_, data_stage_2__466_, data_stage_2__465_, data_stage_2__464_, data_stage_2__463_, data_stage_2__462_, data_stage_2__461_, data_stage_2__460_, data_stage_2__459_, data_stage_2__458_, data_stage_2__457_, data_stage_2__456_, data_stage_2__455_, data_stage_2__454_, data_stage_2__453_, data_stage_2__452_, data_stage_2__451_, data_stage_2__450_, data_stage_2__449_, data_stage_2__448_, data_stage_2__447_, data_stage_2__446_, data_stage_2__445_, data_stage_2__444_, data_stage_2__443_, data_stage_2__442_, data_stage_2__441_, data_stage_2__440_, data_stage_2__439_, data_stage_2__438_, data_stage_2__437_, data_stage_2__436_, data_stage_2__435_, data_stage_2__434_, data_stage_2__433_, data_stage_2__432_, data_stage_2__431_, data_stage_2__430_, data_stage_2__429_, data_stage_2__428_, data_stage_2__427_, data_stage_2__426_, data_stage_2__425_, data_stage_2__424_, data_stage_2__423_, data_stage_2__422_, data_stage_2__421_, data_stage_2__420_, data_stage_2__419_, data_stage_2__418_, data_stage_2__417_, data_stage_2__416_, data_stage_2__415_, data_stage_2__414_, data_stage_2__413_, data_stage_2__412_, data_stage_2__411_, data_stage_2__410_, data_stage_2__409_, data_stage_2__408_, data_stage_2__407_, data_stage_2__406_, data_stage_2__405_, data_stage_2__404_, data_stage_2__403_, data_stage_2__402_, data_stage_2__401_, data_stage_2__400_, data_stage_2__399_, data_stage_2__398_, data_stage_2__397_, data_stage_2__396_, data_stage_2__395_, data_stage_2__394_, data_stage_2__393_, data_stage_2__392_, data_stage_2__391_, data_stage_2__390_, data_stage_2__389_, data_stage_2__388_, data_stage_2__387_, data_stage_2__386_, data_stage_2__385_, data_stage_2__384_, data_stage_2__383_, data_stage_2__382_, data_stage_2__381_, data_stage_2__380_, data_stage_2__379_, data_stage_2__378_, data_stage_2__377_, data_stage_2__376_, data_stage_2__375_, data_stage_2__374_, data_stage_2__373_, data_stage_2__372_, data_stage_2__371_, data_stage_2__370_, data_stage_2__369_, data_stage_2__368_, data_stage_2__367_, data_stage_2__366_, data_stage_2__365_, data_stage_2__364_, data_stage_2__363_, data_stage_2__362_, data_stage_2__361_, data_stage_2__360_, data_stage_2__359_, data_stage_2__358_, data_stage_2__357_, data_stage_2__356_, data_stage_2__355_, data_stage_2__354_, data_stage_2__353_, data_stage_2__352_, data_stage_2__351_, data_stage_2__350_, data_stage_2__349_, data_stage_2__348_, data_stage_2__347_, data_stage_2__346_, data_stage_2__345_, data_stage_2__344_, data_stage_2__343_, data_stage_2__342_, data_stage_2__341_, data_stage_2__340_, data_stage_2__339_, data_stage_2__338_, data_stage_2__337_, data_stage_2__336_, data_stage_2__335_, data_stage_2__334_, data_stage_2__333_, data_stage_2__332_, data_stage_2__331_, data_stage_2__330_, data_stage_2__329_, data_stage_2__328_, data_stage_2__327_, data_stage_2__326_, data_stage_2__325_, data_stage_2__324_, data_stage_2__323_, data_stage_2__322_, data_stage_2__321_, data_stage_2__320_, data_stage_2__319_, data_stage_2__318_, data_stage_2__317_, data_stage_2__316_, data_stage_2__315_, data_stage_2__314_, data_stage_2__313_, data_stage_2__312_, data_stage_2__311_, data_stage_2__310_, data_stage_2__309_, data_stage_2__308_, data_stage_2__307_, data_stage_2__306_, data_stage_2__305_, data_stage_2__304_, data_stage_2__303_, data_stage_2__302_, data_stage_2__301_, data_stage_2__300_, data_stage_2__299_, data_stage_2__298_, data_stage_2__297_, data_stage_2__296_, data_stage_2__295_, data_stage_2__294_, data_stage_2__293_, data_stage_2__292_, data_stage_2__291_, data_stage_2__290_, data_stage_2__289_, data_stage_2__288_, data_stage_2__287_, data_stage_2__286_, data_stage_2__285_, data_stage_2__284_, data_stage_2__283_, data_stage_2__282_, data_stage_2__281_, data_stage_2__280_, data_stage_2__279_, data_stage_2__278_, data_stage_2__277_, data_stage_2__276_, data_stage_2__275_, data_stage_2__274_, data_stage_2__273_, data_stage_2__272_, data_stage_2__271_, data_stage_2__270_, data_stage_2__269_, data_stage_2__268_, data_stage_2__267_, data_stage_2__266_, data_stage_2__265_, data_stage_2__264_, data_stage_2__263_, data_stage_2__262_, data_stage_2__261_, data_stage_2__260_, data_stage_2__259_, data_stage_2__258_, data_stage_2__257_, data_stage_2__256_, data_stage_2__255_, data_stage_2__254_, data_stage_2__253_, data_stage_2__252_, data_stage_2__251_, data_stage_2__250_, data_stage_2__249_, data_stage_2__248_, data_stage_2__247_, data_stage_2__246_, data_stage_2__245_, data_stage_2__244_, data_stage_2__243_, data_stage_2__242_, data_stage_2__241_, data_stage_2__240_, data_stage_2__239_, data_stage_2__238_, data_stage_2__237_, data_stage_2__236_, data_stage_2__235_, data_stage_2__234_, data_stage_2__233_, data_stage_2__232_, data_stage_2__231_, data_stage_2__230_, data_stage_2__229_, data_stage_2__228_, data_stage_2__227_, data_stage_2__226_, data_stage_2__225_, data_stage_2__224_, data_stage_2__223_, data_stage_2__222_, data_stage_2__221_, data_stage_2__220_, data_stage_2__219_, data_stage_2__218_, data_stage_2__217_, data_stage_2__216_, data_stage_2__215_, data_stage_2__214_, data_stage_2__213_, data_stage_2__212_, data_stage_2__211_, data_stage_2__210_, data_stage_2__209_, data_stage_2__208_, data_stage_2__207_, data_stage_2__206_, data_stage_2__205_, data_stage_2__204_, data_stage_2__203_, data_stage_2__202_, data_stage_2__201_, data_stage_2__200_, data_stage_2__199_, data_stage_2__198_, data_stage_2__197_, data_stage_2__196_, data_stage_2__195_, data_stage_2__194_, data_stage_2__193_, data_stage_2__192_, data_stage_2__191_, data_stage_2__190_, data_stage_2__189_, data_stage_2__188_, data_stage_2__187_, data_stage_2__186_, data_stage_2__185_, data_stage_2__184_, data_stage_2__183_, data_stage_2__182_, data_stage_2__181_, data_stage_2__180_, data_stage_2__179_, data_stage_2__178_, data_stage_2__177_, data_stage_2__176_, data_stage_2__175_, data_stage_2__174_, data_stage_2__173_, data_stage_2__172_, data_stage_2__171_, data_stage_2__170_, data_stage_2__169_, data_stage_2__168_, data_stage_2__167_, data_stage_2__166_, data_stage_2__165_, data_stage_2__164_, data_stage_2__163_, data_stage_2__162_, data_stage_2__161_, data_stage_2__160_, data_stage_2__159_, data_stage_2__158_, data_stage_2__157_, data_stage_2__156_, data_stage_2__155_, data_stage_2__154_, data_stage_2__153_, data_stage_2__152_, data_stage_2__151_, data_stage_2__150_, data_stage_2__149_, data_stage_2__148_, data_stage_2__147_, data_stage_2__146_, data_stage_2__145_, data_stage_2__144_, data_stage_2__143_, data_stage_2__142_, data_stage_2__141_, data_stage_2__140_, data_stage_2__139_, data_stage_2__138_, data_stage_2__137_, data_stage_2__136_, data_stage_2__135_, data_stage_2__134_, data_stage_2__133_, data_stage_2__132_, data_stage_2__131_, data_stage_2__130_, data_stage_2__129_, data_stage_2__128_, data_stage_2__127_, data_stage_2__126_, data_stage_2__125_, data_stage_2__124_, data_stage_2__123_, data_stage_2__122_, data_stage_2__121_, data_stage_2__120_, data_stage_2__119_, data_stage_2__118_, data_stage_2__117_, data_stage_2__116_, data_stage_2__115_, data_stage_2__114_, data_stage_2__113_, data_stage_2__112_, data_stage_2__111_, data_stage_2__110_, data_stage_2__109_, data_stage_2__108_, data_stage_2__107_, data_stage_2__106_, data_stage_2__105_, data_stage_2__104_, data_stage_2__103_, data_stage_2__102_, data_stage_2__101_, data_stage_2__100_, data_stage_2__99_, data_stage_2__98_, data_stage_2__97_, data_stage_2__96_, data_stage_2__95_, data_stage_2__94_, data_stage_2__93_, data_stage_2__92_, data_stage_2__91_, data_stage_2__90_, data_stage_2__89_, data_stage_2__88_, data_stage_2__87_, data_stage_2__86_, data_stage_2__85_, data_stage_2__84_, data_stage_2__83_, data_stage_2__82_, data_stage_2__81_, data_stage_2__80_, data_stage_2__79_, data_stage_2__78_, data_stage_2__77_, data_stage_2__76_, data_stage_2__75_, data_stage_2__74_, data_stage_2__73_, data_stage_2__72_, data_stage_2__71_, data_stage_2__70_, data_stage_2__69_, data_stage_2__68_, data_stage_2__67_, data_stage_2__66_, data_stage_2__65_, data_stage_2__64_, data_stage_2__63_, data_stage_2__62_, data_stage_2__61_, data_stage_2__60_, data_stage_2__59_, data_stage_2__58_, data_stage_2__57_, data_stage_2__56_, data_stage_2__55_, data_stage_2__54_, data_stage_2__53_, data_stage_2__52_, data_stage_2__51_, data_stage_2__50_, data_stage_2__49_, data_stage_2__48_, data_stage_2__47_, data_stage_2__46_, data_stage_2__45_, data_stage_2__44_, data_stage_2__43_, data_stage_2__42_, data_stage_2__41_, data_stage_2__40_, data_stage_2__39_, data_stage_2__38_, data_stage_2__37_, data_stage_2__36_, data_stage_2__35_, data_stage_2__34_, data_stage_2__33_, data_stage_2__32_, data_stage_2__31_, data_stage_2__30_, data_stage_2__29_, data_stage_2__28_, data_stage_2__27_, data_stage_2__26_, data_stage_2__25_, data_stage_2__24_, data_stage_2__23_, data_stage_2__22_, data_stage_2__21_, data_stage_2__20_, data_stage_2__19_, data_stage_2__18_, data_stage_2__17_, data_stage_2__16_, data_stage_2__15_, data_stage_2__14_, data_stage_2__13_, data_stage_2__12_, data_stage_2__11_, data_stage_2__10_, data_stage_2__9_, data_stage_2__8_, data_stage_2__7_, data_stage_2__6_, data_stage_2__5_, data_stage_2__4_, data_stage_2__3_, data_stage_2__2_, data_stage_2__1_, data_stage_2__0_ }),
    .swap_i(sel_i[2]),
    .data_o(data_o)
  );


endmodule



module bsg_decode_num_out_p8
(
  i,
  o
);

  input [2:0] i;
  output [7:0] o;
  wire [7:0] o;
  assign o = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << i;

endmodule



module bsg_lru_pseudo_tree_decode_ways_p8
(
  way_id_i,
  data_o,
  mask_o
);

  input [2:0] way_id_i;
  output [6:0] data_o;
  output [6:0] mask_o;
  wire [6:0] data_o,mask_o;
  wire N0,N1,N2;
  assign mask_o[0] = 1'b1;
  assign data_o[0] = 1'b1 & N0;
  assign N0 = ~way_id_i[2];
  assign mask_o[1] = 1'b1 & N0;
  assign data_o[1] = mask_o[1] & N1;
  assign N1 = ~way_id_i[1];
  assign mask_o[2] = 1'b1 & way_id_i[2];
  assign data_o[2] = mask_o[2] & N1;
  assign mask_o[3] = mask_o[1] & N1;
  assign data_o[3] = mask_o[3] & N2;
  assign N2 = ~way_id_i[0];
  assign mask_o[4] = mask_o[1] & way_id_i[1];
  assign data_o[4] = mask_o[4] & N2;
  assign mask_o[5] = mask_o[2] & N1;
  assign data_o[5] = mask_o[5] & N2;
  assign mask_o[6] = mask_o[2] & way_id_i[1];
  assign data_o[6] = mask_o[6] & N2;

endmodule



module bp_fe_icache_02
(
  clk_i,
  reset_i,
  freeze_i,
  id_i,
  cfg_w_v_i,
  cfg_addr_i,
  cfg_data_i,
  pc_gen_icache_vaddr_i,
  pc_gen_icache_vaddr_v_i,
  pc_gen_icache_vaddr_ready_o,
  icache_pc_gen_data_o,
  icache_pc_gen_data_v_o,
  icache_pc_gen_data_ready_i,
  itlb_icache_data_resp_i,
  itlb_icache_data_resp_v_i,
  itlb_icache_data_resp_ready_o,
  itlb_icache_miss_i,
  uncached_i,
  cache_miss_o,
  instr_access_fault_o,
  poison_tl_i,
  lce_req_o,
  lce_req_v_o,
  lce_req_ready_i,
  lce_resp_o,
  lce_resp_v_o,
  lce_resp_ready_i,
  lce_data_resp_o,
  lce_data_resp_v_o,
  lce_data_resp_ready_i,
  lce_cmd_i,
  lce_cmd_v_i,
  lce_cmd_ready_o,
  lce_data_cmd_i,
  lce_data_cmd_v_i,
  lce_data_cmd_ready_o,
  lce_data_cmd_o,
  lce_data_cmd_v_o,
  lce_data_cmd_ready_i
);

  input [0:0] id_i;
  input [15:0] cfg_addr_i;
  input [31:0] cfg_data_i;
  input [38:0] pc_gen_icache_vaddr_i;
  output [70:0] icache_pc_gen_data_o;
  input [26:0] itlb_icache_data_resp_i;
  output [113:0] lce_req_o;
  output [42:0] lce_resp_o;
  output [553:0] lce_data_resp_o;
  input [52:0] lce_cmd_i;
  input [517:0] lce_data_cmd_i;
  output [517:0] lce_data_cmd_o;
  input clk_i;
  input reset_i;
  input freeze_i;
  input cfg_w_v_i;
  input pc_gen_icache_vaddr_v_i;
  input icache_pc_gen_data_ready_i;
  input itlb_icache_data_resp_v_i;
  input itlb_icache_miss_i;
  input uncached_i;
  input poison_tl_i;
  input lce_req_ready_i;
  input lce_resp_ready_i;
  input lce_data_resp_ready_i;
  input lce_cmd_v_i;
  input lce_data_cmd_v_i;
  input lce_data_cmd_ready_i;
  output pc_gen_icache_vaddr_ready_o;
  output icache_pc_gen_data_v_o;
  output itlb_icache_data_resp_ready_o;
  output cache_miss_o;
  output instr_access_fault_o;
  output lce_req_v_o;
  output lce_resp_v_o;
  output lce_data_resp_v_o;
  output lce_cmd_ready_o;
  output lce_data_cmd_ready_o;
  output lce_data_cmd_v_o;
  wire [113:0] lce_req_o;
  wire [42:0] lce_resp_o;
  wire [553:0] lce_data_resp_o;
  wire [517:0] lce_data_cmd_o;
  wire pc_gen_icache_vaddr_ready_o,icache_pc_gen_data_v_o,cache_miss_o,
  instr_access_fault_o,lce_req_v_o,lce_resp_v_o,lce_data_resp_v_o,lce_cmd_ready_o,
  lce_data_cmd_ready_o,lce_data_cmd_v_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,
  N17,N18,N19,N20,N21,N22,tl_we,N23,N24,N25,N26,n_0_net_,tag_mem_w_li,
  tag_mem_v_li,n_1_net_,data_mem_w_li,n_2_net_,n_3_net_,n_4_net_,n_5_net_,n_6_net_,n_7_net_,
  n_8_net_,tv_we,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,
  N43,N44,N45,N46,hit,miss_tv,uncached_req,n_9_net_,stat_mem_w_li,stat_mem_v_li,
  n_10_net__7_,n_10_net__6_,n_10_net__5_,n_10_net__4_,n_10_net__3_,n_10_net__2_,
  n_10_net__1_,n_10_net__0_,invalid_exist,N47,lce_data_mem_pkt_v_lo,
  lce_data_mem_pkt_yumi_li,tag_mem_pkt_v_lo,tag_mem_pkt_yumi_li,stat_mem_pkt_v_lo,stat_mem_pkt_yumi_li,
  lce_mode_lo,N48,N49,N50,n_11_net__2_,n_11_net__1_,n_11_net__0_,N51,N52,
  lce_data_mem_v,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,
  N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,
  N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,
  N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,
  N125,N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,
  N141,N142;
  wire [231:0] tag_mem_data_li,tag_mem_w_mask_li,tag_mem_data_lo;
  wire [5:0] tag_mem_addr_li,stat_mem_addr_li;
  wire [511:0] data_mem_data_li,data_mem_data_lo,lce_data_mem_data_li;
  wire [71:0] data_mem_addr_li;
  wire [7:0] data_mem_v_li,hit_v,lce_tag_mem_way_one_hot;
  wire [2:0] hit_index,lru_encode,way_invalid_index,lru_way_li;
  wire [6:0] stat_mem_data_li,stat_mem_mask_li,stat_mem_data_lo,lru_decode_data_lo,
  lru_decode_mask_lo;
  wire [522:0] lce_data_mem_pkt;
  wire [39:0] tag_mem_pkt;
  wire [9:0] stat_mem_pkt;
  wire [63:0] ld_data_way_picked,final_data;
  reg [38:0] vaddr_tl_r,addr_tv_r;
  reg itlb_icache_data_resp_ready_o,v_tv_r,uncached_tv_r,uncached_load_data_v_r;
  reg [511:0] ld_data_tv_r;
  reg [70:0] icache_pc_gen_data_o;
  reg [215:0] tag_tv_r;
  reg [15:0] state_tv_r;
  reg [2:0] lce_data_mem_pkt_way_r;
  reg [63:0] uncached_load_data_r;

  bsg_mem_1rw_sync_mask_write_bit_width_p232_els_p64
  tag_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(tag_mem_data_li),
    .addr_i(tag_mem_addr_li),
    .v_i(n_0_net_),
    .w_mask_i(tag_mem_w_mask_li),
    .w_i(tag_mem_w_li),
    .data_o(tag_mem_data_lo)
  );


  bsg_mem_1rw_sync_mask_write_byte_els_p512_data_width_p64
  data_mems_0__data_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(n_1_net_),
    .w_i(data_mem_w_li),
    .addr_i(data_mem_addr_li[8:0]),
    .data_i(data_mem_data_li[63:0]),
    .write_mask_i({ 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 }),
    .data_o(data_mem_data_lo[63:0])
  );


  bsg_mem_1rw_sync_mask_write_byte_els_p512_data_width_p64
  data_mems_1__data_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(n_2_net_),
    .w_i(data_mem_w_li),
    .addr_i(data_mem_addr_li[17:9]),
    .data_i(data_mem_data_li[127:64]),
    .write_mask_i({ 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 }),
    .data_o(data_mem_data_lo[127:64])
  );


  bsg_mem_1rw_sync_mask_write_byte_els_p512_data_width_p64
  data_mems_2__data_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(n_3_net_),
    .w_i(data_mem_w_li),
    .addr_i(data_mem_addr_li[26:18]),
    .data_i(data_mem_data_li[191:128]),
    .write_mask_i({ 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 }),
    .data_o(data_mem_data_lo[191:128])
  );


  bsg_mem_1rw_sync_mask_write_byte_els_p512_data_width_p64
  data_mems_3__data_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(n_4_net_),
    .w_i(data_mem_w_li),
    .addr_i(data_mem_addr_li[35:27]),
    .data_i(data_mem_data_li[255:192]),
    .write_mask_i({ 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 }),
    .data_o(data_mem_data_lo[255:192])
  );


  bsg_mem_1rw_sync_mask_write_byte_els_p512_data_width_p64
  data_mems_4__data_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(n_5_net_),
    .w_i(data_mem_w_li),
    .addr_i(data_mem_addr_li[44:36]),
    .data_i(data_mem_data_li[319:256]),
    .write_mask_i({ 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 }),
    .data_o(data_mem_data_lo[319:256])
  );


  bsg_mem_1rw_sync_mask_write_byte_els_p512_data_width_p64
  data_mems_5__data_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(n_6_net_),
    .w_i(data_mem_w_li),
    .addr_i(data_mem_addr_li[53:45]),
    .data_i(data_mem_data_li[383:320]),
    .write_mask_i({ 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 }),
    .data_o(data_mem_data_lo[383:320])
  );


  bsg_mem_1rw_sync_mask_write_byte_els_p512_data_width_p64
  data_mems_6__data_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(n_7_net_),
    .w_i(data_mem_w_li),
    .addr_i(data_mem_addr_li[62:54]),
    .data_i(data_mem_data_li[447:384]),
    .write_mask_i({ 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 }),
    .data_o(data_mem_data_lo[447:384])
  );


  bsg_mem_1rw_sync_mask_write_byte_els_p512_data_width_p64
  data_mems_7__data_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(n_8_net_),
    .w_i(data_mem_w_li),
    .addr_i(data_mem_addr_li[71:63]),
    .data_i(data_mem_data_li[511:448]),
    .write_mask_i({ 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 }),
    .data_o(data_mem_data_lo[511:448])
  );

  assign N39 = tag_tv_r[26:0] == addr_tv_r[38:12];
  assign N40 = tag_tv_r[53:27] == addr_tv_r[38:12];
  assign N41 = tag_tv_r[80:54] == addr_tv_r[38:12];
  assign N42 = tag_tv_r[107:81] == addr_tv_r[38:12];
  assign N43 = tag_tv_r[134:108] == addr_tv_r[38:12];
  assign N44 = tag_tv_r[161:135] == addr_tv_r[38:12];
  assign N45 = tag_tv_r[188:162] == addr_tv_r[38:12];
  assign N46 = tag_tv_r[215:189] == addr_tv_r[38:12];

  bsg_priority_encode_width_p8_lo_to_hi_p1
  pe_load_hit
  (
    .i(hit_v),
    .addr_o(hit_index),
    .v_o(hit)
  );


  bsg_mem_1rw_sync_mask_write_bit_width_p7_els_p64
  stat_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(stat_mem_data_li),
    .addr_i(stat_mem_addr_li),
    .v_i(n_9_net_),
    .w_mask_i(stat_mem_mask_li),
    .w_i(stat_mem_w_li),
    .data_o(stat_mem_data_lo)
  );


  bsg_lru_pseudo_tree_encode_ways_p8
  lru_encoder
  (
    .lru_i(stat_mem_data_lo),
    .way_id_o(lru_encode)
  );


  bsg_priority_encode_width_p8_lo_to_hi_p1
  pe_invalid
  (
    .i({ n_10_net__7_, n_10_net__6_, n_10_net__5_, n_10_net__4_, n_10_net__3_, n_10_net__2_, n_10_net__1_, n_10_net__0_ }),
    .addr_o(way_invalid_index),
    .v_o(invalid_exist)
  );


  bp_fe_lce_02
  lce
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .freeze_i(freeze_i),
    .cfg_w_v_i(cfg_w_v_i),
    .cfg_addr_i(cfg_addr_i),
    .cfg_data_i(cfg_data_i),
    .id_i(id_i[0]),
    .ready_o(pc_gen_icache_vaddr_ready_o),
    .cache_miss_o(cache_miss_o),
    .miss_i(miss_tv),
    .miss_addr_i(addr_tv_r),
    .uncached_req_i(uncached_req),
    .data_mem_data_i(lce_data_mem_data_li),
    .data_mem_pkt_o(lce_data_mem_pkt),
    .data_mem_pkt_v_o(lce_data_mem_pkt_v_lo),
    .data_mem_pkt_yumi_i(lce_data_mem_pkt_yumi_li),
    .tag_mem_pkt_o(tag_mem_pkt),
    .tag_mem_pkt_v_o(tag_mem_pkt_v_lo),
    .tag_mem_pkt_yumi_i(tag_mem_pkt_yumi_li),
    .stat_mem_pkt_v_o(stat_mem_pkt_v_lo),
    .stat_mem_pkt_o(stat_mem_pkt),
    .lru_way_i(lru_way_li),
    .stat_mem_pkt_yumi_i(stat_mem_pkt_yumi_li),
    .lce_req_o(lce_req_o),
    .lce_req_v_o(lce_req_v_o),
    .lce_req_ready_i(lce_req_ready_i),
    .lce_resp_o(lce_resp_o),
    .lce_resp_v_o(lce_resp_v_o),
    .lce_resp_ready_i(lce_resp_ready_i),
    .lce_data_resp_o(lce_data_resp_o),
    .lce_data_resp_v_o(lce_data_resp_v_o),
    .lce_data_resp_ready_i(lce_data_resp_ready_i),
    .lce_cmd_i(lce_cmd_i),
    .lce_cmd_v_i(lce_cmd_v_i),
    .lce_cmd_ready_o(lce_cmd_ready_o),
    .lce_data_cmd_i(lce_data_cmd_i),
    .lce_data_cmd_v_i(lce_data_cmd_v_i),
    .lce_data_cmd_ready_o(lce_data_cmd_ready_o),
    .lce_data_cmd_o(lce_data_cmd_o),
    .lce_data_cmd_v_o(lce_data_cmd_v_o),
    .lce_data_cmd_ready_i(lce_data_cmd_ready_i),
    .lce_mode_o(lce_mode_lo)
  );


  bsg_mux_width_p64_els_p8
  data_set_select_mux
  (
    .data_i(ld_data_tv_r),
    .sel_i({ n_11_net__2_, n_11_net__1_, n_11_net__0_ }),
    .data_o(ld_data_way_picked)
  );


  bsg_mux_width_p64_els_p2
  final_data_mux
  (
    .data_i({ uncached_load_data_r, ld_data_way_picked }),
    .sel_i(uncached_load_data_v_r),
    .data_o(final_data)
  );


  bsg_mux_butterfly_width_p64_els_p8
  write_mux_butterfly
  (
    .data_i(lce_data_mem_pkt[513:2]),
    .sel_i(lce_data_mem_pkt[516:514]),
    .data_o(data_mem_data_li)
  );


  bsg_decode_num_out_p8
  lce_tag_mem_way_decode
  (
    .i(tag_mem_pkt[33:31]),
    .o(lce_tag_mem_way_one_hot)
  );

  assign N68 = N66 & N67;
  assign N69 = tag_mem_pkt[1] | N67;
  assign N71 = N66 | tag_mem_pkt[0];
  assign N73 = tag_mem_pkt[1] & tag_mem_pkt[0];

  bsg_lru_pseudo_tree_decode_ways_p8
  lru_decode
  (
    .way_id_i(hit_index),
    .data_o(lru_decode_data_lo),
    .mask_o(lru_decode_mask_lo)
  );


  bsg_mux_butterfly_width_p64_els_p8
  read_mux_butterfly
  (
    .data_i(data_mem_data_lo),
    .sel_i(lce_data_mem_pkt_way_r),
    .data_o(lce_data_mem_data_li)
  );

  assign N91 = lce_data_mem_pkt[0] | lce_data_mem_pkt[1];
  assign N92 = ~N91;
  assign N93 = state_tv_r[14] | state_tv_r[15];
  assign N94 = state_tv_r[12] | state_tv_r[13];
  assign N95 = state_tv_r[10] | state_tv_r[11];
  assign N96 = state_tv_r[8] | state_tv_r[9];
  assign N97 = state_tv_r[6] | state_tv_r[7];
  assign N98 = state_tv_r[4] | state_tv_r[5];
  assign N99 = state_tv_r[2] | state_tv_r[3];
  assign N100 = state_tv_r[0] | state_tv_r[1];
  assign N101 = state_tv_r[14] | state_tv_r[15];
  assign N102 = state_tv_r[12] | state_tv_r[13];
  assign N103 = state_tv_r[10] | state_tv_r[11];
  assign N104 = state_tv_r[8] | state_tv_r[9];
  assign N105 = state_tv_r[6] | state_tv_r[7];
  assign N106 = state_tv_r[4] | state_tv_r[5];
  assign N107 = state_tv_r[2] | state_tv_r[3];
  assign N108 = state_tv_r[0] | state_tv_r[1];
  assign N109 = ~lce_mode_lo;
  assign N110 = ~stat_mem_pkt[0];
  assign N111 = ~lce_data_mem_pkt[1];
  assign N112 = lce_data_mem_pkt[0] | N111;
  assign N113 = ~lce_data_mem_pkt[0];
  assign N114 = N113 | lce_data_mem_pkt[1];
  assign N115 = ~N114;
  assign N116 = lce_data_mem_pkt[0] | N111;
  assign N117 = ~N116;
  assign N118 = lce_data_mem_pkt[0] | N111;
  assign N119 = ~N118;
  assign N25 = (N0)? 1'b0 : 
               (N1)? tl_we : 1'b0;
  assign N0 = N24;
  assign N1 = N23;
  assign N26 = (N0)? 1'b0 : 
               (N1)? tl_we : 1'b0;
  assign N29 = (N2)? 1'b0 : 
               (N3)? tv_we : 1'b0;
  assign N2 = N28;
  assign N3 = N27;
  assign { N38, N37, N36, N35, N34, N33, N32, N31, N30 } = (N2)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                           (N3)? { tv_we, tv_we, tv_we, tv_we, tv_we, tv_we, tv_we, tv_we, tv_we } : 1'b0;
  assign lru_way_li = (N4)? way_invalid_index : 
                      (N5)? lru_encode : 1'b0;
  assign N4 = invalid_exist;
  assign N5 = N47;
  assign instr_access_fault_o = (N6)? N135 : 
                                (N7)? 1'b0 : 1'b0;
  assign N6 = N109;
  assign N7 = lce_mode_lo;
  assign N50 = (N8)? uncached_load_data_v_r : 
               (N9)? N49 : 1'b0;
  assign N8 = uncached_tv_r;
  assign N9 = N135;
  assign icache_pc_gen_data_v_o = (N10)? N50 : 
                                  (N11)? 1'b0 : 1'b0;
  assign N10 = v_tv_r;
  assign N11 = N48;
  assign icache_pc_gen_data_o[70:39] = (N12)? final_data[63:32] : 
                                       (N13)? final_data[31:0] : 1'b0;
  assign N12 = N52;
  assign N13 = N51;
  assign data_mem_v_li = (N14)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                         (N15)? { lce_data_mem_v, lce_data_mem_v, lce_data_mem_v, lce_data_mem_v, lce_data_mem_v, lce_data_mem_v, lce_data_mem_v, lce_data_mem_v } : 1'b0;
  assign N14 = tl_we;
  assign N15 = N53;
  assign data_mem_addr_li[8:0] = (N14)? pc_gen_icache_vaddr_i[11:3] : 
                                 (N15)? lce_data_mem_pkt[522:514] : 1'b0;
  assign data_mem_addr_li[17:9] = (N14)? pc_gen_icache_vaddr_i[11:3] : 
                                  (N15)? { lce_data_mem_pkt[522:515], N54 } : 1'b0;
  assign data_mem_addr_li[26:18] = (N14)? pc_gen_icache_vaddr_i[11:3] : 
                                   (N15)? { lce_data_mem_pkt[522:516], N55, lce_data_mem_pkt[514:514] } : 1'b0;
  assign data_mem_addr_li[35:27] = (N14)? pc_gen_icache_vaddr_i[11:3] : 
                                   (N15)? { lce_data_mem_pkt[522:516], N56, N57 } : 1'b0;
  assign data_mem_addr_li[44:36] = (N14)? pc_gen_icache_vaddr_i[11:3] : 
                                   (N15)? { lce_data_mem_pkt[522:517], N58, lce_data_mem_pkt[515:514] } : 1'b0;
  assign data_mem_addr_li[53:45] = (N14)? pc_gen_icache_vaddr_i[11:3] : 
                                   (N15)? { lce_data_mem_pkt[522:517], N59, lce_data_mem_pkt[515:515], N60 } : 1'b0;
  assign data_mem_addr_li[62:54] = (N14)? pc_gen_icache_vaddr_i[11:3] : 
                                   (N15)? { lce_data_mem_pkt[522:517], N61, N62, lce_data_mem_pkt[514:514] } : 1'b0;
  assign data_mem_addr_li[71:63] = (N14)? pc_gen_icache_vaddr_i[11:3] : 
                                   (N15)? { lce_data_mem_pkt[522:517], N63, N64, N65 } : 1'b0;
  assign tag_mem_addr_li = (N14)? pc_gen_icache_vaddr_i[11:6] : 
                           (N15)? tag_mem_pkt[39:34] : 1'b0;
  assign tag_mem_w_mask_li = (N16)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                             (N17)? { lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                             (N18)? { lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0] } : 
                             (N19)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N16 = N68;
  assign N17 = N70;
  assign N18 = N72;
  assign N19 = N73;
  assign tag_mem_data_li = (N16)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                           (N17)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                           (N18)? { tag_mem_pkt[30:2], tag_mem_pkt[30:2], tag_mem_pkt[30:2], tag_mem_pkt[30:2], tag_mem_pkt[30:2], tag_mem_pkt[30:2], tag_mem_pkt[30:2], tag_mem_pkt[30:2] } : 
                           (N19)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign stat_mem_w_li = (N10)? N74 : 
                         (N11)? N75 : 1'b0;
  assign stat_mem_addr_li = (N10)? addr_tv_r[11:6] : 
                            (N11)? stat_mem_pkt[9:4] : 1'b0;
  assign stat_mem_data_li = (N10)? lru_decode_data_lo : 
                            (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign stat_mem_mask_li = (N10)? lru_decode_mask_lo : 
                            (N11)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign lce_data_mem_pkt_yumi_li = (N20)? lce_data_mem_pkt_v_lo : 
                                    (N21)? N77 : 1'b0;
  assign N20 = N119;
  assign N21 = N118;
  assign N83 = (N22)? 1'b1 : 
               (N87)? 1'b1 : 
               (N90)? 1'b1 : 
               (N82)? 1'b0 : 1'b0;
  assign N22 = N79;
  assign N84 = (N22)? 1'b0 : 
               (N87)? 1'b1 : 
               (N90)? 1'b0 : 1'b0;
  assign N85 = (N22)? 1'b0 : 
               (N87)? 1'b1 : 
               (N90)? 1'b0 : 
               (N82)? 1'b0 : 1'b0;
  assign tl_we = pc_gen_icache_vaddr_v_i & pc_gen_icache_vaddr_ready_o;
  assign N23 = ~reset_i;
  assign N24 = reset_i;
  assign n_0_net_ = N120 & tag_mem_v_li;
  assign N120 = ~reset_i;
  assign n_1_net_ = N121 & data_mem_v_li[0];
  assign N121 = ~reset_i;
  assign n_2_net_ = N122 & data_mem_v_li[1];
  assign N122 = ~reset_i;
  assign n_3_net_ = N123 & data_mem_v_li[2];
  assign N123 = ~reset_i;
  assign n_4_net_ = N124 & data_mem_v_li[3];
  assign N124 = ~reset_i;
  assign n_5_net_ = N125 & data_mem_v_li[4];
  assign N125 = ~reset_i;
  assign n_6_net_ = N126 & data_mem_v_li[5];
  assign N126 = ~reset_i;
  assign n_7_net_ = N127 & data_mem_v_li[6];
  assign N127 = ~reset_i;
  assign n_8_net_ = N128 & data_mem_v_li[7];
  assign N128 = ~reset_i;
  assign tv_we = N131 & N132;
  assign N131 = N130 & itlb_icache_data_resp_v_i;
  assign N130 = itlb_icache_data_resp_ready_o & N129;
  assign N129 = ~poison_tl_i;
  assign N132 = ~itlb_icache_miss_i;
  assign N27 = ~reset_i;
  assign N28 = reset_i;
  assign hit_v[0] = N39 & N100;
  assign hit_v[1] = N40 & N99;
  assign hit_v[2] = N41 & N98;
  assign hit_v[3] = N42 & N97;
  assign hit_v[4] = N43 & N96;
  assign hit_v[5] = N44 & N95;
  assign hit_v[6] = N45 & N94;
  assign hit_v[7] = N46 & N93;
  assign miss_tv = N134 & N135;
  assign N134 = N133 & v_tv_r;
  assign N133 = ~hit;
  assign N135 = ~uncached_tv_r;
  assign uncached_req = N136 & N137;
  assign N136 = v_tv_r & uncached_tv_r;
  assign N137 = ~uncached_load_data_v_r;
  assign n_9_net_ = N138 & stat_mem_v_li;
  assign N138 = ~reset_i;
  assign n_10_net__7_ = ~N101;
  assign n_10_net__6_ = ~N102;
  assign n_10_net__5_ = ~N103;
  assign n_10_net__4_ = ~N104;
  assign n_10_net__3_ = ~N105;
  assign n_10_net__2_ = ~N106;
  assign n_10_net__1_ = ~N107;
  assign n_10_net__0_ = ~N108;
  assign N47 = ~invalid_exist;
  assign N48 = ~v_tv_r;
  assign N49 = v_tv_r & N139;
  assign N139 = ~cache_miss_o;
  assign n_11_net__2_ = hit_index[2] ^ addr_tv_r[5];
  assign n_11_net__1_ = hit_index[1] ^ addr_tv_r[4];
  assign n_11_net__0_ = hit_index[0] ^ addr_tv_r[3];
  assign N51 = ~addr_tv_r[2];
  assign N52 = addr_tv_r[2];
  assign lce_data_mem_v = N112 & lce_data_mem_pkt_yumi_li;
  assign N53 = ~tl_we;
  assign data_mem_w_li = lce_data_mem_pkt_yumi_li & N92;
  assign N54 = ~lce_data_mem_pkt[514];
  assign N55 = ~lce_data_mem_pkt[515];
  assign N56 = ~lce_data_mem_pkt[515];
  assign N57 = ~lce_data_mem_pkt[514];
  assign N58 = ~lce_data_mem_pkt[516];
  assign N59 = ~lce_data_mem_pkt[516];
  assign N60 = ~lce_data_mem_pkt[514];
  assign N61 = ~lce_data_mem_pkt[516];
  assign N62 = ~lce_data_mem_pkt[515];
  assign N63 = ~lce_data_mem_pkt[516];
  assign N64 = ~lce_data_mem_pkt[515];
  assign N65 = ~lce_data_mem_pkt[514];
  assign tag_mem_v_li = tl_we | tag_mem_pkt_yumi_li;
  assign tag_mem_w_li = N53 & tag_mem_pkt_v_lo;
  assign N66 = ~tag_mem_pkt[1];
  assign N67 = ~tag_mem_pkt[0];
  assign N70 = ~N69;
  assign N72 = ~N71;
  assign stat_mem_v_li = N140 | stat_mem_pkt_yumi_li;
  assign N140 = v_tv_r & N135;
  assign N74 = ~miss_tv;
  assign N75 = stat_mem_pkt_yumi_li & N110;
  assign N76 = lce_data_mem_pkt_yumi_li & N115;
  assign N77 = lce_data_mem_pkt_v_lo & N53;
  assign N78 = lce_data_mem_pkt_yumi_li & N117;
  assign N79 = reset_i;
  assign N80 = N78 | N79;
  assign N81 = icache_pc_gen_data_v_o | N80;
  assign N82 = ~N81;
  assign N86 = ~N79;
  assign N87 = N78 & N86;
  assign N88 = ~N78;
  assign N89 = N86 & N88;
  assign N90 = icache_pc_gen_data_v_o & N89;
  assign tag_mem_pkt_yumi_li = tag_mem_pkt_v_lo & N53;
  assign stat_mem_pkt_yumi_li = N142 & stat_mem_pkt_v_lo;
  assign N142 = ~N141;
  assign N141 = v_tv_r & N135;

  always @(posedge clk_i) begin
    if(N26) begin
      { vaddr_tl_r[38:0] } <= { pc_gen_icache_vaddr_i[38:0] };
    end 
    if(1'b1) begin
      itlb_icache_data_resp_ready_o <= N25;
      v_tv_r <= N29;
    end 
    if(N30) begin
      { ld_data_tv_r[511:414] } <= { data_mem_data_lo[511:414] };
      uncached_tv_r <= uncached_i;
      { addr_tv_r[0:0] } <= { vaddr_tl_r[0:0] };
    end 
    if(N31) begin
      { ld_data_tv_r[413:315] } <= { data_mem_data_lo[413:315] };
      { addr_tv_r[1:1] } <= { vaddr_tl_r[1:1] };
    end 
    if(N32) begin
      { ld_data_tv_r[314:216] } <= { data_mem_data_lo[314:216] };
      { addr_tv_r[2:2] } <= { vaddr_tl_r[2:2] };
    end 
    if(N33) begin
      { ld_data_tv_r[215:117] } <= { data_mem_data_lo[215:117] };
      { addr_tv_r[3:3] } <= { vaddr_tl_r[3:3] };
    end 
    if(N34) begin
      { ld_data_tv_r[116:18] } <= { data_mem_data_lo[116:18] };
      { addr_tv_r[4:4] } <= { vaddr_tl_r[4:4] };
    end 
    if(N35) begin
      { ld_data_tv_r[17:0] } <= { data_mem_data_lo[17:0] };
      { addr_tv_r[5:5] } <= { vaddr_tl_r[5:5] };
      { tag_tv_r[215:151] } <= { tag_mem_data_lo[229:203], tag_mem_data_lo[200:174], tag_mem_data_lo[171:161] };
      { state_tv_r[15:0] } <= { tag_mem_data_lo[231:230], tag_mem_data_lo[202:201], tag_mem_data_lo[173:172], tag_mem_data_lo[144:143], tag_mem_data_lo[115:114], tag_mem_data_lo[86:85], tag_mem_data_lo[57:56], tag_mem_data_lo[28:27] };
    end 
    if(N37) begin
      { addr_tv_r[38:31], addr_tv_r[7:7] } <= { itlb_icache_data_resp_i[26:19], vaddr_tl_r[7:7] };
      { icache_pc_gen_data_o[38:0] } <= { vaddr_tl_r[38:0] };
      { tag_tv_r[51:0] } <= { tag_mem_data_lo[53:29], tag_mem_data_lo[26:0] };
    end 
    if(N38) begin
      { addr_tv_r[30:8] } <= { itlb_icache_data_resp_i[18:0], vaddr_tl_r[11:8] };
    end 
    if(N36) begin
      { addr_tv_r[6:6] } <= { vaddr_tl_r[6:6] };
      { tag_tv_r[150:52] } <= { tag_mem_data_lo[160:145], tag_mem_data_lo[142:116], tag_mem_data_lo[113:87], tag_mem_data_lo[84:58], tag_mem_data_lo[55:54] };
    end 
    if(N76) begin
      { lce_data_mem_pkt_way_r[2:0] } <= { lce_data_mem_pkt[516:514] };
    end 
    if(N85) begin
      { uncached_load_data_r[63:0] } <= { lce_data_mem_pkt[65:2] };
    end 
    if(N83) begin
      uncached_load_data_v_r <= N84;
    end 
  end


endmodule



module bsg_dff_reset_width_p1
(
  clk_i,
  reset_i,
  data_i,
  data_o
);

  input [0:0] data_i;
  output [0:0] data_o;
  input clk_i;
  input reset_i;
  wire N0,N1,N2,N3;
  reg [0:0] data_o;
  assign N3 = (N0)? 1'b0 : 
              (N1)? data_i[0] : 1'b0;
  assign N0 = reset_i;
  assign N1 = N2;
  assign N2 = ~reset_i;

  always @(posedge clk_i) begin
    if(1'b1) begin
      { data_o[0:0] } <= { N3 };
    end 
  end


endmodule



module bsg_dff_reset_width_p27
(
  clk_i,
  reset_i,
  data_i,
  data_o
);

  input [26:0] data_i;
  output [26:0] data_o;
  input clk_i;
  input reset_i;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29;
  reg [26:0] data_o;
  assign { N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3 } = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                              (N1)? data_i : 1'b0;
  assign N0 = reset_i;
  assign N1 = N2;
  assign N2 = ~reset_i;

  always @(posedge clk_i) begin
    if(1'b1) begin
      { data_o[26:0] } <= { N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3 };
    end 
  end


endmodule



module bp_be_dtlb_replacement_ways_p8
(
  clk_i,
  reset_i,
  v_i,
  way_i,
  way_o
);

  input [2:0] way_i;
  output [2:0] way_o;
  input clk_i;
  input reset_i;
  input v_i;
  wire [2:0] way_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26;
  wire [6:0] update_mask,update_data,lru_n;
  reg [6:0] lru_r;

  bsg_lru_pseudo_tree_decode_ways_p8
  decoder
  (
    .way_id_i(way_i),
    .data_o(update_data),
    .mask_o(update_mask)
  );


  bsg_lru_pseudo_tree_encode_ways_p8
  encoder
  (
    .lru_i(lru_r),
    .way_id_o(way_o)
  );

  assign lru_n[0] = (N0)? update_data[0] : 
                    (N8)? lru_r[0] : 1'b0;
  assign N0 = update_mask[0];
  assign lru_n[1] = (N1)? update_data[1] : 
                    (N9)? lru_r[1] : 1'b0;
  assign N1 = update_mask[1];
  assign lru_n[2] = (N2)? update_data[2] : 
                    (N10)? lru_r[2] : 1'b0;
  assign N2 = update_mask[2];
  assign lru_n[3] = (N3)? update_data[3] : 
                    (N11)? lru_r[3] : 1'b0;
  assign N3 = update_mask[3];
  assign lru_n[4] = (N4)? update_data[4] : 
                    (N12)? lru_r[4] : 1'b0;
  assign N4 = update_mask[4];
  assign lru_n[5] = (N5)? update_data[5] : 
                    (N13)? lru_r[5] : 1'b0;
  assign N5 = update_mask[5];
  assign lru_n[6] = (N6)? update_data[6] : 
                    (N14)? lru_r[6] : 1'b0;
  assign N6 = update_mask[6];
  assign N17 = (N7)? 1'b1 : 
               (N26)? 1'b1 : 
               (N16)? 1'b0 : 1'b0;
  assign N7 = reset_i;
  assign { N24, N23, N22, N21, N20, N19, N18 } = (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                 (N26)? lru_n : 1'b0;
  assign N8 = ~update_mask[0];
  assign N9 = ~update_mask[1];
  assign N10 = ~update_mask[2];
  assign N11 = ~update_mask[3];
  assign N12 = ~update_mask[4];
  assign N13 = ~update_mask[5];
  assign N14 = ~update_mask[6];
  assign N15 = v_i | reset_i;
  assign N16 = ~N15;
  assign N25 = ~reset_i;
  assign N26 = v_i & N25;

  always @(posedge clk_i) begin
    if(N17) begin
      { lru_r[6:0] } <= { N24, N23, N22, N21, N20, N19, N18 };
    end 
  end


endmodule



module bsg_cam_1r1w_els_p8_width_p27_multiple_entries_p0_find_empty_entry_p1
(
  clk_i,
  reset_i,
  en_i,
  w_v_i,
  w_set_not_clear_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_data_i,
  r_v_o,
  r_addr_o,
  empty_v_o,
  empty_addr_o
);

  input [2:0] w_addr_i;
  input [26:0] w_data_i;
  input [26:0] r_data_i;
  output [2:0] r_addr_o;
  output [2:0] empty_addr_o;
  input clk_i;
  input reset_i;
  input en_i;
  input w_v_i;
  input w_set_not_clear_i;
  input r_v_i;
  output r_v_o;
  output empty_v_o;
  wire [2:0] r_addr_o,empty_addr_o;
  wire r_v_o,empty_v_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,matched,empty_found,N9,N10,N11,N12,
  N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,
  N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,
  N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,
  N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84;
  wire [7:0] match_array,empty_array;
  reg [215:0] mem;
  reg [7:0] valid;
  assign N39 = mem[215:189] == r_data_i;
  assign N40 = mem[188:162] == r_data_i;
  assign N41 = mem[161:135] == r_data_i;
  assign N42 = mem[134:108] == r_data_i;
  assign N43 = mem[107:81] == r_data_i;
  assign N44 = mem[80:54] == r_data_i;
  assign N45 = mem[53:27] == r_data_i;
  assign N46 = mem[26:0] == r_data_i;

  bsg_encode_one_hot_width_p8_lo_to_hi_p1
  fi4_ohe
  (
    .i(match_array),
    .addr_o(r_addr_o),
    .v_o(matched)
  );


  bsg_priority_encode_width_p8_lo_to_hi_p1
  fi5_epe
  (
    .i(empty_array),
    .addr_o(empty_addr_o),
    .v_o(empty_found)
  );

  assign N19 = N47 & w_addr_i[2];
  assign N18 = N48 & w_addr_i[2];
  assign N17 = N49 & w_addr_i[2];
  assign N16 = N50 & w_addr_i[2];
  assign N47 = w_addr_i[0] & w_addr_i[1];
  assign N15 = N47 & N0;
  assign N0 = ~w_addr_i[2];
  assign N48 = N1 & w_addr_i[1];
  assign N1 = ~w_addr_i[0];
  assign N14 = N48 & N2;
  assign N2 = ~w_addr_i[2];
  assign N49 = w_addr_i[0] & N3;
  assign N3 = ~w_addr_i[1];
  assign N13 = N49 & N4;
  assign N4 = ~w_addr_i[2];
  assign N50 = N5 & N6;
  assign N5 = ~w_addr_i[0];
  assign N6 = ~w_addr_i[1];
  assign N12 = N50 & N7;
  assign N7 = ~w_addr_i[2];
  assign { N28, N27, N26, N25, N24, N23, N22, N20 } = (N8)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                                                      (N38)? { N19, N18, N17, N16, N15, N14, N13, N12 } : 
                                                      (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N8 = reset_i;
  assign N21 = (N8)? 1'b0 : 
               (N38)? w_set_not_clear_i : 1'b0;
  assign { N36, N35, N34, N33, N32, N31, N30, N29 } = (N8)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                      (N38)? { N12, N13, N14, N15, N16, N17, N18, N19 } : 
                                                      (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign r_v_o = N51 & matched;
  assign N51 = en_i & r_v_i;
  assign empty_v_o = en_i & empty_found;
  assign N9 = en_i & w_v_i;
  assign N10 = N9 | reset_i;
  assign N11 = ~N10;
  assign N37 = ~reset_i;
  assign N38 = N9 & N37;
  assign match_array[0] = N54 & valid[0];
  assign N54 = N53 & N39;
  assign N53 = N52 & en_i;
  assign N52 = ~reset_i;
  assign empty_array[0] = N55 & N56;
  assign N55 = N52 & en_i;
  assign N56 = ~valid[0];
  assign match_array[1] = N58 & valid[1];
  assign N58 = N57 & N40;
  assign N57 = N52 & en_i;
  assign empty_array[1] = N59 & N60;
  assign N59 = N52 & en_i;
  assign N60 = ~valid[1];
  assign match_array[2] = N62 & valid[2];
  assign N62 = N61 & N41;
  assign N61 = N52 & en_i;
  assign empty_array[2] = N63 & N64;
  assign N63 = N52 & en_i;
  assign N64 = ~valid[2];
  assign match_array[3] = N66 & valid[3];
  assign N66 = N65 & N42;
  assign N65 = N52 & en_i;
  assign empty_array[3] = N67 & N68;
  assign N67 = N52 & en_i;
  assign N68 = ~valid[3];
  assign match_array[4] = N70 & valid[4];
  assign N70 = N69 & N43;
  assign N69 = N52 & en_i;
  assign empty_array[4] = N71 & N72;
  assign N71 = N52 & en_i;
  assign N72 = ~valid[4];
  assign match_array[5] = N74 & valid[5];
  assign N74 = N73 & N44;
  assign N73 = N52 & en_i;
  assign empty_array[5] = N75 & N76;
  assign N75 = N52 & en_i;
  assign N76 = ~valid[5];
  assign match_array[6] = N78 & valid[6];
  assign N78 = N77 & N45;
  assign N77 = N52 & en_i;
  assign empty_array[6] = N79 & N80;
  assign N79 = N52 & en_i;
  assign N80 = ~valid[6];
  assign match_array[7] = N82 & valid[7];
  assign N82 = N81 & N46;
  assign N81 = N52 & en_i;
  assign empty_array[7] = N83 & N84;
  assign N83 = N52 & en_i;
  assign N84 = ~valid[7];

  always @(posedge clk_i) begin
    if(N36) begin
      { mem[215:189] } <= { w_data_i[26:0] };
    end 
    if(N35) begin
      { mem[188:162] } <= { w_data_i[26:0] };
    end 
    if(N34) begin
      { mem[161:135] } <= { w_data_i[26:0] };
    end 
    if(N33) begin
      { mem[134:108] } <= { w_data_i[26:0] };
    end 
    if(N32) begin
      { mem[107:81] } <= { w_data_i[26:0] };
    end 
    if(N31) begin
      { mem[80:54] } <= { w_data_i[26:0] };
    end 
    if(N30) begin
      { mem[53:27] } <= { w_data_i[26:0] };
    end 
    if(N29) begin
      { mem[26:0] } <= { w_data_i[26:0] };
    end 
    if(N28) begin
      { valid[7:7] } <= { N21 };
    end 
    if(N27) begin
      { valid[6:6] } <= { N21 };
    end 
    if(N26) begin
      { valid[5:5] } <= { N21 };
    end 
    if(N25) begin
      { valid[4:4] } <= { N21 };
    end 
    if(N24) begin
      { valid[3:3] } <= { N21 };
    end 
    if(N23) begin
      { valid[2:2] } <= { N21 };
    end 
    if(N22) begin
      { valid[1:1] } <= { N21 };
    end 
    if(N20) begin
      { valid[0:0] } <= { N21 };
    end 
  end


endmodule



module bsg_mem_1r1w_synth_width_p33_els_p8_read_write_same_addr_p0_harden_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [2:0] w_addr_i;
  input [32:0] w_data_i;
  input [2:0] r_addr_i;
  output [32:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [32:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45;
  reg [263:0] mem;
  assign r_data_o[32] = (N17)? mem[32] : 
                        (N19)? mem[65] : 
                        (N21)? mem[98] : 
                        (N23)? mem[131] : 
                        (N18)? mem[164] : 
                        (N20)? mem[197] : 
                        (N22)? mem[230] : 
                        (N24)? mem[263] : 1'b0;
  assign r_data_o[31] = (N17)? mem[31] : 
                        (N19)? mem[64] : 
                        (N21)? mem[97] : 
                        (N23)? mem[130] : 
                        (N18)? mem[163] : 
                        (N20)? mem[196] : 
                        (N22)? mem[229] : 
                        (N24)? mem[262] : 1'b0;
  assign r_data_o[30] = (N17)? mem[30] : 
                        (N19)? mem[63] : 
                        (N21)? mem[96] : 
                        (N23)? mem[129] : 
                        (N18)? mem[162] : 
                        (N20)? mem[195] : 
                        (N22)? mem[228] : 
                        (N24)? mem[261] : 1'b0;
  assign r_data_o[29] = (N17)? mem[29] : 
                        (N19)? mem[62] : 
                        (N21)? mem[95] : 
                        (N23)? mem[128] : 
                        (N18)? mem[161] : 
                        (N20)? mem[194] : 
                        (N22)? mem[227] : 
                        (N24)? mem[260] : 1'b0;
  assign r_data_o[28] = (N17)? mem[28] : 
                        (N19)? mem[61] : 
                        (N21)? mem[94] : 
                        (N23)? mem[127] : 
                        (N18)? mem[160] : 
                        (N20)? mem[193] : 
                        (N22)? mem[226] : 
                        (N24)? mem[259] : 1'b0;
  assign r_data_o[27] = (N17)? mem[27] : 
                        (N19)? mem[60] : 
                        (N21)? mem[93] : 
                        (N23)? mem[126] : 
                        (N18)? mem[159] : 
                        (N20)? mem[192] : 
                        (N22)? mem[225] : 
                        (N24)? mem[258] : 1'b0;
  assign r_data_o[26] = (N17)? mem[26] : 
                        (N19)? mem[59] : 
                        (N21)? mem[92] : 
                        (N23)? mem[125] : 
                        (N18)? mem[158] : 
                        (N20)? mem[191] : 
                        (N22)? mem[224] : 
                        (N24)? mem[257] : 1'b0;
  assign r_data_o[25] = (N17)? mem[25] : 
                        (N19)? mem[58] : 
                        (N21)? mem[91] : 
                        (N23)? mem[124] : 
                        (N18)? mem[157] : 
                        (N20)? mem[190] : 
                        (N22)? mem[223] : 
                        (N24)? mem[256] : 1'b0;
  assign r_data_o[24] = (N17)? mem[24] : 
                        (N19)? mem[57] : 
                        (N21)? mem[90] : 
                        (N23)? mem[123] : 
                        (N18)? mem[156] : 
                        (N20)? mem[189] : 
                        (N22)? mem[222] : 
                        (N24)? mem[255] : 1'b0;
  assign r_data_o[23] = (N17)? mem[23] : 
                        (N19)? mem[56] : 
                        (N21)? mem[89] : 
                        (N23)? mem[122] : 
                        (N18)? mem[155] : 
                        (N20)? mem[188] : 
                        (N22)? mem[221] : 
                        (N24)? mem[254] : 1'b0;
  assign r_data_o[22] = (N17)? mem[22] : 
                        (N19)? mem[55] : 
                        (N21)? mem[88] : 
                        (N23)? mem[121] : 
                        (N18)? mem[154] : 
                        (N20)? mem[187] : 
                        (N22)? mem[220] : 
                        (N24)? mem[253] : 1'b0;
  assign r_data_o[21] = (N17)? mem[21] : 
                        (N19)? mem[54] : 
                        (N21)? mem[87] : 
                        (N23)? mem[120] : 
                        (N18)? mem[153] : 
                        (N20)? mem[186] : 
                        (N22)? mem[219] : 
                        (N24)? mem[252] : 1'b0;
  assign r_data_o[20] = (N17)? mem[20] : 
                        (N19)? mem[53] : 
                        (N21)? mem[86] : 
                        (N23)? mem[119] : 
                        (N18)? mem[152] : 
                        (N20)? mem[185] : 
                        (N22)? mem[218] : 
                        (N24)? mem[251] : 1'b0;
  assign r_data_o[19] = (N17)? mem[19] : 
                        (N19)? mem[52] : 
                        (N21)? mem[85] : 
                        (N23)? mem[118] : 
                        (N18)? mem[151] : 
                        (N20)? mem[184] : 
                        (N22)? mem[217] : 
                        (N24)? mem[250] : 1'b0;
  assign r_data_o[18] = (N17)? mem[18] : 
                        (N19)? mem[51] : 
                        (N21)? mem[84] : 
                        (N23)? mem[117] : 
                        (N18)? mem[150] : 
                        (N20)? mem[183] : 
                        (N22)? mem[216] : 
                        (N24)? mem[249] : 1'b0;
  assign r_data_o[17] = (N17)? mem[17] : 
                        (N19)? mem[50] : 
                        (N21)? mem[83] : 
                        (N23)? mem[116] : 
                        (N18)? mem[149] : 
                        (N20)? mem[182] : 
                        (N22)? mem[215] : 
                        (N24)? mem[248] : 1'b0;
  assign r_data_o[16] = (N17)? mem[16] : 
                        (N19)? mem[49] : 
                        (N21)? mem[82] : 
                        (N23)? mem[115] : 
                        (N18)? mem[148] : 
                        (N20)? mem[181] : 
                        (N22)? mem[214] : 
                        (N24)? mem[247] : 1'b0;
  assign r_data_o[15] = (N17)? mem[15] : 
                        (N19)? mem[48] : 
                        (N21)? mem[81] : 
                        (N23)? mem[114] : 
                        (N18)? mem[147] : 
                        (N20)? mem[180] : 
                        (N22)? mem[213] : 
                        (N24)? mem[246] : 1'b0;
  assign r_data_o[14] = (N17)? mem[14] : 
                        (N19)? mem[47] : 
                        (N21)? mem[80] : 
                        (N23)? mem[113] : 
                        (N18)? mem[146] : 
                        (N20)? mem[179] : 
                        (N22)? mem[212] : 
                        (N24)? mem[245] : 1'b0;
  assign r_data_o[13] = (N17)? mem[13] : 
                        (N19)? mem[46] : 
                        (N21)? mem[79] : 
                        (N23)? mem[112] : 
                        (N18)? mem[145] : 
                        (N20)? mem[178] : 
                        (N22)? mem[211] : 
                        (N24)? mem[244] : 1'b0;
  assign r_data_o[12] = (N17)? mem[12] : 
                        (N19)? mem[45] : 
                        (N21)? mem[78] : 
                        (N23)? mem[111] : 
                        (N18)? mem[144] : 
                        (N20)? mem[177] : 
                        (N22)? mem[210] : 
                        (N24)? mem[243] : 1'b0;
  assign r_data_o[11] = (N17)? mem[11] : 
                        (N19)? mem[44] : 
                        (N21)? mem[77] : 
                        (N23)? mem[110] : 
                        (N18)? mem[143] : 
                        (N20)? mem[176] : 
                        (N22)? mem[209] : 
                        (N24)? mem[242] : 1'b0;
  assign r_data_o[10] = (N17)? mem[10] : 
                        (N19)? mem[43] : 
                        (N21)? mem[76] : 
                        (N23)? mem[109] : 
                        (N18)? mem[142] : 
                        (N20)? mem[175] : 
                        (N22)? mem[208] : 
                        (N24)? mem[241] : 1'b0;
  assign r_data_o[9] = (N17)? mem[9] : 
                       (N19)? mem[42] : 
                       (N21)? mem[75] : 
                       (N23)? mem[108] : 
                       (N18)? mem[141] : 
                       (N20)? mem[174] : 
                       (N22)? mem[207] : 
                       (N24)? mem[240] : 1'b0;
  assign r_data_o[8] = (N17)? mem[8] : 
                       (N19)? mem[41] : 
                       (N21)? mem[74] : 
                       (N23)? mem[107] : 
                       (N18)? mem[140] : 
                       (N20)? mem[173] : 
                       (N22)? mem[206] : 
                       (N24)? mem[239] : 1'b0;
  assign r_data_o[7] = (N17)? mem[7] : 
                       (N19)? mem[40] : 
                       (N21)? mem[73] : 
                       (N23)? mem[106] : 
                       (N18)? mem[139] : 
                       (N20)? mem[172] : 
                       (N22)? mem[205] : 
                       (N24)? mem[238] : 1'b0;
  assign r_data_o[6] = (N17)? mem[6] : 
                       (N19)? mem[39] : 
                       (N21)? mem[72] : 
                       (N23)? mem[105] : 
                       (N18)? mem[138] : 
                       (N20)? mem[171] : 
                       (N22)? mem[204] : 
                       (N24)? mem[237] : 1'b0;
  assign r_data_o[5] = (N17)? mem[5] : 
                       (N19)? mem[38] : 
                       (N21)? mem[71] : 
                       (N23)? mem[104] : 
                       (N18)? mem[137] : 
                       (N20)? mem[170] : 
                       (N22)? mem[203] : 
                       (N24)? mem[236] : 1'b0;
  assign r_data_o[4] = (N17)? mem[4] : 
                       (N19)? mem[37] : 
                       (N21)? mem[70] : 
                       (N23)? mem[103] : 
                       (N18)? mem[136] : 
                       (N20)? mem[169] : 
                       (N22)? mem[202] : 
                       (N24)? mem[235] : 1'b0;
  assign r_data_o[3] = (N17)? mem[3] : 
                       (N19)? mem[36] : 
                       (N21)? mem[69] : 
                       (N23)? mem[102] : 
                       (N18)? mem[135] : 
                       (N20)? mem[168] : 
                       (N22)? mem[201] : 
                       (N24)? mem[234] : 1'b0;
  assign r_data_o[2] = (N17)? mem[2] : 
                       (N19)? mem[35] : 
                       (N21)? mem[68] : 
                       (N23)? mem[101] : 
                       (N18)? mem[134] : 
                       (N20)? mem[167] : 
                       (N22)? mem[200] : 
                       (N24)? mem[233] : 1'b0;
  assign r_data_o[1] = (N17)? mem[1] : 
                       (N19)? mem[34] : 
                       (N21)? mem[67] : 
                       (N23)? mem[100] : 
                       (N18)? mem[133] : 
                       (N20)? mem[166] : 
                       (N22)? mem[199] : 
                       (N24)? mem[232] : 1'b0;
  assign r_data_o[0] = (N17)? mem[0] : 
                       (N19)? mem[33] : 
                       (N21)? mem[66] : 
                       (N23)? mem[99] : 
                       (N18)? mem[132] : 
                       (N20)? mem[165] : 
                       (N22)? mem[198] : 
                       (N24)? mem[231] : 1'b0;
  assign N42 = w_addr_i[0] & w_addr_i[1];
  assign N33 = N42 & w_addr_i[2];
  assign N43 = N0 & w_addr_i[1];
  assign N0 = ~w_addr_i[0];
  assign N32 = N43 & w_addr_i[2];
  assign N44 = w_addr_i[0] & N1;
  assign N1 = ~w_addr_i[1];
  assign N31 = N44 & w_addr_i[2];
  assign N45 = N2 & N3;
  assign N2 = ~w_addr_i[0];
  assign N3 = ~w_addr_i[1];
  assign N30 = N45 & w_addr_i[2];
  assign N29 = N42 & N4;
  assign N4 = ~w_addr_i[2];
  assign N28 = N43 & N5;
  assign N5 = ~w_addr_i[2];
  assign N27 = N44 & N6;
  assign N6 = ~w_addr_i[2];
  assign N26 = N45 & N7;
  assign N7 = ~w_addr_i[2];
  assign { N41, N40, N39, N38, N37, N36, N35, N34 } = (N8)? { N33, N32, N31, N30, N29, N28, N27, N26 } : 
                                                      (N9)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N8 = w_v_i;
  assign N9 = N25;
  assign N10 = ~r_addr_i[0];
  assign N11 = ~r_addr_i[1];
  assign N12 = N10 & N11;
  assign N13 = N10 & r_addr_i[1];
  assign N14 = r_addr_i[0] & N11;
  assign N15 = r_addr_i[0] & r_addr_i[1];
  assign N16 = ~r_addr_i[2];
  assign N17 = N12 & N16;
  assign N18 = N12 & r_addr_i[2];
  assign N19 = N14 & N16;
  assign N20 = N14 & r_addr_i[2];
  assign N21 = N13 & N16;
  assign N22 = N13 & r_addr_i[2];
  assign N23 = N15 & N16;
  assign N24 = N15 & r_addr_i[2];
  assign N25 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N41) begin
      { mem[263:231] } <= { w_data_i[32:0] };
    end 
    if(N40) begin
      { mem[230:198] } <= { w_data_i[32:0] };
    end 
    if(N39) begin
      { mem[197:165] } <= { w_data_i[32:0] };
    end 
    if(N38) begin
      { mem[164:132] } <= { w_data_i[32:0] };
    end 
    if(N37) begin
      { mem[131:99] } <= { w_data_i[32:0] };
    end 
    if(N36) begin
      { mem[98:66] } <= { w_data_i[32:0] };
    end 
    if(N35) begin
      { mem[65:33] } <= { w_data_i[32:0] };
    end 
    if(N34) begin
      { mem[32:0] } <= { w_data_i[32:0] };
    end 
  end


endmodule



module bsg_mem_1r1w_width_p33_els_p8_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [2:0] w_addr_i;
  input [32:0] w_data_i;
  input [2:0] r_addr_i;
  output [32:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [32:0] r_data_o;

  bsg_mem_1r1w_synth_width_p33_els_p8_read_write_same_addr_p0_harden_p0
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_mem_1rw_sync_width_p33_els_p8
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_i,
  data_o
);

  input [32:0] data_i;
  input [2:0] addr_i;
  output [32:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire n_0_net_,n_1_net_,N0;
  wire [32:0] z_s1r1w_data_lo;
  reg [32:0] data_o;

  bsg_mem_1r1w_width_p33_els_p8_read_write_same_addr_p0
  z_s1r1w_mem
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(n_0_net_),
    .w_addr_i(addr_i),
    .w_data_i(data_i),
    .r_v_i(n_1_net_),
    .r_addr_i(addr_i),
    .r_data_o(z_s1r1w_data_lo)
  );

  assign n_1_net_ = v_i & N0;
  assign N0 = ~w_i;
  assign n_0_net_ = v_i & w_i;

  always @(posedge clk_i) begin
    if(1'b1) begin
      { data_o[32:0] } <= { z_s1r1w_data_lo[32:0] };
    end 
  end


endmodule



module bp_be_dtlb_02
(
  clk_i,
  reset_i,
  flush_i,
  r_v_i,
  r_ready_o,
  r_vtag_i,
  r_v_o,
  r_entry_o,
  w_v_i,
  w_vtag_i,
  w_entry_i,
  miss_v_o,
  miss_vtag_o
);

  input [26:0] r_vtag_i;
  output [32:0] r_entry_o;
  input [26:0] w_vtag_i;
  input [32:0] w_entry_i;
  output [26:0] miss_vtag_o;
  input clk_i;
  input reset_i;
  input flush_i;
  input r_v_i;
  input w_v_i;
  output r_ready_o;
  output r_v_o;
  output miss_v_o;
  wire [32:0] r_entry_o;
  wire [26:0] miss_vtag_o;
  wire r_ready_o,r_v_o,miss_v_o,N0,N1,N2,N3,cam_r_v,r_v_n,miss_v_n,n_0_net_,n_1_net_,
  n_4_net_,N4,SYNOPSYS_UNCONNECTED_1,SYNOPSYS_UNCONNECTED_2,SYNOPSYS_UNCONNECTED_3;
  wire [2:0] cam_w_addr,ram_addr,cam_r_addr;

  bsg_dff_reset_width_p1
  r_v_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(r_v_n),
    .data_o(r_v_o)
  );


  bsg_dff_reset_width_p1
  miss_v_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(miss_v_n),
    .data_o(miss_v_o)
  );


  bsg_dff_reset_width_p27
  miss_vtag_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(r_vtag_i),
    .data_o(miss_vtag_o)
  );


  bp_be_dtlb_replacement_ways_p8
  plru
  (
    .clk_i(clk_i),
    .reset_i(n_0_net_),
    .v_i(cam_r_v),
    .way_i(cam_r_addr),
    .way_o(cam_w_addr)
  );


  bsg_cam_1r1w_els_p8_width_p27_multiple_entries_p0_find_empty_entry_p1
  vtag_cam
  (
    .clk_i(clk_i),
    .reset_i(n_1_net_),
    .en_i(1'b1),
    .w_v_i(w_v_i),
    .w_set_not_clear_i(1'b1),
    .w_addr_i(cam_w_addr),
    .w_data_i(w_vtag_i),
    .r_v_i(r_v_i),
    .r_data_i(r_vtag_i),
    .r_v_o(cam_r_v),
    .r_addr_o(cam_r_addr),
    .empty_addr_o({ SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3 })
  );


  bsg_mem_1rw_sync_width_p33_els_p8
  entry_ram
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(w_entry_i),
    .addr_i(ram_addr),
    .v_i(n_4_net_),
    .w_i(w_v_i),
    .data_o(r_entry_o)
  );

  assign ram_addr = (N0)? cam_w_addr : 
                    (N1)? cam_r_addr : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign r_ready_o = ~w_v_i;
  assign N2 = ~w_v_i;
  assign N3 = w_v_i;
  assign r_v_n = r_v_i & cam_r_v;
  assign miss_v_n = r_v_i & N4;
  assign N4 = ~cam_r_v;
  assign n_0_net_ = reset_i | flush_i;
  assign n_1_net_ = reset_i | flush_i;
  assign n_4_net_ = cam_r_v | w_v_i;

endmodule



module bp_fe_top
(
  clk_i,
  reset_i,
  freeze_i,
  icache_id_i,
  cfg_w_v_i,
  cfg_addr_i,
  cfg_data_i,
  fe_cmd_i,
  fe_cmd_v_i,
  fe_cmd_ready_o,
  fe_queue_o,
  fe_queue_v_o,
  fe_queue_ready_i,
  lce_req_o,
  lce_req_v_o,
  lce_req_ready_i,
  lce_resp_o,
  lce_resp_v_o,
  lce_resp_ready_i,
  lce_data_resp_o,
  lce_data_resp_v_o,
  lce_data_resp_ready_i,
  lce_cmd_i,
  lce_cmd_v_i,
  lce_cmd_ready_o,
  lce_data_cmd_i,
  lce_data_cmd_v_i,
  lce_data_cmd_ready_o,
  lce_data_cmd_o,
  lce_data_cmd_v_o,
  lce_data_cmd_ready_i
);

  input [0:0] icache_id_i;
  input [15:0] cfg_addr_i;
  input [31:0] cfg_data_i;
  input [75:0] fe_cmd_i;
  output [99:0] fe_queue_o;
  output [113:0] lce_req_o;
  output [42:0] lce_resp_o;
  output [553:0] lce_data_resp_o;
  input [52:0] lce_cmd_i;
  input [517:0] lce_data_cmd_i;
  output [517:0] lce_data_cmd_o;
  input clk_i;
  input reset_i;
  input freeze_i;
  input cfg_w_v_i;
  input fe_cmd_v_i;
  input fe_queue_ready_i;
  input lce_req_ready_i;
  input lce_resp_ready_i;
  input lce_data_resp_ready_i;
  input lce_cmd_v_i;
  input lce_data_cmd_v_i;
  input lce_data_cmd_ready_i;
  output fe_cmd_ready_o;
  output fe_queue_v_o;
  output lce_req_v_o;
  output lce_resp_v_o;
  output lce_data_resp_v_o;
  output lce_cmd_ready_o;
  output lce_data_cmd_ready_o;
  output lce_data_cmd_v_o;
  wire [99:0] fe_queue_o;
  wire [113:0] lce_req_o;
  wire [42:0] lce_resp_o;
  wire [553:0] lce_data_resp_o;
  wire [517:0] lce_data_cmd_o;
  wire fe_cmd_ready_o,fe_queue_v_o,lce_req_v_o,lce_resp_v_o,lce_data_resp_v_o,
  lce_cmd_ready_o,lce_data_cmd_ready_o,lce_data_cmd_v_o,N0,N1,N2,N3,
  pc_gen_queue_scan_instr__68_,pc_gen_queue_scan_instr__67_,pc_gen_queue_scan_instr__66_,
  pc_gen_queue_scan_instr__65_,pc_gen_queue_scan_instr__64_,pc_gen_queue_scan_instr__63_,
  pc_gen_queue_scan_instr__62_,pc_gen_queue_scan_instr__61_,pc_gen_queue_scan_instr__60_,
  pc_gen_queue_scan_instr__59_,pc_gen_queue_scan_instr__58_,
  pc_gen_queue_scan_instr__57_,pc_gen_queue_scan_instr__56_,pc_gen_queue_scan_instr__55_,
  pc_gen_queue_scan_instr__54_,pc_gen_queue_scan_instr__53_,pc_gen_queue_scan_instr__52_,
  pc_gen_queue_scan_instr__51_,pc_gen_queue_scan_instr__50_,pc_gen_queue_scan_instr__49_,
  pc_gen_queue_scan_instr__48_,pc_gen_queue_scan_instr__47_,
  pc_gen_queue_scan_instr__46_,pc_gen_queue_scan_instr__45_,pc_gen_queue_scan_instr__44_,
  pc_gen_queue_scan_instr__43_,pc_gen_queue_scan_instr__42_,pc_gen_queue_scan_instr__41_,
  pc_gen_queue_scan_instr__40_,pc_gen_queue_scan_instr__39_,pc_gen_queue_scan_instr__38_,
  pc_gen_queue_scan_instr__37_,pc_gen_queue_scan_instr__36_,
  pc_gen_queue_scan_instr__35_,pc_gen_queue_scan_instr__34_,pc_gen_queue_scan_instr__33_,
  pc_gen_queue_scan_instr__32_,pc_gen_queue_scan_instr__31_,pc_gen_queue_scan_instr__30_,
  pc_gen_queue_scan_instr__29_,pc_gen_queue_scan_instr__28_,pc_gen_queue_scan_instr__27_,
  pc_gen_queue_scan_instr__26_,pc_gen_queue_scan_instr__25_,
  pc_gen_queue_scan_instr__24_,pc_gen_queue_scan_instr__23_,pc_gen_queue_scan_instr__22_,
  pc_gen_queue_scan_instr__21_,pc_gen_queue_scan_instr__20_,pc_gen_queue_scan_instr__19_,
  pc_gen_queue_scan_instr__18_,pc_gen_queue_scan_instr__17_,pc_gen_queue_scan_instr__16_,
  pc_gen_queue_scan_instr__15_,pc_gen_queue_scan_instr__14_,
  pc_gen_queue_scan_instr__13_,pc_gen_queue_scan_instr__12_,pc_gen_queue_scan_instr__11_,
  pc_gen_queue_scan_instr__10_,pc_gen_queue_scan_instr__9_,pc_gen_queue_scan_instr__8_,
  pc_gen_queue_scan_instr__7_,pc_gen_queue_scan_instr__6_,pc_gen_queue_scan_instr__5_,
  pc_gen_queue_scan_instr__4_,pc_gen_queue_scan_instr__3_,pc_gen_queue_scan_instr__2_,
  pc_gen_queue_scan_instr__1_,pc_gen_queue_scan_instr__0_,
  fe_pc_gen_branch_metadata_fwd__26_,fe_pc_gen_branch_metadata_fwd__25_,fe_pc_gen_branch_metadata_fwd__24_,
  fe_pc_gen_branch_metadata_fwd__23_,fe_pc_gen_branch_metadata_fwd__22_,
  fe_pc_gen_branch_metadata_fwd__21_,fe_pc_gen_branch_metadata_fwd__20_,
  fe_pc_gen_branch_metadata_fwd__19_,fe_pc_gen_branch_metadata_fwd__18_,fe_pc_gen_branch_metadata_fwd__17_,
  fe_pc_gen_branch_metadata_fwd__16_,fe_pc_gen_branch_metadata_fwd__15_,
  fe_pc_gen_branch_metadata_fwd__14_,fe_pc_gen_branch_metadata_fwd__13_,
  fe_pc_gen_branch_metadata_fwd__12_,fe_pc_gen_branch_metadata_fwd__11_,
  fe_pc_gen_branch_metadata_fwd__10_,fe_pc_gen_branch_metadata_fwd__9_,fe_pc_gen_branch_metadata_fwd__8_,
  fe_pc_gen_branch_metadata_fwd__7_,fe_pc_gen_branch_metadata_fwd__6_,
  fe_pc_gen_branch_metadata_fwd__5_,fe_pc_gen_branch_metadata_fwd__4_,
  fe_pc_gen_branch_metadata_fwd__3_,fe_pc_gen_branch_metadata_fwd__2_,fe_pc_gen_branch_metadata_fwd__1_,
  fe_pc_gen_branch_metadata_fwd__0_,fe_pc_gen_pc_redirect_valid_,N4,N5,icache_miss,poison_tl,
  itlb_entry_r_g_,itlb_entry_r_u_,itlb_entry_r_x_,itlb_entry_r_w_,itlb_entry_r_r_,
  itlb_entry_r_uc_,itlb_fill_v,itlb_w_v,itlb_fence_v,N6,N7,N8,pc_gen_icache_v,
  pc_gen_icache_ready,icache_pc_gen_v,icache_pc_gen_ready,instr_access_fault,
  pc_gen_itlb_v,pc_gen_itlb_ready,itlb_miss,itlb_icache_data_resp_v,
  itlb_icache_data_resp_ready,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,
  N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43;
  wire [38:0] itlb_vaddr,pc_gen_icache;
  wire [26:0] itlb_icache,itlb_miss_vtag;
  wire [70:0] icache_pc_gen;
  reg itlb_fill_r;

  bp_fe_pc_gen_02
  bp_fe_pc_gen_1
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .pc_gen_icache_o(pc_gen_icache),
    .pc_gen_icache_v_o(pc_gen_icache_v),
    .pc_gen_icache_ready_i(pc_gen_icache_ready),
    .icache_pc_gen_i(icache_pc_gen),
    .icache_pc_gen_v_i(icache_pc_gen_v),
    .icache_pc_gen_ready_o(icache_pc_gen_ready),
    .icache_miss_i(icache_miss),
    .instr_access_fault_i(instr_access_fault),
    .pc_gen_itlb_o(itlb_vaddr),
    .pc_gen_itlb_v_o(pc_gen_itlb_v),
    .pc_gen_itlb_ready_i(pc_gen_itlb_ready),
    .pc_gen_fe_o({ fe_queue_o[99:99], pc_gen_queue_scan_instr__68_, pc_gen_queue_scan_instr__67_, pc_gen_queue_scan_instr__66_, pc_gen_queue_scan_instr__65_, pc_gen_queue_scan_instr__64_, pc_gen_queue_scan_instr__63_, pc_gen_queue_scan_instr__62_, pc_gen_queue_scan_instr__61_, pc_gen_queue_scan_instr__60_, pc_gen_queue_scan_instr__59_, pc_gen_queue_scan_instr__58_, pc_gen_queue_scan_instr__57_, pc_gen_queue_scan_instr__56_, pc_gen_queue_scan_instr__55_, pc_gen_queue_scan_instr__54_, pc_gen_queue_scan_instr__53_, pc_gen_queue_scan_instr__52_, pc_gen_queue_scan_instr__51_, pc_gen_queue_scan_instr__50_, pc_gen_queue_scan_instr__49_, pc_gen_queue_scan_instr__48_, pc_gen_queue_scan_instr__47_, pc_gen_queue_scan_instr__46_, pc_gen_queue_scan_instr__45_, pc_gen_queue_scan_instr__44_, pc_gen_queue_scan_instr__43_, pc_gen_queue_scan_instr__42_, pc_gen_queue_scan_instr__41_, pc_gen_queue_scan_instr__40_, pc_gen_queue_scan_instr__39_, pc_gen_queue_scan_instr__38_, pc_gen_queue_scan_instr__37_, pc_gen_queue_scan_instr__36_, pc_gen_queue_scan_instr__35_, pc_gen_queue_scan_instr__34_, pc_gen_queue_scan_instr__33_, pc_gen_queue_scan_instr__32_, pc_gen_queue_scan_instr__31_, pc_gen_queue_scan_instr__30_, pc_gen_queue_scan_instr__29_, pc_gen_queue_scan_instr__28_, pc_gen_queue_scan_instr__27_, pc_gen_queue_scan_instr__26_, pc_gen_queue_scan_instr__25_, pc_gen_queue_scan_instr__24_, pc_gen_queue_scan_instr__23_, pc_gen_queue_scan_instr__22_, pc_gen_queue_scan_instr__21_, pc_gen_queue_scan_instr__20_, pc_gen_queue_scan_instr__19_, pc_gen_queue_scan_instr__18_, pc_gen_queue_scan_instr__17_, pc_gen_queue_scan_instr__16_, pc_gen_queue_scan_instr__15_, pc_gen_queue_scan_instr__14_, pc_gen_queue_scan_instr__13_, pc_gen_queue_scan_instr__12_, pc_gen_queue_scan_instr__11_, pc_gen_queue_scan_instr__10_, pc_gen_queue_scan_instr__9_, pc_gen_queue_scan_instr__8_, pc_gen_queue_scan_instr__7_, pc_gen_queue_scan_instr__6_, pc_gen_queue_scan_instr__5_, pc_gen_queue_scan_instr__4_, pc_gen_queue_scan_instr__3_, pc_gen_queue_scan_instr__2_, pc_gen_queue_scan_instr__1_, pc_gen_queue_scan_instr__0_, fe_queue_o[98:0] }),
    .pc_gen_fe_v_o(fe_queue_v_o),
    .pc_gen_fe_ready_i(fe_queue_ready_i),
    .fe_pc_gen_i({ fe_cmd_i[72:34], fe_pc_gen_branch_metadata_fwd__26_, fe_pc_gen_branch_metadata_fwd__25_, fe_pc_gen_branch_metadata_fwd__24_, fe_pc_gen_branch_metadata_fwd__23_, fe_pc_gen_branch_metadata_fwd__22_, fe_pc_gen_branch_metadata_fwd__21_, fe_pc_gen_branch_metadata_fwd__20_, fe_pc_gen_branch_metadata_fwd__19_, fe_pc_gen_branch_metadata_fwd__18_, fe_pc_gen_branch_metadata_fwd__17_, fe_pc_gen_branch_metadata_fwd__16_, fe_pc_gen_branch_metadata_fwd__15_, fe_pc_gen_branch_metadata_fwd__14_, fe_pc_gen_branch_metadata_fwd__13_, fe_pc_gen_branch_metadata_fwd__12_, fe_pc_gen_branch_metadata_fwd__11_, fe_pc_gen_branch_metadata_fwd__10_, fe_pc_gen_branch_metadata_fwd__9_, fe_pc_gen_branch_metadata_fwd__8_, fe_pc_gen_branch_metadata_fwd__7_, fe_pc_gen_branch_metadata_fwd__6_, fe_pc_gen_branch_metadata_fwd__5_, fe_pc_gen_branch_metadata_fwd__4_, fe_pc_gen_branch_metadata_fwd__3_, fe_pc_gen_branch_metadata_fwd__2_, fe_pc_gen_branch_metadata_fwd__1_, fe_pc_gen_branch_metadata_fwd__0_, N11, fe_pc_gen_pc_redirect_valid_, N27, N35, N15, N18 }),
    .fe_pc_gen_v_i(fe_cmd_v_i),
    .fe_pc_gen_ready_o(fe_cmd_ready_o),
    .itlb_miss_i(itlb_miss)
  );


  bp_fe_icache_02
  icache
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .freeze_i(freeze_i),
    .id_i(icache_id_i[0]),
    .cfg_w_v_i(cfg_w_v_i),
    .cfg_addr_i(cfg_addr_i),
    .cfg_data_i(cfg_data_i),
    .pc_gen_icache_vaddr_i(pc_gen_icache),
    .pc_gen_icache_vaddr_v_i(pc_gen_icache_v),
    .pc_gen_icache_vaddr_ready_o(pc_gen_icache_ready),
    .icache_pc_gen_data_o(icache_pc_gen),
    .icache_pc_gen_data_v_o(icache_pc_gen_v),
    .icache_pc_gen_data_ready_i(icache_pc_gen_ready),
    .itlb_icache_data_resp_i(itlb_icache),
    .itlb_icache_data_resp_v_i(itlb_icache_data_resp_v),
    .itlb_icache_data_resp_ready_o(itlb_icache_data_resp_ready),
    .itlb_icache_miss_i(itlb_miss),
    .uncached_i(itlb_entry_r_uc_),
    .cache_miss_o(icache_miss),
    .instr_access_fault_o(instr_access_fault),
    .poison_tl_i(poison_tl),
    .lce_req_o(lce_req_o),
    .lce_req_v_o(lce_req_v_o),
    .lce_req_ready_i(lce_req_ready_i),
    .lce_resp_o(lce_resp_o),
    .lce_resp_v_o(lce_resp_v_o),
    .lce_resp_ready_i(lce_resp_ready_i),
    .lce_data_resp_o(lce_data_resp_o),
    .lce_data_resp_v_o(lce_data_resp_v_o),
    .lce_data_resp_ready_i(lce_data_resp_ready_i),
    .lce_cmd_i(lce_cmd_i),
    .lce_cmd_v_i(lce_cmd_v_i),
    .lce_cmd_ready_o(lce_cmd_ready_o),
    .lce_data_cmd_i(lce_data_cmd_i),
    .lce_data_cmd_v_i(lce_data_cmd_v_i),
    .lce_data_cmd_ready_o(lce_data_cmd_ready_o),
    .lce_data_cmd_o(lce_data_cmd_o),
    .lce_data_cmd_v_o(lce_data_cmd_v_o),
    .lce_data_cmd_ready_i(lce_data_cmd_ready_i)
  );


  bp_be_dtlb_02
  itlb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .flush_i(itlb_fence_v),
    .r_v_i(pc_gen_itlb_v),
    .r_ready_o(pc_gen_itlb_ready),
    .r_vtag_i(itlb_vaddr[38:12]),
    .r_v_o(itlb_icache_data_resp_v),
    .r_entry_o({ itlb_icache, itlb_entry_r_g_, itlb_entry_r_u_, itlb_entry_r_x_, itlb_entry_r_w_, itlb_entry_r_r_, itlb_entry_r_uc_ }),
    .w_v_i(itlb_w_v),
    .w_vtag_i(fe_cmd_i[72:46]),
    .w_entry_i(fe_cmd_i[33:1]),
    .miss_v_o(itlb_miss),
    .miss_vtag_o(itlb_miss_vtag)
  );

  assign N9 = fe_cmd_i[74] | fe_cmd_i[75];
  assign N10 = fe_cmd_i[73] | N9;
  assign N11 = ~N10;
  assign N12 = ~fe_cmd_i[74];
  assign N13 = N12 | fe_cmd_i[75];
  assign N14 = N32 | N13;
  assign N15 = ~N14;
  assign N16 = N12 | N31;
  assign N17 = fe_cmd_i[73] | N16;
  assign N18 = ~N17;
  assign N19 = fe_cmd_i[74] | fe_cmd_i[75];
  assign N20 = N32 | N19;
  assign N21 = ~N20;
  assign N22 = ~fe_cmd_i[33];
  assign N23 = fe_cmd_i[32] | N22;
  assign N24 = fe_cmd_i[31] | N23;
  assign N25 = ~N24;
  assign N26 = fe_cmd_i[73] | N33;
  assign N27 = ~N26;
  assign N28 = N12 | N31;
  assign N29 = fe_cmd_i[73] | N28;
  assign N30 = ~N29;
  assign N31 = ~fe_cmd_i[75];
  assign N32 = ~fe_cmd_i[73];
  assign N33 = fe_cmd_i[74] | N31;
  assign N34 = N32 | N33;
  assign N35 = ~N34;
  assign N36 = fe_cmd_i[74] | fe_cmd_i[75];
  assign N37 = N32 | N36;
  assign N38 = ~N37;
  assign N39 = fe_cmd_i[73] | N33;
  assign N40 = ~N39;
  assign { fe_pc_gen_branch_metadata_fwd__26_, fe_pc_gen_branch_metadata_fwd__25_, fe_pc_gen_branch_metadata_fwd__24_, fe_pc_gen_branch_metadata_fwd__23_, fe_pc_gen_branch_metadata_fwd__22_, fe_pc_gen_branch_metadata_fwd__21_, fe_pc_gen_branch_metadata_fwd__20_, fe_pc_gen_branch_metadata_fwd__19_, fe_pc_gen_branch_metadata_fwd__18_, fe_pc_gen_branch_metadata_fwd__17_, fe_pc_gen_branch_metadata_fwd__16_, fe_pc_gen_branch_metadata_fwd__15_, fe_pc_gen_branch_metadata_fwd__14_, fe_pc_gen_branch_metadata_fwd__13_, fe_pc_gen_branch_metadata_fwd__12_, fe_pc_gen_branch_metadata_fwd__11_, fe_pc_gen_branch_metadata_fwd__10_, fe_pc_gen_branch_metadata_fwd__9_, fe_pc_gen_branch_metadata_fwd__8_, fe_pc_gen_branch_metadata_fwd__7_, fe_pc_gen_branch_metadata_fwd__6_, fe_pc_gen_branch_metadata_fwd__5_, fe_pc_gen_branch_metadata_fwd__4_, fe_pc_gen_branch_metadata_fwd__3_, fe_pc_gen_branch_metadata_fwd__2_, fe_pc_gen_branch_metadata_fwd__1_, fe_pc_gen_branch_metadata_fwd__0_ } = (N0)? fe_cmd_i[33:7] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                (N1)? fe_cmd_i[30:4] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N0 = N40;
  assign N1 = N38;
  assign N8 = (N2)? 1'b0 : 
              (N3)? itlb_fill_v : 1'b0;
  assign N2 = N7;
  assign N3 = N6;
  assign fe_pc_gen_pc_redirect_valid_ = N21 & N25;
  assign N4 = N38 | N40;
  assign N5 = ~N4;
  assign poison_tl = icache_miss | N42;
  assign N42 = fe_cmd_v_i & N41;
  assign N41 = ~N27;
  assign itlb_fill_v = fe_cmd_v_i & N35;
  assign itlb_w_v = itlb_fill_v & N43;
  assign N43 = ~itlb_fill_r;
  assign itlb_fence_v = fe_cmd_v_i & N30;
  assign N6 = ~reset_i;
  assign N7 = reset_i;

  always @(posedge clk_i) begin
    if(1'b1) begin
      itlb_fill_r <= N8;
    end 
  end


endmodule
