BUSBITCHARS "[]" ;

MACRO nangate45_8x64_1P_bit
  FOREIGN nangate45_8x64_1P_bit 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 100.0 BY 100.0 ;
  CLASS RING ;
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 8.5 89.79 9.0 90.0 ;
      LAYER metal2 ;
      RECT 8.5 89.79 9.0 90.0 ;
      LAYER metal3 ;
      RECT 8.5 89.79 9.0 90.0 ;
      LAYER metal4 ;
      RECT 8.5 89.79 9.0 90.0 ;
      END
    END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 8.5 86.3117391304 9.0 86.5217391304 ;
      LAYER metal2 ;
      RECT 8.5 86.3117391304 9.0 86.5217391304 ;
      LAYER metal3 ;
      RECT 8.5 86.3117391304 9.0 86.5217391304 ;
      LAYER metal4 ;
      RECT 8.5 86.3117391304 9.0 86.5217391304 ;
      END
    END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 8.5 82.8334782609 9.0 83.0434782609 ;
      LAYER metal2 ;
      RECT 8.5 82.8334782609 9.0 83.0434782609 ;
      LAYER metal3 ;
      RECT 8.5 82.8334782609 9.0 83.0434782609 ;
      LAYER metal4 ;
      RECT 8.5 82.8334782609 9.0 83.0434782609 ;
      END
    END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 8.5 79.3552173913 9.0 79.5652173913 ;
      LAYER metal2 ;
      RECT 8.5 79.3552173913 9.0 79.5652173913 ;
      LAYER metal3 ;
      RECT 8.5 79.3552173913 9.0 79.5652173913 ;
      LAYER metal4 ;
      RECT 8.5 79.3552173913 9.0 79.5652173913 ;
      END
    END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 8.5 75.8769565217 9.0 76.0869565217 ;
      LAYER metal2 ;
      RECT 8.5 75.8769565217 9.0 76.0869565217 ;
      LAYER metal3 ;
      RECT 8.5 75.8769565217 9.0 76.0869565217 ;
      LAYER metal4 ;
      RECT 8.5 75.8769565217 9.0 76.0869565217 ;
      END
    END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 8.5 72.3986956522 9.0 72.6086956522 ;
      LAYER metal2 ;
      RECT 8.5 72.3986956522 9.0 72.6086956522 ;
      LAYER metal3 ;
      RECT 8.5 72.3986956522 9.0 72.6086956522 ;
      LAYER metal4 ;
      RECT 8.5 72.3986956522 9.0 72.6086956522 ;
      END
    END addr_in[5]
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 8.5 68.9204347826 9.0 69.1304347826 ;
      LAYER metal2 ;
      RECT 8.5 68.9204347826 9.0 69.1304347826 ;
      LAYER metal3 ;
      RECT 8.5 68.9204347826 9.0 69.1304347826 ;
      LAYER metal4 ;
      RECT 8.5 68.9204347826 9.0 69.1304347826 ;
      END
    END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 8.5 65.442173913 9.0 65.652173913 ;
      LAYER metal2 ;
      RECT 8.5 65.442173913 9.0 65.652173913 ;
      LAYER metal3 ;
      RECT 8.5 65.442173913 9.0 65.652173913 ;
      LAYER metal4 ;
      RECT 8.5 65.442173913 9.0 65.652173913 ;
      END
    END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 8.5 61.9639130435 9.0 62.1739130435 ;
      LAYER metal2 ;
      RECT 8.5 61.9639130435 9.0 62.1739130435 ;
      LAYER metal3 ;
      RECT 8.5 61.9639130435 9.0 62.1739130435 ;
      LAYER metal4 ;
      RECT 8.5 61.9639130435 9.0 62.1739130435 ;
      END
    END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 8.5 58.4856521739 9.0 58.6956521739 ;
      LAYER metal2 ;
      RECT 8.5 58.4856521739 9.0 58.6956521739 ;
      LAYER metal3 ;
      RECT 8.5 58.4856521739 9.0 58.6956521739 ;
      LAYER metal4 ;
      RECT 8.5 58.4856521739 9.0 58.6956521739 ;
      END
    END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 8.5 55.0073913043 9.0 55.2173913043 ;
      LAYER metal2 ;
      RECT 8.5 55.0073913043 9.0 55.2173913043 ;
      LAYER metal3 ;
      RECT 8.5 55.0073913043 9.0 55.2173913043 ;
      LAYER metal4 ;
      RECT 8.5 55.0073913043 9.0 55.2173913043 ;
      END
    END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 8.5 51.5291304348 9.0 51.7391304348 ;
      LAYER metal2 ;
      RECT 8.5 51.5291304348 9.0 51.7391304348 ;
      LAYER metal3 ;
      RECT 8.5 51.5291304348 9.0 51.7391304348 ;
      LAYER metal4 ;
      RECT 8.5 51.5291304348 9.0 51.7391304348 ;
      END
    END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 8.5 48.0508695652 9.0 48.2608695652 ;
      LAYER metal2 ;
      RECT 8.5 48.0508695652 9.0 48.2608695652 ;
      LAYER metal3 ;
      RECT 8.5 48.0508695652 9.0 48.2608695652 ;
      LAYER metal4 ;
      RECT 8.5 48.0508695652 9.0 48.2608695652 ;
      END
    END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 8.5 44.5726086957 9.0 44.7826086957 ;
      LAYER metal2 ;
      RECT 8.5 44.5726086957 9.0 44.7826086957 ;
      LAYER metal3 ;
      RECT 8.5 44.5726086957 9.0 44.7826086957 ;
      LAYER metal4 ;
      RECT 8.5 44.5726086957 9.0 44.7826086957 ;
      END
    END w_mask_in[7]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 8.5 41.0943478261 9.0 41.3043478261 ;
      LAYER metal2 ;
      RECT 8.5 41.0943478261 9.0 41.3043478261 ;
      LAYER metal3 ;
      RECT 8.5 41.0943478261 9.0 41.3043478261 ;
      LAYER metal4 ;
      RECT 8.5 41.0943478261 9.0 41.3043478261 ;
      END
    END we_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 8.5 37.6160869565 9.0 37.8260869565 ;
      LAYER metal2 ;
      RECT 8.5 37.6160869565 9.0 37.8260869565 ;
      LAYER metal3 ;
      RECT 8.5 37.6160869565 9.0 37.8260869565 ;
      LAYER metal4 ;
      RECT 8.5 37.6160869565 9.0 37.8260869565 ;
      END
    END clk
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 8.5 34.137826087 9.0 34.347826087 ;
      LAYER metal2 ;
      RECT 8.5 34.137826087 9.0 34.347826087 ;
      LAYER metal3 ;
      RECT 8.5 34.137826087 9.0 34.347826087 ;
      LAYER metal4 ;
      RECT 8.5 34.137826087 9.0 34.347826087 ;
      END
    END ce_in
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 89.5 59.79 90.0 60.0 ;
      LAYER metal2 ;
      RECT 89.5 59.79 90.0 60.0 ;
      LAYER metal3 ;
      RECT 89.5 59.79 90.0 60.0 ;
      LAYER metal4 ;
      RECT 89.5 59.79 90.0 60.0 ;
      END
    END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 80.125 59.79 80.625 60.0 ;
      LAYER metal2 ;
      RECT 80.125 59.79 80.625 60.0 ;
      LAYER metal3 ;
      RECT 80.125 59.79 80.625 60.0 ;
      LAYER metal4 ;
      RECT 80.125 59.79 80.625 60.0 ;
      END
    END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 70.75 59.79 71.25 60.0 ;
      LAYER metal2 ;
      RECT 70.75 59.79 71.25 60.0 ;
      LAYER metal3 ;
      RECT 70.75 59.79 71.25 60.0 ;
      LAYER metal4 ;
      RECT 70.75 59.79 71.25 60.0 ;
      END
    END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 61.375 59.79 61.875 60.0 ;
      LAYER metal2 ;
      RECT 61.375 59.79 61.875 60.0 ;
      LAYER metal3 ;
      RECT 61.375 59.79 61.875 60.0 ;
      LAYER metal4 ;
      RECT 61.375 59.79 61.875 60.0 ;
      END
    END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 52.0 59.79 52.5 60.0 ;
      LAYER metal2 ;
      RECT 52.0 59.79 52.5 60.0 ;
      LAYER metal3 ;
      RECT 52.0 59.79 52.5 60.0 ;
      LAYER metal4 ;
      RECT 52.0 59.79 52.5 60.0 ;
      END
    END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 42.625 59.79 43.125 60.0 ;
      LAYER metal2 ;
      RECT 42.625 59.79 43.125 60.0 ;
      LAYER metal3 ;
      RECT 42.625 59.79 43.125 60.0 ;
      LAYER metal4 ;
      RECT 42.625 59.79 43.125 60.0 ;
      END
    END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 33.25 59.79 33.75 60.0 ;
      LAYER metal2 ;
      RECT 33.25 59.79 33.75 60.0 ;
      LAYER metal3 ;
      RECT 33.25 59.79 33.75 60.0 ;
      LAYER metal4 ;
      RECT 33.25 59.79 33.75 60.0 ;
      END
    END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 23.875 59.79 24.375 60.0 ;
      LAYER metal2 ;
      RECT 23.875 59.79 24.375 60.0 ;
      LAYER metal3 ;
      RECT 23.875 59.79 24.375 60.0 ;
      LAYER metal4 ;
      RECT 23.875 59.79 24.375 60.0 ;
      END
    END rd_out[7]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 89.5 39.79 90.0 40.0 ;
      LAYER metal2 ;
      RECT 89.5 39.79 90.0 40.0 ;
      LAYER metal3 ;
      RECT 89.5 39.79 90.0 40.0 ;
      LAYER metal4 ;
      RECT 89.5 39.79 90.0 40.0 ;
      END
    END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 80.125 39.79 80.625 40.0 ;
      LAYER metal2 ;
      RECT 80.125 39.79 80.625 40.0 ;
      LAYER metal3 ;
      RECT 80.125 39.79 80.625 40.0 ;
      LAYER metal4 ;
      RECT 80.125 39.79 80.625 40.0 ;
      END
    END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 70.75 39.79 71.25 40.0 ;
      LAYER metal2 ;
      RECT 70.75 39.79 71.25 40.0 ;
      LAYER metal3 ;
      RECT 70.75 39.79 71.25 40.0 ;
      LAYER metal4 ;
      RECT 70.75 39.79 71.25 40.0 ;
      END
    END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 61.375 39.79 61.875 40.0 ;
      LAYER metal2 ;
      RECT 61.375 39.79 61.875 40.0 ;
      LAYER metal3 ;
      RECT 61.375 39.79 61.875 40.0 ;
      LAYER metal4 ;
      RECT 61.375 39.79 61.875 40.0 ;
      END
    END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 52.0 39.79 52.5 40.0 ;
      LAYER metal2 ;
      RECT 52.0 39.79 52.5 40.0 ;
      LAYER metal3 ;
      RECT 52.0 39.79 52.5 40.0 ;
      LAYER metal4 ;
      RECT 52.0 39.79 52.5 40.0 ;
      END
    END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 42.625 39.79 43.125 40.0 ;
      LAYER metal2 ;
      RECT 42.625 39.79 43.125 40.0 ;
      LAYER metal3 ;
      RECT 42.625 39.79 43.125 40.0 ;
      LAYER metal4 ;
      RECT 42.625 39.79 43.125 40.0 ;
      END
    END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 33.25 39.79 33.75 40.0 ;
      LAYER metal2 ;
      RECT 33.25 39.79 33.75 40.0 ;
      LAYER metal3 ;
      RECT 33.25 39.79 33.75 40.0 ;
      LAYER metal4 ;
      RECT 33.25 39.79 33.75 40.0 ;
      END
    END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 23.875 39.79 24.375 40.0 ;
      LAYER metal2 ;
      RECT 23.875 39.79 24.375 40.0 ;
      LAYER metal3 ;
      RECT 23.875 39.79 24.375 40.0 ;
      LAYER metal4 ;
      RECT 23.875 39.79 24.375 40.0 ;
      END
    END wd_in[7]
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE RING ;
    PORT
      LAYER metal3 ;
      RECT 3.5 3.5 5.5 96.5 ;
      END
    PORT
      LAYER metal4 ;
      RECT 3.5 3.5 5.5 96.5 ;
      END
    END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE RING ;
    PORT
      LAYER metal3 ;
      RECT 0.0 0.0 98.0 2.0 ;
      END
    PORT
      LAYER metal4 ;
      RECT 0.0 0.0 98.0 2.0 ;
      END
    END VDD
  OBS
    #core
    LAYER VIA1 ;
    RECT 8.5 8.5 91.5 91.5 ;
    LAYER VIA2 ;
    RECT 8.5 8.5 91.5 91.5 ;
    LAYER VIA3 ;
    RECT 8.5 8.5 91.5 91.5 ;
    LAYER OVERLAP ;
    RECT 8.5 8.5 91.5 91.5 ;
    END
  END nangate45_8x64_1P_bit

END LIBRARY
