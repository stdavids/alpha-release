BUSBITCHARS "[]" ;

MACRO nangate45_64x512_1P_BM
  FOREIGN nangate45_64x512_1P_BM 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 100.0 BY 100.0 ;
  CLASS RING ;
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 89.79 9.0 90.0 ;
      LAYER M2 ;
      RECT 8.5 89.79 9.0 90.0 ;
      LAYER M3 ;
      RECT 8.5 89.79 9.0 90.0 ;
      LAYER M4 ;
      RECT 8.5 89.79 9.0 90.0 ;
      END
    END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 88.8488235294 9.0 89.0588235294 ;
      LAYER M2 ;
      RECT 8.5 88.8488235294 9.0 89.0588235294 ;
      LAYER M3 ;
      RECT 8.5 88.8488235294 9.0 89.0588235294 ;
      LAYER M4 ;
      RECT 8.5 88.8488235294 9.0 89.0588235294 ;
      END
    END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 87.9076470588 9.0 88.1176470588 ;
      LAYER M2 ;
      RECT 8.5 87.9076470588 9.0 88.1176470588 ;
      LAYER M3 ;
      RECT 8.5 87.9076470588 9.0 88.1176470588 ;
      LAYER M4 ;
      RECT 8.5 87.9076470588 9.0 88.1176470588 ;
      END
    END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 86.9664705882 9.0 87.1764705882 ;
      LAYER M2 ;
      RECT 8.5 86.9664705882 9.0 87.1764705882 ;
      LAYER M3 ;
      RECT 8.5 86.9664705882 9.0 87.1764705882 ;
      LAYER M4 ;
      RECT 8.5 86.9664705882 9.0 87.1764705882 ;
      END
    END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 86.0252941176 9.0 86.2352941176 ;
      LAYER M2 ;
      RECT 8.5 86.0252941176 9.0 86.2352941176 ;
      LAYER M3 ;
      RECT 8.5 86.0252941176 9.0 86.2352941176 ;
      LAYER M4 ;
      RECT 8.5 86.0252941176 9.0 86.2352941176 ;
      END
    END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 85.0841176471 9.0 85.2941176471 ;
      LAYER M2 ;
      RECT 8.5 85.0841176471 9.0 85.2941176471 ;
      LAYER M3 ;
      RECT 8.5 85.0841176471 9.0 85.2941176471 ;
      LAYER M4 ;
      RECT 8.5 85.0841176471 9.0 85.2941176471 ;
      END
    END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 84.1429411765 9.0 84.3529411765 ;
      LAYER M2 ;
      RECT 8.5 84.1429411765 9.0 84.3529411765 ;
      LAYER M3 ;
      RECT 8.5 84.1429411765 9.0 84.3529411765 ;
      LAYER M4 ;
      RECT 8.5 84.1429411765 9.0 84.3529411765 ;
      END
    END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 83.2017647059 9.0 83.4117647059 ;
      LAYER M2 ;
      RECT 8.5 83.2017647059 9.0 83.4117647059 ;
      LAYER M3 ;
      RECT 8.5 83.2017647059 9.0 83.4117647059 ;
      LAYER M4 ;
      RECT 8.5 83.2017647059 9.0 83.4117647059 ;
      END
    END addr_in[7]
  PIN addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 82.2605882353 9.0 82.4705882353 ;
      LAYER M2 ;
      RECT 8.5 82.2605882353 9.0 82.4705882353 ;
      LAYER M3 ;
      RECT 8.5 82.2605882353 9.0 82.4705882353 ;
      LAYER M4 ;
      RECT 8.5 82.2605882353 9.0 82.4705882353 ;
      END
    END addr_in[8]
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 81.3194117647 9.0 81.5294117647 ;
      LAYER M2 ;
      RECT 8.5 81.3194117647 9.0 81.5294117647 ;
      LAYER M3 ;
      RECT 8.5 81.3194117647 9.0 81.5294117647 ;
      LAYER M4 ;
      RECT 8.5 81.3194117647 9.0 81.5294117647 ;
      END
    END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 80.3782352941 9.0 80.5882352941 ;
      LAYER M2 ;
      RECT 8.5 80.3782352941 9.0 80.5882352941 ;
      LAYER M3 ;
      RECT 8.5 80.3782352941 9.0 80.5882352941 ;
      LAYER M4 ;
      RECT 8.5 80.3782352941 9.0 80.5882352941 ;
      END
    END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 79.4370588235 9.0 79.6470588235 ;
      LAYER M2 ;
      RECT 8.5 79.4370588235 9.0 79.6470588235 ;
      LAYER M3 ;
      RECT 8.5 79.4370588235 9.0 79.6470588235 ;
      LAYER M4 ;
      RECT 8.5 79.4370588235 9.0 79.6470588235 ;
      END
    END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 78.4958823529 9.0 78.7058823529 ;
      LAYER M2 ;
      RECT 8.5 78.4958823529 9.0 78.7058823529 ;
      LAYER M3 ;
      RECT 8.5 78.4958823529 9.0 78.7058823529 ;
      LAYER M4 ;
      RECT 8.5 78.4958823529 9.0 78.7058823529 ;
      END
    END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 77.5547058824 9.0 77.7647058824 ;
      LAYER M2 ;
      RECT 8.5 77.5547058824 9.0 77.7647058824 ;
      LAYER M3 ;
      RECT 8.5 77.5547058824 9.0 77.7647058824 ;
      LAYER M4 ;
      RECT 8.5 77.5547058824 9.0 77.7647058824 ;
      END
    END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 76.6135294118 9.0 76.8235294118 ;
      LAYER M2 ;
      RECT 8.5 76.6135294118 9.0 76.8235294118 ;
      LAYER M3 ;
      RECT 8.5 76.6135294118 9.0 76.8235294118 ;
      LAYER M4 ;
      RECT 8.5 76.6135294118 9.0 76.8235294118 ;
      END
    END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 75.6723529412 9.0 75.8823529412 ;
      LAYER M2 ;
      RECT 8.5 75.6723529412 9.0 75.8823529412 ;
      LAYER M3 ;
      RECT 8.5 75.6723529412 9.0 75.8823529412 ;
      LAYER M4 ;
      RECT 8.5 75.6723529412 9.0 75.8823529412 ;
      END
    END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 74.7311764706 9.0 74.9411764706 ;
      LAYER M2 ;
      RECT 8.5 74.7311764706 9.0 74.9411764706 ;
      LAYER M3 ;
      RECT 8.5 74.7311764706 9.0 74.9411764706 ;
      LAYER M4 ;
      RECT 8.5 74.7311764706 9.0 74.9411764706 ;
      END
    END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 73.79 9.0 74.0 ;
      LAYER M2 ;
      RECT 8.5 73.79 9.0 74.0 ;
      LAYER M3 ;
      RECT 8.5 73.79 9.0 74.0 ;
      LAYER M4 ;
      RECT 8.5 73.79 9.0 74.0 ;
      END
    END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 72.8488235294 9.0 73.0588235294 ;
      LAYER M2 ;
      RECT 8.5 72.8488235294 9.0 73.0588235294 ;
      LAYER M3 ;
      RECT 8.5 72.8488235294 9.0 73.0588235294 ;
      LAYER M4 ;
      RECT 8.5 72.8488235294 9.0 73.0588235294 ;
      END
    END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 71.9076470588 9.0 72.1176470588 ;
      LAYER M2 ;
      RECT 8.5 71.9076470588 9.0 72.1176470588 ;
      LAYER M3 ;
      RECT 8.5 71.9076470588 9.0 72.1176470588 ;
      LAYER M4 ;
      RECT 8.5 71.9076470588 9.0 72.1176470588 ;
      END
    END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 70.9664705882 9.0 71.1764705882 ;
      LAYER M2 ;
      RECT 8.5 70.9664705882 9.0 71.1764705882 ;
      LAYER M3 ;
      RECT 8.5 70.9664705882 9.0 71.1764705882 ;
      LAYER M4 ;
      RECT 8.5 70.9664705882 9.0 71.1764705882 ;
      END
    END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 70.0252941176 9.0 70.2352941176 ;
      LAYER M2 ;
      RECT 8.5 70.0252941176 9.0 70.2352941176 ;
      LAYER M3 ;
      RECT 8.5 70.0252941176 9.0 70.2352941176 ;
      LAYER M4 ;
      RECT 8.5 70.0252941176 9.0 70.2352941176 ;
      END
    END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 69.0841176471 9.0 69.2941176471 ;
      LAYER M2 ;
      RECT 8.5 69.0841176471 9.0 69.2941176471 ;
      LAYER M3 ;
      RECT 8.5 69.0841176471 9.0 69.2941176471 ;
      LAYER M4 ;
      RECT 8.5 69.0841176471 9.0 69.2941176471 ;
      END
    END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 68.1429411765 9.0 68.3529411765 ;
      LAYER M2 ;
      RECT 8.5 68.1429411765 9.0 68.3529411765 ;
      LAYER M3 ;
      RECT 8.5 68.1429411765 9.0 68.3529411765 ;
      LAYER M4 ;
      RECT 8.5 68.1429411765 9.0 68.3529411765 ;
      END
    END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 67.2017647059 9.0 67.4117647059 ;
      LAYER M2 ;
      RECT 8.5 67.2017647059 9.0 67.4117647059 ;
      LAYER M3 ;
      RECT 8.5 67.2017647059 9.0 67.4117647059 ;
      LAYER M4 ;
      RECT 8.5 67.2017647059 9.0 67.4117647059 ;
      END
    END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 66.2605882353 9.0 66.4705882353 ;
      LAYER M2 ;
      RECT 8.5 66.2605882353 9.0 66.4705882353 ;
      LAYER M3 ;
      RECT 8.5 66.2605882353 9.0 66.4705882353 ;
      LAYER M4 ;
      RECT 8.5 66.2605882353 9.0 66.4705882353 ;
      END
    END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 65.3194117647 9.0 65.5294117647 ;
      LAYER M2 ;
      RECT 8.5 65.3194117647 9.0 65.5294117647 ;
      LAYER M3 ;
      RECT 8.5 65.3194117647 9.0 65.5294117647 ;
      LAYER M4 ;
      RECT 8.5 65.3194117647 9.0 65.5294117647 ;
      END
    END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 64.3782352941 9.0 64.5882352941 ;
      LAYER M2 ;
      RECT 8.5 64.3782352941 9.0 64.5882352941 ;
      LAYER M3 ;
      RECT 8.5 64.3782352941 9.0 64.5882352941 ;
      LAYER M4 ;
      RECT 8.5 64.3782352941 9.0 64.5882352941 ;
      END
    END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 63.4370588235 9.0 63.6470588235 ;
      LAYER M2 ;
      RECT 8.5 63.4370588235 9.0 63.6470588235 ;
      LAYER M3 ;
      RECT 8.5 63.4370588235 9.0 63.6470588235 ;
      LAYER M4 ;
      RECT 8.5 63.4370588235 9.0 63.6470588235 ;
      END
    END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 62.4958823529 9.0 62.7058823529 ;
      LAYER M2 ;
      RECT 8.5 62.4958823529 9.0 62.7058823529 ;
      LAYER M3 ;
      RECT 8.5 62.4958823529 9.0 62.7058823529 ;
      LAYER M4 ;
      RECT 8.5 62.4958823529 9.0 62.7058823529 ;
      END
    END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 61.5547058824 9.0 61.7647058824 ;
      LAYER M2 ;
      RECT 8.5 61.5547058824 9.0 61.7647058824 ;
      LAYER M3 ;
      RECT 8.5 61.5547058824 9.0 61.7647058824 ;
      LAYER M4 ;
      RECT 8.5 61.5547058824 9.0 61.7647058824 ;
      END
    END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 60.6135294118 9.0 60.8235294118 ;
      LAYER M2 ;
      RECT 8.5 60.6135294118 9.0 60.8235294118 ;
      LAYER M3 ;
      RECT 8.5 60.6135294118 9.0 60.8235294118 ;
      LAYER M4 ;
      RECT 8.5 60.6135294118 9.0 60.8235294118 ;
      END
    END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 59.6723529412 9.0 59.8823529412 ;
      LAYER M2 ;
      RECT 8.5 59.6723529412 9.0 59.8823529412 ;
      LAYER M3 ;
      RECT 8.5 59.6723529412 9.0 59.8823529412 ;
      LAYER M4 ;
      RECT 8.5 59.6723529412 9.0 59.8823529412 ;
      END
    END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 58.7311764706 9.0 58.9411764706 ;
      LAYER M2 ;
      RECT 8.5 58.7311764706 9.0 58.9411764706 ;
      LAYER M3 ;
      RECT 8.5 58.7311764706 9.0 58.9411764706 ;
      LAYER M4 ;
      RECT 8.5 58.7311764706 9.0 58.9411764706 ;
      END
    END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 57.79 9.0 58.0 ;
      LAYER M2 ;
      RECT 8.5 57.79 9.0 58.0 ;
      LAYER M3 ;
      RECT 8.5 57.79 9.0 58.0 ;
      LAYER M4 ;
      RECT 8.5 57.79 9.0 58.0 ;
      END
    END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 56.8488235294 9.0 57.0588235294 ;
      LAYER M2 ;
      RECT 8.5 56.8488235294 9.0 57.0588235294 ;
      LAYER M3 ;
      RECT 8.5 56.8488235294 9.0 57.0588235294 ;
      LAYER M4 ;
      RECT 8.5 56.8488235294 9.0 57.0588235294 ;
      END
    END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 55.9076470588 9.0 56.1176470588 ;
      LAYER M2 ;
      RECT 8.5 55.9076470588 9.0 56.1176470588 ;
      LAYER M3 ;
      RECT 8.5 55.9076470588 9.0 56.1176470588 ;
      LAYER M4 ;
      RECT 8.5 55.9076470588 9.0 56.1176470588 ;
      END
    END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 54.9664705882 9.0 55.1764705882 ;
      LAYER M2 ;
      RECT 8.5 54.9664705882 9.0 55.1764705882 ;
      LAYER M3 ;
      RECT 8.5 54.9664705882 9.0 55.1764705882 ;
      LAYER M4 ;
      RECT 8.5 54.9664705882 9.0 55.1764705882 ;
      END
    END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 54.0252941176 9.0 54.2352941176 ;
      LAYER M2 ;
      RECT 8.5 54.0252941176 9.0 54.2352941176 ;
      LAYER M3 ;
      RECT 8.5 54.0252941176 9.0 54.2352941176 ;
      LAYER M4 ;
      RECT 8.5 54.0252941176 9.0 54.2352941176 ;
      END
    END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 53.0841176471 9.0 53.2941176471 ;
      LAYER M2 ;
      RECT 8.5 53.0841176471 9.0 53.2941176471 ;
      LAYER M3 ;
      RECT 8.5 53.0841176471 9.0 53.2941176471 ;
      LAYER M4 ;
      RECT 8.5 53.0841176471 9.0 53.2941176471 ;
      END
    END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 52.1429411765 9.0 52.3529411765 ;
      LAYER M2 ;
      RECT 8.5 52.1429411765 9.0 52.3529411765 ;
      LAYER M3 ;
      RECT 8.5 52.1429411765 9.0 52.3529411765 ;
      LAYER M4 ;
      RECT 8.5 52.1429411765 9.0 52.3529411765 ;
      END
    END w_mask_in[31]
  PIN w_mask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 51.2017647059 9.0 51.4117647059 ;
      LAYER M2 ;
      RECT 8.5 51.2017647059 9.0 51.4117647059 ;
      LAYER M3 ;
      RECT 8.5 51.2017647059 9.0 51.4117647059 ;
      LAYER M4 ;
      RECT 8.5 51.2017647059 9.0 51.4117647059 ;
      END
    END w_mask_in[32]
  PIN w_mask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 50.2605882353 9.0 50.4705882353 ;
      LAYER M2 ;
      RECT 8.5 50.2605882353 9.0 50.4705882353 ;
      LAYER M3 ;
      RECT 8.5 50.2605882353 9.0 50.4705882353 ;
      LAYER M4 ;
      RECT 8.5 50.2605882353 9.0 50.4705882353 ;
      END
    END w_mask_in[33]
  PIN w_mask_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 49.3194117647 9.0 49.5294117647 ;
      LAYER M2 ;
      RECT 8.5 49.3194117647 9.0 49.5294117647 ;
      LAYER M3 ;
      RECT 8.5 49.3194117647 9.0 49.5294117647 ;
      LAYER M4 ;
      RECT 8.5 49.3194117647 9.0 49.5294117647 ;
      END
    END w_mask_in[34]
  PIN w_mask_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 48.3782352941 9.0 48.5882352941 ;
      LAYER M2 ;
      RECT 8.5 48.3782352941 9.0 48.5882352941 ;
      LAYER M3 ;
      RECT 8.5 48.3782352941 9.0 48.5882352941 ;
      LAYER M4 ;
      RECT 8.5 48.3782352941 9.0 48.5882352941 ;
      END
    END w_mask_in[35]
  PIN w_mask_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 47.4370588235 9.0 47.6470588235 ;
      LAYER M2 ;
      RECT 8.5 47.4370588235 9.0 47.6470588235 ;
      LAYER M3 ;
      RECT 8.5 47.4370588235 9.0 47.6470588235 ;
      LAYER M4 ;
      RECT 8.5 47.4370588235 9.0 47.6470588235 ;
      END
    END w_mask_in[36]
  PIN w_mask_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 46.4958823529 9.0 46.7058823529 ;
      LAYER M2 ;
      RECT 8.5 46.4958823529 9.0 46.7058823529 ;
      LAYER M3 ;
      RECT 8.5 46.4958823529 9.0 46.7058823529 ;
      LAYER M4 ;
      RECT 8.5 46.4958823529 9.0 46.7058823529 ;
      END
    END w_mask_in[37]
  PIN w_mask_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 45.5547058824 9.0 45.7647058824 ;
      LAYER M2 ;
      RECT 8.5 45.5547058824 9.0 45.7647058824 ;
      LAYER M3 ;
      RECT 8.5 45.5547058824 9.0 45.7647058824 ;
      LAYER M4 ;
      RECT 8.5 45.5547058824 9.0 45.7647058824 ;
      END
    END w_mask_in[38]
  PIN w_mask_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 44.6135294118 9.0 44.8235294118 ;
      LAYER M2 ;
      RECT 8.5 44.6135294118 9.0 44.8235294118 ;
      LAYER M3 ;
      RECT 8.5 44.6135294118 9.0 44.8235294118 ;
      LAYER M4 ;
      RECT 8.5 44.6135294118 9.0 44.8235294118 ;
      END
    END w_mask_in[39]
  PIN w_mask_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 43.6723529412 9.0 43.8823529412 ;
      LAYER M2 ;
      RECT 8.5 43.6723529412 9.0 43.8823529412 ;
      LAYER M3 ;
      RECT 8.5 43.6723529412 9.0 43.8823529412 ;
      LAYER M4 ;
      RECT 8.5 43.6723529412 9.0 43.8823529412 ;
      END
    END w_mask_in[40]
  PIN w_mask_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 42.7311764706 9.0 42.9411764706 ;
      LAYER M2 ;
      RECT 8.5 42.7311764706 9.0 42.9411764706 ;
      LAYER M3 ;
      RECT 8.5 42.7311764706 9.0 42.9411764706 ;
      LAYER M4 ;
      RECT 8.5 42.7311764706 9.0 42.9411764706 ;
      END
    END w_mask_in[41]
  PIN w_mask_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 41.79 9.0 42.0 ;
      LAYER M2 ;
      RECT 8.5 41.79 9.0 42.0 ;
      LAYER M3 ;
      RECT 8.5 41.79 9.0 42.0 ;
      LAYER M4 ;
      RECT 8.5 41.79 9.0 42.0 ;
      END
    END w_mask_in[42]
  PIN w_mask_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 40.8488235294 9.0 41.0588235294 ;
      LAYER M2 ;
      RECT 8.5 40.8488235294 9.0 41.0588235294 ;
      LAYER M3 ;
      RECT 8.5 40.8488235294 9.0 41.0588235294 ;
      LAYER M4 ;
      RECT 8.5 40.8488235294 9.0 41.0588235294 ;
      END
    END w_mask_in[43]
  PIN w_mask_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 39.9076470588 9.0 40.1176470588 ;
      LAYER M2 ;
      RECT 8.5 39.9076470588 9.0 40.1176470588 ;
      LAYER M3 ;
      RECT 8.5 39.9076470588 9.0 40.1176470588 ;
      LAYER M4 ;
      RECT 8.5 39.9076470588 9.0 40.1176470588 ;
      END
    END w_mask_in[44]
  PIN w_mask_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 38.9664705882 9.0 39.1764705882 ;
      LAYER M2 ;
      RECT 8.5 38.9664705882 9.0 39.1764705882 ;
      LAYER M3 ;
      RECT 8.5 38.9664705882 9.0 39.1764705882 ;
      LAYER M4 ;
      RECT 8.5 38.9664705882 9.0 39.1764705882 ;
      END
    END w_mask_in[45]
  PIN w_mask_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 38.0252941176 9.0 38.2352941176 ;
      LAYER M2 ;
      RECT 8.5 38.0252941176 9.0 38.2352941176 ;
      LAYER M3 ;
      RECT 8.5 38.0252941176 9.0 38.2352941176 ;
      LAYER M4 ;
      RECT 8.5 38.0252941176 9.0 38.2352941176 ;
      END
    END w_mask_in[46]
  PIN w_mask_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 37.0841176471 9.0 37.2941176471 ;
      LAYER M2 ;
      RECT 8.5 37.0841176471 9.0 37.2941176471 ;
      LAYER M3 ;
      RECT 8.5 37.0841176471 9.0 37.2941176471 ;
      LAYER M4 ;
      RECT 8.5 37.0841176471 9.0 37.2941176471 ;
      END
    END w_mask_in[47]
  PIN w_mask_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 36.1429411765 9.0 36.3529411765 ;
      LAYER M2 ;
      RECT 8.5 36.1429411765 9.0 36.3529411765 ;
      LAYER M3 ;
      RECT 8.5 36.1429411765 9.0 36.3529411765 ;
      LAYER M4 ;
      RECT 8.5 36.1429411765 9.0 36.3529411765 ;
      END
    END w_mask_in[48]
  PIN w_mask_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 35.2017647059 9.0 35.4117647059 ;
      LAYER M2 ;
      RECT 8.5 35.2017647059 9.0 35.4117647059 ;
      LAYER M3 ;
      RECT 8.5 35.2017647059 9.0 35.4117647059 ;
      LAYER M4 ;
      RECT 8.5 35.2017647059 9.0 35.4117647059 ;
      END
    END w_mask_in[49]
  PIN w_mask_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 34.2605882353 9.0 34.4705882353 ;
      LAYER M2 ;
      RECT 8.5 34.2605882353 9.0 34.4705882353 ;
      LAYER M3 ;
      RECT 8.5 34.2605882353 9.0 34.4705882353 ;
      LAYER M4 ;
      RECT 8.5 34.2605882353 9.0 34.4705882353 ;
      END
    END w_mask_in[50]
  PIN w_mask_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 33.3194117647 9.0 33.5294117647 ;
      LAYER M2 ;
      RECT 8.5 33.3194117647 9.0 33.5294117647 ;
      LAYER M3 ;
      RECT 8.5 33.3194117647 9.0 33.5294117647 ;
      LAYER M4 ;
      RECT 8.5 33.3194117647 9.0 33.5294117647 ;
      END
    END w_mask_in[51]
  PIN w_mask_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 32.3782352941 9.0 32.5882352941 ;
      LAYER M2 ;
      RECT 8.5 32.3782352941 9.0 32.5882352941 ;
      LAYER M3 ;
      RECT 8.5 32.3782352941 9.0 32.5882352941 ;
      LAYER M4 ;
      RECT 8.5 32.3782352941 9.0 32.5882352941 ;
      END
    END w_mask_in[52]
  PIN w_mask_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 31.4370588235 9.0 31.6470588235 ;
      LAYER M2 ;
      RECT 8.5 31.4370588235 9.0 31.6470588235 ;
      LAYER M3 ;
      RECT 8.5 31.4370588235 9.0 31.6470588235 ;
      LAYER M4 ;
      RECT 8.5 31.4370588235 9.0 31.6470588235 ;
      END
    END w_mask_in[53]
  PIN w_mask_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 30.4958823529 9.0 30.7058823529 ;
      LAYER M2 ;
      RECT 8.5 30.4958823529 9.0 30.7058823529 ;
      LAYER M3 ;
      RECT 8.5 30.4958823529 9.0 30.7058823529 ;
      LAYER M4 ;
      RECT 8.5 30.4958823529 9.0 30.7058823529 ;
      END
    END w_mask_in[54]
  PIN w_mask_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 29.5547058824 9.0 29.7647058824 ;
      LAYER M2 ;
      RECT 8.5 29.5547058824 9.0 29.7647058824 ;
      LAYER M3 ;
      RECT 8.5 29.5547058824 9.0 29.7647058824 ;
      LAYER M4 ;
      RECT 8.5 29.5547058824 9.0 29.7647058824 ;
      END
    END w_mask_in[55]
  PIN w_mask_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 28.6135294118 9.0 28.8235294118 ;
      LAYER M2 ;
      RECT 8.5 28.6135294118 9.0 28.8235294118 ;
      LAYER M3 ;
      RECT 8.5 28.6135294118 9.0 28.8235294118 ;
      LAYER M4 ;
      RECT 8.5 28.6135294118 9.0 28.8235294118 ;
      END
    END w_mask_in[56]
  PIN w_mask_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 27.6723529412 9.0 27.8823529412 ;
      LAYER M2 ;
      RECT 8.5 27.6723529412 9.0 27.8823529412 ;
      LAYER M3 ;
      RECT 8.5 27.6723529412 9.0 27.8823529412 ;
      LAYER M4 ;
      RECT 8.5 27.6723529412 9.0 27.8823529412 ;
      END
    END w_mask_in[57]
  PIN w_mask_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 26.7311764706 9.0 26.9411764706 ;
      LAYER M2 ;
      RECT 8.5 26.7311764706 9.0 26.9411764706 ;
      LAYER M3 ;
      RECT 8.5 26.7311764706 9.0 26.9411764706 ;
      LAYER M4 ;
      RECT 8.5 26.7311764706 9.0 26.9411764706 ;
      END
    END w_mask_in[58]
  PIN w_mask_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 25.79 9.0 26.0 ;
      LAYER M2 ;
      RECT 8.5 25.79 9.0 26.0 ;
      LAYER M3 ;
      RECT 8.5 25.79 9.0 26.0 ;
      LAYER M4 ;
      RECT 8.5 25.79 9.0 26.0 ;
      END
    END w_mask_in[59]
  PIN w_mask_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 24.8488235294 9.0 25.0588235294 ;
      LAYER M2 ;
      RECT 8.5 24.8488235294 9.0 25.0588235294 ;
      LAYER M3 ;
      RECT 8.5 24.8488235294 9.0 25.0588235294 ;
      LAYER M4 ;
      RECT 8.5 24.8488235294 9.0 25.0588235294 ;
      END
    END w_mask_in[60]
  PIN w_mask_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 23.9076470588 9.0 24.1176470588 ;
      LAYER M2 ;
      RECT 8.5 23.9076470588 9.0 24.1176470588 ;
      LAYER M3 ;
      RECT 8.5 23.9076470588 9.0 24.1176470588 ;
      LAYER M4 ;
      RECT 8.5 23.9076470588 9.0 24.1176470588 ;
      END
    END w_mask_in[61]
  PIN w_mask_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 22.9664705882 9.0 23.1764705882 ;
      LAYER M2 ;
      RECT 8.5 22.9664705882 9.0 23.1764705882 ;
      LAYER M3 ;
      RECT 8.5 22.9664705882 9.0 23.1764705882 ;
      LAYER M4 ;
      RECT 8.5 22.9664705882 9.0 23.1764705882 ;
      END
    END w_mask_in[62]
  PIN w_mask_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 22.0252941176 9.0 22.2352941176 ;
      LAYER M2 ;
      RECT 8.5 22.0252941176 9.0 22.2352941176 ;
      LAYER M3 ;
      RECT 8.5 22.0252941176 9.0 22.2352941176 ;
      LAYER M4 ;
      RECT 8.5 22.0252941176 9.0 22.2352941176 ;
      END
    END w_mask_in[63]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 21.0841176471 9.0 21.2941176471 ;
      LAYER M2 ;
      RECT 8.5 21.0841176471 9.0 21.2941176471 ;
      LAYER M3 ;
      RECT 8.5 21.0841176471 9.0 21.2941176471 ;
      LAYER M4 ;
      RECT 8.5 21.0841176471 9.0 21.2941176471 ;
      END
    END we_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 20.1429411765 9.0 20.3529411765 ;
      LAYER M2 ;
      RECT 8.5 20.1429411765 9.0 20.3529411765 ;
      LAYER M3 ;
      RECT 8.5 20.1429411765 9.0 20.3529411765 ;
      LAYER M4 ;
      RECT 8.5 20.1429411765 9.0 20.3529411765 ;
      END
    END clk
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 8.5 19.2017647059 9.0 19.4117647059 ;
      LAYER M2 ;
      RECT 8.5 19.2017647059 9.0 19.4117647059 ;
      LAYER M3 ;
      RECT 8.5 19.2017647059 9.0 19.4117647059 ;
      LAYER M4 ;
      RECT 8.5 19.2017647059 9.0 19.4117647059 ;
      END
    END ce_in
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 89.5 59.79 90.0 60.0 ;
      LAYER M2 ;
      RECT 89.5 59.79 90.0 60.0 ;
      LAYER M3 ;
      RECT 89.5 59.79 90.0 60.0 ;
      LAYER M4 ;
      RECT 89.5 59.79 90.0 60.0 ;
      END
    END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 88.328125 59.79 88.828125 60.0 ;
      LAYER M2 ;
      RECT 88.328125 59.79 88.828125 60.0 ;
      LAYER M3 ;
      RECT 88.328125 59.79 88.828125 60.0 ;
      LAYER M4 ;
      RECT 88.328125 59.79 88.828125 60.0 ;
      END
    END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 87.15625 59.79 87.65625 60.0 ;
      LAYER M2 ;
      RECT 87.15625 59.79 87.65625 60.0 ;
      LAYER M3 ;
      RECT 87.15625 59.79 87.65625 60.0 ;
      LAYER M4 ;
      RECT 87.15625 59.79 87.65625 60.0 ;
      END
    END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 85.984375 59.79 86.484375 60.0 ;
      LAYER M2 ;
      RECT 85.984375 59.79 86.484375 60.0 ;
      LAYER M3 ;
      RECT 85.984375 59.79 86.484375 60.0 ;
      LAYER M4 ;
      RECT 85.984375 59.79 86.484375 60.0 ;
      END
    END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 84.8125 59.79 85.3125 60.0 ;
      LAYER M2 ;
      RECT 84.8125 59.79 85.3125 60.0 ;
      LAYER M3 ;
      RECT 84.8125 59.79 85.3125 60.0 ;
      LAYER M4 ;
      RECT 84.8125 59.79 85.3125 60.0 ;
      END
    END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 83.640625 59.79 84.140625 60.0 ;
      LAYER M2 ;
      RECT 83.640625 59.79 84.140625 60.0 ;
      LAYER M3 ;
      RECT 83.640625 59.79 84.140625 60.0 ;
      LAYER M4 ;
      RECT 83.640625 59.79 84.140625 60.0 ;
      END
    END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 82.46875 59.79 82.96875 60.0 ;
      LAYER M2 ;
      RECT 82.46875 59.79 82.96875 60.0 ;
      LAYER M3 ;
      RECT 82.46875 59.79 82.96875 60.0 ;
      LAYER M4 ;
      RECT 82.46875 59.79 82.96875 60.0 ;
      END
    END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 81.296875 59.79 81.796875 60.0 ;
      LAYER M2 ;
      RECT 81.296875 59.79 81.796875 60.0 ;
      LAYER M3 ;
      RECT 81.296875 59.79 81.796875 60.0 ;
      LAYER M4 ;
      RECT 81.296875 59.79 81.796875 60.0 ;
      END
    END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 80.125 59.79 80.625 60.0 ;
      LAYER M2 ;
      RECT 80.125 59.79 80.625 60.0 ;
      LAYER M3 ;
      RECT 80.125 59.79 80.625 60.0 ;
      LAYER M4 ;
      RECT 80.125 59.79 80.625 60.0 ;
      END
    END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 78.953125 59.79 79.453125 60.0 ;
      LAYER M2 ;
      RECT 78.953125 59.79 79.453125 60.0 ;
      LAYER M3 ;
      RECT 78.953125 59.79 79.453125 60.0 ;
      LAYER M4 ;
      RECT 78.953125 59.79 79.453125 60.0 ;
      END
    END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 77.78125 59.79 78.28125 60.0 ;
      LAYER M2 ;
      RECT 77.78125 59.79 78.28125 60.0 ;
      LAYER M3 ;
      RECT 77.78125 59.79 78.28125 60.0 ;
      LAYER M4 ;
      RECT 77.78125 59.79 78.28125 60.0 ;
      END
    END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 76.609375 59.79 77.109375 60.0 ;
      LAYER M2 ;
      RECT 76.609375 59.79 77.109375 60.0 ;
      LAYER M3 ;
      RECT 76.609375 59.79 77.109375 60.0 ;
      LAYER M4 ;
      RECT 76.609375 59.79 77.109375 60.0 ;
      END
    END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 75.4375 59.79 75.9375 60.0 ;
      LAYER M2 ;
      RECT 75.4375 59.79 75.9375 60.0 ;
      LAYER M3 ;
      RECT 75.4375 59.79 75.9375 60.0 ;
      LAYER M4 ;
      RECT 75.4375 59.79 75.9375 60.0 ;
      END
    END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 74.265625 59.79 74.765625 60.0 ;
      LAYER M2 ;
      RECT 74.265625 59.79 74.765625 60.0 ;
      LAYER M3 ;
      RECT 74.265625 59.79 74.765625 60.0 ;
      LAYER M4 ;
      RECT 74.265625 59.79 74.765625 60.0 ;
      END
    END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 73.09375 59.79 73.59375 60.0 ;
      LAYER M2 ;
      RECT 73.09375 59.79 73.59375 60.0 ;
      LAYER M3 ;
      RECT 73.09375 59.79 73.59375 60.0 ;
      LAYER M4 ;
      RECT 73.09375 59.79 73.59375 60.0 ;
      END
    END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 71.921875 59.79 72.421875 60.0 ;
      LAYER M2 ;
      RECT 71.921875 59.79 72.421875 60.0 ;
      LAYER M3 ;
      RECT 71.921875 59.79 72.421875 60.0 ;
      LAYER M4 ;
      RECT 71.921875 59.79 72.421875 60.0 ;
      END
    END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 70.75 59.79 71.25 60.0 ;
      LAYER M2 ;
      RECT 70.75 59.79 71.25 60.0 ;
      LAYER M3 ;
      RECT 70.75 59.79 71.25 60.0 ;
      LAYER M4 ;
      RECT 70.75 59.79 71.25 60.0 ;
      END
    END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 69.578125 59.79 70.078125 60.0 ;
      LAYER M2 ;
      RECT 69.578125 59.79 70.078125 60.0 ;
      LAYER M3 ;
      RECT 69.578125 59.79 70.078125 60.0 ;
      LAYER M4 ;
      RECT 69.578125 59.79 70.078125 60.0 ;
      END
    END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 68.40625 59.79 68.90625 60.0 ;
      LAYER M2 ;
      RECT 68.40625 59.79 68.90625 60.0 ;
      LAYER M3 ;
      RECT 68.40625 59.79 68.90625 60.0 ;
      LAYER M4 ;
      RECT 68.40625 59.79 68.90625 60.0 ;
      END
    END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 67.234375 59.79 67.734375 60.0 ;
      LAYER M2 ;
      RECT 67.234375 59.79 67.734375 60.0 ;
      LAYER M3 ;
      RECT 67.234375 59.79 67.734375 60.0 ;
      LAYER M4 ;
      RECT 67.234375 59.79 67.734375 60.0 ;
      END
    END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 66.0625 59.79 66.5625 60.0 ;
      LAYER M2 ;
      RECT 66.0625 59.79 66.5625 60.0 ;
      LAYER M3 ;
      RECT 66.0625 59.79 66.5625 60.0 ;
      LAYER M4 ;
      RECT 66.0625 59.79 66.5625 60.0 ;
      END
    END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 64.890625 59.79 65.390625 60.0 ;
      LAYER M2 ;
      RECT 64.890625 59.79 65.390625 60.0 ;
      LAYER M3 ;
      RECT 64.890625 59.79 65.390625 60.0 ;
      LAYER M4 ;
      RECT 64.890625 59.79 65.390625 60.0 ;
      END
    END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 63.71875 59.79 64.21875 60.0 ;
      LAYER M2 ;
      RECT 63.71875 59.79 64.21875 60.0 ;
      LAYER M3 ;
      RECT 63.71875 59.79 64.21875 60.0 ;
      LAYER M4 ;
      RECT 63.71875 59.79 64.21875 60.0 ;
      END
    END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 62.546875 59.79 63.046875 60.0 ;
      LAYER M2 ;
      RECT 62.546875 59.79 63.046875 60.0 ;
      LAYER M3 ;
      RECT 62.546875 59.79 63.046875 60.0 ;
      LAYER M4 ;
      RECT 62.546875 59.79 63.046875 60.0 ;
      END
    END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 61.375 59.79 61.875 60.0 ;
      LAYER M2 ;
      RECT 61.375 59.79 61.875 60.0 ;
      LAYER M3 ;
      RECT 61.375 59.79 61.875 60.0 ;
      LAYER M4 ;
      RECT 61.375 59.79 61.875 60.0 ;
      END
    END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 60.203125 59.79 60.703125 60.0 ;
      LAYER M2 ;
      RECT 60.203125 59.79 60.703125 60.0 ;
      LAYER M3 ;
      RECT 60.203125 59.79 60.703125 60.0 ;
      LAYER M4 ;
      RECT 60.203125 59.79 60.703125 60.0 ;
      END
    END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 59.03125 59.79 59.53125 60.0 ;
      LAYER M2 ;
      RECT 59.03125 59.79 59.53125 60.0 ;
      LAYER M3 ;
      RECT 59.03125 59.79 59.53125 60.0 ;
      LAYER M4 ;
      RECT 59.03125 59.79 59.53125 60.0 ;
      END
    END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 57.859375 59.79 58.359375 60.0 ;
      LAYER M2 ;
      RECT 57.859375 59.79 58.359375 60.0 ;
      LAYER M3 ;
      RECT 57.859375 59.79 58.359375 60.0 ;
      LAYER M4 ;
      RECT 57.859375 59.79 58.359375 60.0 ;
      END
    END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 56.6875 59.79 57.1875 60.0 ;
      LAYER M2 ;
      RECT 56.6875 59.79 57.1875 60.0 ;
      LAYER M3 ;
      RECT 56.6875 59.79 57.1875 60.0 ;
      LAYER M4 ;
      RECT 56.6875 59.79 57.1875 60.0 ;
      END
    END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 55.515625 59.79 56.015625 60.0 ;
      LAYER M2 ;
      RECT 55.515625 59.79 56.015625 60.0 ;
      LAYER M3 ;
      RECT 55.515625 59.79 56.015625 60.0 ;
      LAYER M4 ;
      RECT 55.515625 59.79 56.015625 60.0 ;
      END
    END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 54.34375 59.79 54.84375 60.0 ;
      LAYER M2 ;
      RECT 54.34375 59.79 54.84375 60.0 ;
      LAYER M3 ;
      RECT 54.34375 59.79 54.84375 60.0 ;
      LAYER M4 ;
      RECT 54.34375 59.79 54.84375 60.0 ;
      END
    END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 53.171875 59.79 53.671875 60.0 ;
      LAYER M2 ;
      RECT 53.171875 59.79 53.671875 60.0 ;
      LAYER M3 ;
      RECT 53.171875 59.79 53.671875 60.0 ;
      LAYER M4 ;
      RECT 53.171875 59.79 53.671875 60.0 ;
      END
    END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 52.0 59.79 52.5 60.0 ;
      LAYER M2 ;
      RECT 52.0 59.79 52.5 60.0 ;
      LAYER M3 ;
      RECT 52.0 59.79 52.5 60.0 ;
      LAYER M4 ;
      RECT 52.0 59.79 52.5 60.0 ;
      END
    END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 50.828125 59.79 51.328125 60.0 ;
      LAYER M2 ;
      RECT 50.828125 59.79 51.328125 60.0 ;
      LAYER M3 ;
      RECT 50.828125 59.79 51.328125 60.0 ;
      LAYER M4 ;
      RECT 50.828125 59.79 51.328125 60.0 ;
      END
    END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 49.65625 59.79 50.15625 60.0 ;
      LAYER M2 ;
      RECT 49.65625 59.79 50.15625 60.0 ;
      LAYER M3 ;
      RECT 49.65625 59.79 50.15625 60.0 ;
      LAYER M4 ;
      RECT 49.65625 59.79 50.15625 60.0 ;
      END
    END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 48.484375 59.79 48.984375 60.0 ;
      LAYER M2 ;
      RECT 48.484375 59.79 48.984375 60.0 ;
      LAYER M3 ;
      RECT 48.484375 59.79 48.984375 60.0 ;
      LAYER M4 ;
      RECT 48.484375 59.79 48.984375 60.0 ;
      END
    END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 47.3125 59.79 47.8125 60.0 ;
      LAYER M2 ;
      RECT 47.3125 59.79 47.8125 60.0 ;
      LAYER M3 ;
      RECT 47.3125 59.79 47.8125 60.0 ;
      LAYER M4 ;
      RECT 47.3125 59.79 47.8125 60.0 ;
      END
    END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 46.140625 59.79 46.640625 60.0 ;
      LAYER M2 ;
      RECT 46.140625 59.79 46.640625 60.0 ;
      LAYER M3 ;
      RECT 46.140625 59.79 46.640625 60.0 ;
      LAYER M4 ;
      RECT 46.140625 59.79 46.640625 60.0 ;
      END
    END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 44.96875 59.79 45.46875 60.0 ;
      LAYER M2 ;
      RECT 44.96875 59.79 45.46875 60.0 ;
      LAYER M3 ;
      RECT 44.96875 59.79 45.46875 60.0 ;
      LAYER M4 ;
      RECT 44.96875 59.79 45.46875 60.0 ;
      END
    END rd_out[38]
  PIN rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 43.796875 59.79 44.296875 60.0 ;
      LAYER M2 ;
      RECT 43.796875 59.79 44.296875 60.0 ;
      LAYER M3 ;
      RECT 43.796875 59.79 44.296875 60.0 ;
      LAYER M4 ;
      RECT 43.796875 59.79 44.296875 60.0 ;
      END
    END rd_out[39]
  PIN rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 42.625 59.79 43.125 60.0 ;
      LAYER M2 ;
      RECT 42.625 59.79 43.125 60.0 ;
      LAYER M3 ;
      RECT 42.625 59.79 43.125 60.0 ;
      LAYER M4 ;
      RECT 42.625 59.79 43.125 60.0 ;
      END
    END rd_out[40]
  PIN rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 41.453125 59.79 41.953125 60.0 ;
      LAYER M2 ;
      RECT 41.453125 59.79 41.953125 60.0 ;
      LAYER M3 ;
      RECT 41.453125 59.79 41.953125 60.0 ;
      LAYER M4 ;
      RECT 41.453125 59.79 41.953125 60.0 ;
      END
    END rd_out[41]
  PIN rd_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 40.28125 59.79 40.78125 60.0 ;
      LAYER M2 ;
      RECT 40.28125 59.79 40.78125 60.0 ;
      LAYER M3 ;
      RECT 40.28125 59.79 40.78125 60.0 ;
      LAYER M4 ;
      RECT 40.28125 59.79 40.78125 60.0 ;
      END
    END rd_out[42]
  PIN rd_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 39.109375 59.79 39.609375 60.0 ;
      LAYER M2 ;
      RECT 39.109375 59.79 39.609375 60.0 ;
      LAYER M3 ;
      RECT 39.109375 59.79 39.609375 60.0 ;
      LAYER M4 ;
      RECT 39.109375 59.79 39.609375 60.0 ;
      END
    END rd_out[43]
  PIN rd_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 37.9375 59.79 38.4375 60.0 ;
      LAYER M2 ;
      RECT 37.9375 59.79 38.4375 60.0 ;
      LAYER M3 ;
      RECT 37.9375 59.79 38.4375 60.0 ;
      LAYER M4 ;
      RECT 37.9375 59.79 38.4375 60.0 ;
      END
    END rd_out[44]
  PIN rd_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 36.765625 59.79 37.265625 60.0 ;
      LAYER M2 ;
      RECT 36.765625 59.79 37.265625 60.0 ;
      LAYER M3 ;
      RECT 36.765625 59.79 37.265625 60.0 ;
      LAYER M4 ;
      RECT 36.765625 59.79 37.265625 60.0 ;
      END
    END rd_out[45]
  PIN rd_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 35.59375 59.79 36.09375 60.0 ;
      LAYER M2 ;
      RECT 35.59375 59.79 36.09375 60.0 ;
      LAYER M3 ;
      RECT 35.59375 59.79 36.09375 60.0 ;
      LAYER M4 ;
      RECT 35.59375 59.79 36.09375 60.0 ;
      END
    END rd_out[46]
  PIN rd_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 34.421875 59.79 34.921875 60.0 ;
      LAYER M2 ;
      RECT 34.421875 59.79 34.921875 60.0 ;
      LAYER M3 ;
      RECT 34.421875 59.79 34.921875 60.0 ;
      LAYER M4 ;
      RECT 34.421875 59.79 34.921875 60.0 ;
      END
    END rd_out[47]
  PIN rd_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 33.25 59.79 33.75 60.0 ;
      LAYER M2 ;
      RECT 33.25 59.79 33.75 60.0 ;
      LAYER M3 ;
      RECT 33.25 59.79 33.75 60.0 ;
      LAYER M4 ;
      RECT 33.25 59.79 33.75 60.0 ;
      END
    END rd_out[48]
  PIN rd_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 32.078125 59.79 32.578125 60.0 ;
      LAYER M2 ;
      RECT 32.078125 59.79 32.578125 60.0 ;
      LAYER M3 ;
      RECT 32.078125 59.79 32.578125 60.0 ;
      LAYER M4 ;
      RECT 32.078125 59.79 32.578125 60.0 ;
      END
    END rd_out[49]
  PIN rd_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 30.90625 59.79 31.40625 60.0 ;
      LAYER M2 ;
      RECT 30.90625 59.79 31.40625 60.0 ;
      LAYER M3 ;
      RECT 30.90625 59.79 31.40625 60.0 ;
      LAYER M4 ;
      RECT 30.90625 59.79 31.40625 60.0 ;
      END
    END rd_out[50]
  PIN rd_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 29.734375 59.79 30.234375 60.0 ;
      LAYER M2 ;
      RECT 29.734375 59.79 30.234375 60.0 ;
      LAYER M3 ;
      RECT 29.734375 59.79 30.234375 60.0 ;
      LAYER M4 ;
      RECT 29.734375 59.79 30.234375 60.0 ;
      END
    END rd_out[51]
  PIN rd_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 28.5625 59.79 29.0625 60.0 ;
      LAYER M2 ;
      RECT 28.5625 59.79 29.0625 60.0 ;
      LAYER M3 ;
      RECT 28.5625 59.79 29.0625 60.0 ;
      LAYER M4 ;
      RECT 28.5625 59.79 29.0625 60.0 ;
      END
    END rd_out[52]
  PIN rd_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 27.390625 59.79 27.890625 60.0 ;
      LAYER M2 ;
      RECT 27.390625 59.79 27.890625 60.0 ;
      LAYER M3 ;
      RECT 27.390625 59.79 27.890625 60.0 ;
      LAYER M4 ;
      RECT 27.390625 59.79 27.890625 60.0 ;
      END
    END rd_out[53]
  PIN rd_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 26.21875 59.79 26.71875 60.0 ;
      LAYER M2 ;
      RECT 26.21875 59.79 26.71875 60.0 ;
      LAYER M3 ;
      RECT 26.21875 59.79 26.71875 60.0 ;
      LAYER M4 ;
      RECT 26.21875 59.79 26.71875 60.0 ;
      END
    END rd_out[54]
  PIN rd_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 25.046875 59.79 25.546875 60.0 ;
      LAYER M2 ;
      RECT 25.046875 59.79 25.546875 60.0 ;
      LAYER M3 ;
      RECT 25.046875 59.79 25.546875 60.0 ;
      LAYER M4 ;
      RECT 25.046875 59.79 25.546875 60.0 ;
      END
    END rd_out[55]
  PIN rd_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 23.875 59.79 24.375 60.0 ;
      LAYER M2 ;
      RECT 23.875 59.79 24.375 60.0 ;
      LAYER M3 ;
      RECT 23.875 59.79 24.375 60.0 ;
      LAYER M4 ;
      RECT 23.875 59.79 24.375 60.0 ;
      END
    END rd_out[56]
  PIN rd_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 22.703125 59.79 23.203125 60.0 ;
      LAYER M2 ;
      RECT 22.703125 59.79 23.203125 60.0 ;
      LAYER M3 ;
      RECT 22.703125 59.79 23.203125 60.0 ;
      LAYER M4 ;
      RECT 22.703125 59.79 23.203125 60.0 ;
      END
    END rd_out[57]
  PIN rd_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 21.53125 59.79 22.03125 60.0 ;
      LAYER M2 ;
      RECT 21.53125 59.79 22.03125 60.0 ;
      LAYER M3 ;
      RECT 21.53125 59.79 22.03125 60.0 ;
      LAYER M4 ;
      RECT 21.53125 59.79 22.03125 60.0 ;
      END
    END rd_out[58]
  PIN rd_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 20.359375 59.79 20.859375 60.0 ;
      LAYER M2 ;
      RECT 20.359375 59.79 20.859375 60.0 ;
      LAYER M3 ;
      RECT 20.359375 59.79 20.859375 60.0 ;
      LAYER M4 ;
      RECT 20.359375 59.79 20.859375 60.0 ;
      END
    END rd_out[59]
  PIN rd_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 19.1875 59.79 19.6875 60.0 ;
      LAYER M2 ;
      RECT 19.1875 59.79 19.6875 60.0 ;
      LAYER M3 ;
      RECT 19.1875 59.79 19.6875 60.0 ;
      LAYER M4 ;
      RECT 19.1875 59.79 19.6875 60.0 ;
      END
    END rd_out[60]
  PIN rd_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 18.015625 59.79 18.515625 60.0 ;
      LAYER M2 ;
      RECT 18.015625 59.79 18.515625 60.0 ;
      LAYER M3 ;
      RECT 18.015625 59.79 18.515625 60.0 ;
      LAYER M4 ;
      RECT 18.015625 59.79 18.515625 60.0 ;
      END
    END rd_out[61]
  PIN rd_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 16.84375 59.79 17.34375 60.0 ;
      LAYER M2 ;
      RECT 16.84375 59.79 17.34375 60.0 ;
      LAYER M3 ;
      RECT 16.84375 59.79 17.34375 60.0 ;
      LAYER M4 ;
      RECT 16.84375 59.79 17.34375 60.0 ;
      END
    END rd_out[62]
  PIN rd_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 15.671875 59.79 16.171875 60.0 ;
      LAYER M2 ;
      RECT 15.671875 59.79 16.171875 60.0 ;
      LAYER M3 ;
      RECT 15.671875 59.79 16.171875 60.0 ;
      LAYER M4 ;
      RECT 15.671875 59.79 16.171875 60.0 ;
      END
    END rd_out[63]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 89.5 39.79 90.0 40.0 ;
      LAYER M2 ;
      RECT 89.5 39.79 90.0 40.0 ;
      LAYER M3 ;
      RECT 89.5 39.79 90.0 40.0 ;
      LAYER M4 ;
      RECT 89.5 39.79 90.0 40.0 ;
      END
    END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 88.328125 39.79 88.828125 40.0 ;
      LAYER M2 ;
      RECT 88.328125 39.79 88.828125 40.0 ;
      LAYER M3 ;
      RECT 88.328125 39.79 88.828125 40.0 ;
      LAYER M4 ;
      RECT 88.328125 39.79 88.828125 40.0 ;
      END
    END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 87.15625 39.79 87.65625 40.0 ;
      LAYER M2 ;
      RECT 87.15625 39.79 87.65625 40.0 ;
      LAYER M3 ;
      RECT 87.15625 39.79 87.65625 40.0 ;
      LAYER M4 ;
      RECT 87.15625 39.79 87.65625 40.0 ;
      END
    END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 85.984375 39.79 86.484375 40.0 ;
      LAYER M2 ;
      RECT 85.984375 39.79 86.484375 40.0 ;
      LAYER M3 ;
      RECT 85.984375 39.79 86.484375 40.0 ;
      LAYER M4 ;
      RECT 85.984375 39.79 86.484375 40.0 ;
      END
    END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 84.8125 39.79 85.3125 40.0 ;
      LAYER M2 ;
      RECT 84.8125 39.79 85.3125 40.0 ;
      LAYER M3 ;
      RECT 84.8125 39.79 85.3125 40.0 ;
      LAYER M4 ;
      RECT 84.8125 39.79 85.3125 40.0 ;
      END
    END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 83.640625 39.79 84.140625 40.0 ;
      LAYER M2 ;
      RECT 83.640625 39.79 84.140625 40.0 ;
      LAYER M3 ;
      RECT 83.640625 39.79 84.140625 40.0 ;
      LAYER M4 ;
      RECT 83.640625 39.79 84.140625 40.0 ;
      END
    END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 82.46875 39.79 82.96875 40.0 ;
      LAYER M2 ;
      RECT 82.46875 39.79 82.96875 40.0 ;
      LAYER M3 ;
      RECT 82.46875 39.79 82.96875 40.0 ;
      LAYER M4 ;
      RECT 82.46875 39.79 82.96875 40.0 ;
      END
    END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 81.296875 39.79 81.796875 40.0 ;
      LAYER M2 ;
      RECT 81.296875 39.79 81.796875 40.0 ;
      LAYER M3 ;
      RECT 81.296875 39.79 81.796875 40.0 ;
      LAYER M4 ;
      RECT 81.296875 39.79 81.796875 40.0 ;
      END
    END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 80.125 39.79 80.625 40.0 ;
      LAYER M2 ;
      RECT 80.125 39.79 80.625 40.0 ;
      LAYER M3 ;
      RECT 80.125 39.79 80.625 40.0 ;
      LAYER M4 ;
      RECT 80.125 39.79 80.625 40.0 ;
      END
    END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 78.953125 39.79 79.453125 40.0 ;
      LAYER M2 ;
      RECT 78.953125 39.79 79.453125 40.0 ;
      LAYER M3 ;
      RECT 78.953125 39.79 79.453125 40.0 ;
      LAYER M4 ;
      RECT 78.953125 39.79 79.453125 40.0 ;
      END
    END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 77.78125 39.79 78.28125 40.0 ;
      LAYER M2 ;
      RECT 77.78125 39.79 78.28125 40.0 ;
      LAYER M3 ;
      RECT 77.78125 39.79 78.28125 40.0 ;
      LAYER M4 ;
      RECT 77.78125 39.79 78.28125 40.0 ;
      END
    END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 76.609375 39.79 77.109375 40.0 ;
      LAYER M2 ;
      RECT 76.609375 39.79 77.109375 40.0 ;
      LAYER M3 ;
      RECT 76.609375 39.79 77.109375 40.0 ;
      LAYER M4 ;
      RECT 76.609375 39.79 77.109375 40.0 ;
      END
    END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 75.4375 39.79 75.9375 40.0 ;
      LAYER M2 ;
      RECT 75.4375 39.79 75.9375 40.0 ;
      LAYER M3 ;
      RECT 75.4375 39.79 75.9375 40.0 ;
      LAYER M4 ;
      RECT 75.4375 39.79 75.9375 40.0 ;
      END
    END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 74.265625 39.79 74.765625 40.0 ;
      LAYER M2 ;
      RECT 74.265625 39.79 74.765625 40.0 ;
      LAYER M3 ;
      RECT 74.265625 39.79 74.765625 40.0 ;
      LAYER M4 ;
      RECT 74.265625 39.79 74.765625 40.0 ;
      END
    END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 73.09375 39.79 73.59375 40.0 ;
      LAYER M2 ;
      RECT 73.09375 39.79 73.59375 40.0 ;
      LAYER M3 ;
      RECT 73.09375 39.79 73.59375 40.0 ;
      LAYER M4 ;
      RECT 73.09375 39.79 73.59375 40.0 ;
      END
    END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 71.921875 39.79 72.421875 40.0 ;
      LAYER M2 ;
      RECT 71.921875 39.79 72.421875 40.0 ;
      LAYER M3 ;
      RECT 71.921875 39.79 72.421875 40.0 ;
      LAYER M4 ;
      RECT 71.921875 39.79 72.421875 40.0 ;
      END
    END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 70.75 39.79 71.25 40.0 ;
      LAYER M2 ;
      RECT 70.75 39.79 71.25 40.0 ;
      LAYER M3 ;
      RECT 70.75 39.79 71.25 40.0 ;
      LAYER M4 ;
      RECT 70.75 39.79 71.25 40.0 ;
      END
    END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 69.578125 39.79 70.078125 40.0 ;
      LAYER M2 ;
      RECT 69.578125 39.79 70.078125 40.0 ;
      LAYER M3 ;
      RECT 69.578125 39.79 70.078125 40.0 ;
      LAYER M4 ;
      RECT 69.578125 39.79 70.078125 40.0 ;
      END
    END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 68.40625 39.79 68.90625 40.0 ;
      LAYER M2 ;
      RECT 68.40625 39.79 68.90625 40.0 ;
      LAYER M3 ;
      RECT 68.40625 39.79 68.90625 40.0 ;
      LAYER M4 ;
      RECT 68.40625 39.79 68.90625 40.0 ;
      END
    END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 67.234375 39.79 67.734375 40.0 ;
      LAYER M2 ;
      RECT 67.234375 39.79 67.734375 40.0 ;
      LAYER M3 ;
      RECT 67.234375 39.79 67.734375 40.0 ;
      LAYER M4 ;
      RECT 67.234375 39.79 67.734375 40.0 ;
      END
    END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 66.0625 39.79 66.5625 40.0 ;
      LAYER M2 ;
      RECT 66.0625 39.79 66.5625 40.0 ;
      LAYER M3 ;
      RECT 66.0625 39.79 66.5625 40.0 ;
      LAYER M4 ;
      RECT 66.0625 39.79 66.5625 40.0 ;
      END
    END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 64.890625 39.79 65.390625 40.0 ;
      LAYER M2 ;
      RECT 64.890625 39.79 65.390625 40.0 ;
      LAYER M3 ;
      RECT 64.890625 39.79 65.390625 40.0 ;
      LAYER M4 ;
      RECT 64.890625 39.79 65.390625 40.0 ;
      END
    END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 63.71875 39.79 64.21875 40.0 ;
      LAYER M2 ;
      RECT 63.71875 39.79 64.21875 40.0 ;
      LAYER M3 ;
      RECT 63.71875 39.79 64.21875 40.0 ;
      LAYER M4 ;
      RECT 63.71875 39.79 64.21875 40.0 ;
      END
    END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 62.546875 39.79 63.046875 40.0 ;
      LAYER M2 ;
      RECT 62.546875 39.79 63.046875 40.0 ;
      LAYER M3 ;
      RECT 62.546875 39.79 63.046875 40.0 ;
      LAYER M4 ;
      RECT 62.546875 39.79 63.046875 40.0 ;
      END
    END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 61.375 39.79 61.875 40.0 ;
      LAYER M2 ;
      RECT 61.375 39.79 61.875 40.0 ;
      LAYER M3 ;
      RECT 61.375 39.79 61.875 40.0 ;
      LAYER M4 ;
      RECT 61.375 39.79 61.875 40.0 ;
      END
    END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 60.203125 39.79 60.703125 40.0 ;
      LAYER M2 ;
      RECT 60.203125 39.79 60.703125 40.0 ;
      LAYER M3 ;
      RECT 60.203125 39.79 60.703125 40.0 ;
      LAYER M4 ;
      RECT 60.203125 39.79 60.703125 40.0 ;
      END
    END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 59.03125 39.79 59.53125 40.0 ;
      LAYER M2 ;
      RECT 59.03125 39.79 59.53125 40.0 ;
      LAYER M3 ;
      RECT 59.03125 39.79 59.53125 40.0 ;
      LAYER M4 ;
      RECT 59.03125 39.79 59.53125 40.0 ;
      END
    END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 57.859375 39.79 58.359375 40.0 ;
      LAYER M2 ;
      RECT 57.859375 39.79 58.359375 40.0 ;
      LAYER M3 ;
      RECT 57.859375 39.79 58.359375 40.0 ;
      LAYER M4 ;
      RECT 57.859375 39.79 58.359375 40.0 ;
      END
    END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 56.6875 39.79 57.1875 40.0 ;
      LAYER M2 ;
      RECT 56.6875 39.79 57.1875 40.0 ;
      LAYER M3 ;
      RECT 56.6875 39.79 57.1875 40.0 ;
      LAYER M4 ;
      RECT 56.6875 39.79 57.1875 40.0 ;
      END
    END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 55.515625 39.79 56.015625 40.0 ;
      LAYER M2 ;
      RECT 55.515625 39.79 56.015625 40.0 ;
      LAYER M3 ;
      RECT 55.515625 39.79 56.015625 40.0 ;
      LAYER M4 ;
      RECT 55.515625 39.79 56.015625 40.0 ;
      END
    END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 54.34375 39.79 54.84375 40.0 ;
      LAYER M2 ;
      RECT 54.34375 39.79 54.84375 40.0 ;
      LAYER M3 ;
      RECT 54.34375 39.79 54.84375 40.0 ;
      LAYER M4 ;
      RECT 54.34375 39.79 54.84375 40.0 ;
      END
    END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 53.171875 39.79 53.671875 40.0 ;
      LAYER M2 ;
      RECT 53.171875 39.79 53.671875 40.0 ;
      LAYER M3 ;
      RECT 53.171875 39.79 53.671875 40.0 ;
      LAYER M4 ;
      RECT 53.171875 39.79 53.671875 40.0 ;
      END
    END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 52.0 39.79 52.5 40.0 ;
      LAYER M2 ;
      RECT 52.0 39.79 52.5 40.0 ;
      LAYER M3 ;
      RECT 52.0 39.79 52.5 40.0 ;
      LAYER M4 ;
      RECT 52.0 39.79 52.5 40.0 ;
      END
    END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 50.828125 39.79 51.328125 40.0 ;
      LAYER M2 ;
      RECT 50.828125 39.79 51.328125 40.0 ;
      LAYER M3 ;
      RECT 50.828125 39.79 51.328125 40.0 ;
      LAYER M4 ;
      RECT 50.828125 39.79 51.328125 40.0 ;
      END
    END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 49.65625 39.79 50.15625 40.0 ;
      LAYER M2 ;
      RECT 49.65625 39.79 50.15625 40.0 ;
      LAYER M3 ;
      RECT 49.65625 39.79 50.15625 40.0 ;
      LAYER M4 ;
      RECT 49.65625 39.79 50.15625 40.0 ;
      END
    END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 48.484375 39.79 48.984375 40.0 ;
      LAYER M2 ;
      RECT 48.484375 39.79 48.984375 40.0 ;
      LAYER M3 ;
      RECT 48.484375 39.79 48.984375 40.0 ;
      LAYER M4 ;
      RECT 48.484375 39.79 48.984375 40.0 ;
      END
    END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 47.3125 39.79 47.8125 40.0 ;
      LAYER M2 ;
      RECT 47.3125 39.79 47.8125 40.0 ;
      LAYER M3 ;
      RECT 47.3125 39.79 47.8125 40.0 ;
      LAYER M4 ;
      RECT 47.3125 39.79 47.8125 40.0 ;
      END
    END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 46.140625 39.79 46.640625 40.0 ;
      LAYER M2 ;
      RECT 46.140625 39.79 46.640625 40.0 ;
      LAYER M3 ;
      RECT 46.140625 39.79 46.640625 40.0 ;
      LAYER M4 ;
      RECT 46.140625 39.79 46.640625 40.0 ;
      END
    END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 44.96875 39.79 45.46875 40.0 ;
      LAYER M2 ;
      RECT 44.96875 39.79 45.46875 40.0 ;
      LAYER M3 ;
      RECT 44.96875 39.79 45.46875 40.0 ;
      LAYER M4 ;
      RECT 44.96875 39.79 45.46875 40.0 ;
      END
    END wd_in[38]
  PIN wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 43.796875 39.79 44.296875 40.0 ;
      LAYER M2 ;
      RECT 43.796875 39.79 44.296875 40.0 ;
      LAYER M3 ;
      RECT 43.796875 39.79 44.296875 40.0 ;
      LAYER M4 ;
      RECT 43.796875 39.79 44.296875 40.0 ;
      END
    END wd_in[39]
  PIN wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 42.625 39.79 43.125 40.0 ;
      LAYER M2 ;
      RECT 42.625 39.79 43.125 40.0 ;
      LAYER M3 ;
      RECT 42.625 39.79 43.125 40.0 ;
      LAYER M4 ;
      RECT 42.625 39.79 43.125 40.0 ;
      END
    END wd_in[40]
  PIN wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 41.453125 39.79 41.953125 40.0 ;
      LAYER M2 ;
      RECT 41.453125 39.79 41.953125 40.0 ;
      LAYER M3 ;
      RECT 41.453125 39.79 41.953125 40.0 ;
      LAYER M4 ;
      RECT 41.453125 39.79 41.953125 40.0 ;
      END
    END wd_in[41]
  PIN wd_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 40.28125 39.79 40.78125 40.0 ;
      LAYER M2 ;
      RECT 40.28125 39.79 40.78125 40.0 ;
      LAYER M3 ;
      RECT 40.28125 39.79 40.78125 40.0 ;
      LAYER M4 ;
      RECT 40.28125 39.79 40.78125 40.0 ;
      END
    END wd_in[42]
  PIN wd_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 39.109375 39.79 39.609375 40.0 ;
      LAYER M2 ;
      RECT 39.109375 39.79 39.609375 40.0 ;
      LAYER M3 ;
      RECT 39.109375 39.79 39.609375 40.0 ;
      LAYER M4 ;
      RECT 39.109375 39.79 39.609375 40.0 ;
      END
    END wd_in[43]
  PIN wd_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 37.9375 39.79 38.4375 40.0 ;
      LAYER M2 ;
      RECT 37.9375 39.79 38.4375 40.0 ;
      LAYER M3 ;
      RECT 37.9375 39.79 38.4375 40.0 ;
      LAYER M4 ;
      RECT 37.9375 39.79 38.4375 40.0 ;
      END
    END wd_in[44]
  PIN wd_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 36.765625 39.79 37.265625 40.0 ;
      LAYER M2 ;
      RECT 36.765625 39.79 37.265625 40.0 ;
      LAYER M3 ;
      RECT 36.765625 39.79 37.265625 40.0 ;
      LAYER M4 ;
      RECT 36.765625 39.79 37.265625 40.0 ;
      END
    END wd_in[45]
  PIN wd_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 35.59375 39.79 36.09375 40.0 ;
      LAYER M2 ;
      RECT 35.59375 39.79 36.09375 40.0 ;
      LAYER M3 ;
      RECT 35.59375 39.79 36.09375 40.0 ;
      LAYER M4 ;
      RECT 35.59375 39.79 36.09375 40.0 ;
      END
    END wd_in[46]
  PIN wd_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 34.421875 39.79 34.921875 40.0 ;
      LAYER M2 ;
      RECT 34.421875 39.79 34.921875 40.0 ;
      LAYER M3 ;
      RECT 34.421875 39.79 34.921875 40.0 ;
      LAYER M4 ;
      RECT 34.421875 39.79 34.921875 40.0 ;
      END
    END wd_in[47]
  PIN wd_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 33.25 39.79 33.75 40.0 ;
      LAYER M2 ;
      RECT 33.25 39.79 33.75 40.0 ;
      LAYER M3 ;
      RECT 33.25 39.79 33.75 40.0 ;
      LAYER M4 ;
      RECT 33.25 39.79 33.75 40.0 ;
      END
    END wd_in[48]
  PIN wd_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 32.078125 39.79 32.578125 40.0 ;
      LAYER M2 ;
      RECT 32.078125 39.79 32.578125 40.0 ;
      LAYER M3 ;
      RECT 32.078125 39.79 32.578125 40.0 ;
      LAYER M4 ;
      RECT 32.078125 39.79 32.578125 40.0 ;
      END
    END wd_in[49]
  PIN wd_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 30.90625 39.79 31.40625 40.0 ;
      LAYER M2 ;
      RECT 30.90625 39.79 31.40625 40.0 ;
      LAYER M3 ;
      RECT 30.90625 39.79 31.40625 40.0 ;
      LAYER M4 ;
      RECT 30.90625 39.79 31.40625 40.0 ;
      END
    END wd_in[50]
  PIN wd_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 29.734375 39.79 30.234375 40.0 ;
      LAYER M2 ;
      RECT 29.734375 39.79 30.234375 40.0 ;
      LAYER M3 ;
      RECT 29.734375 39.79 30.234375 40.0 ;
      LAYER M4 ;
      RECT 29.734375 39.79 30.234375 40.0 ;
      END
    END wd_in[51]
  PIN wd_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 28.5625 39.79 29.0625 40.0 ;
      LAYER M2 ;
      RECT 28.5625 39.79 29.0625 40.0 ;
      LAYER M3 ;
      RECT 28.5625 39.79 29.0625 40.0 ;
      LAYER M4 ;
      RECT 28.5625 39.79 29.0625 40.0 ;
      END
    END wd_in[52]
  PIN wd_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 27.390625 39.79 27.890625 40.0 ;
      LAYER M2 ;
      RECT 27.390625 39.79 27.890625 40.0 ;
      LAYER M3 ;
      RECT 27.390625 39.79 27.890625 40.0 ;
      LAYER M4 ;
      RECT 27.390625 39.79 27.890625 40.0 ;
      END
    END wd_in[53]
  PIN wd_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 26.21875 39.79 26.71875 40.0 ;
      LAYER M2 ;
      RECT 26.21875 39.79 26.71875 40.0 ;
      LAYER M3 ;
      RECT 26.21875 39.79 26.71875 40.0 ;
      LAYER M4 ;
      RECT 26.21875 39.79 26.71875 40.0 ;
      END
    END wd_in[54]
  PIN wd_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 25.046875 39.79 25.546875 40.0 ;
      LAYER M2 ;
      RECT 25.046875 39.79 25.546875 40.0 ;
      LAYER M3 ;
      RECT 25.046875 39.79 25.546875 40.0 ;
      LAYER M4 ;
      RECT 25.046875 39.79 25.546875 40.0 ;
      END
    END wd_in[55]
  PIN wd_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 23.875 39.79 24.375 40.0 ;
      LAYER M2 ;
      RECT 23.875 39.79 24.375 40.0 ;
      LAYER M3 ;
      RECT 23.875 39.79 24.375 40.0 ;
      LAYER M4 ;
      RECT 23.875 39.79 24.375 40.0 ;
      END
    END wd_in[56]
  PIN wd_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 22.703125 39.79 23.203125 40.0 ;
      LAYER M2 ;
      RECT 22.703125 39.79 23.203125 40.0 ;
      LAYER M3 ;
      RECT 22.703125 39.79 23.203125 40.0 ;
      LAYER M4 ;
      RECT 22.703125 39.79 23.203125 40.0 ;
      END
    END wd_in[57]
  PIN wd_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 21.53125 39.79 22.03125 40.0 ;
      LAYER M2 ;
      RECT 21.53125 39.79 22.03125 40.0 ;
      LAYER M3 ;
      RECT 21.53125 39.79 22.03125 40.0 ;
      LAYER M4 ;
      RECT 21.53125 39.79 22.03125 40.0 ;
      END
    END wd_in[58]
  PIN wd_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 20.359375 39.79 20.859375 40.0 ;
      LAYER M2 ;
      RECT 20.359375 39.79 20.859375 40.0 ;
      LAYER M3 ;
      RECT 20.359375 39.79 20.859375 40.0 ;
      LAYER M4 ;
      RECT 20.359375 39.79 20.859375 40.0 ;
      END
    END wd_in[59]
  PIN wd_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 19.1875 39.79 19.6875 40.0 ;
      LAYER M2 ;
      RECT 19.1875 39.79 19.6875 40.0 ;
      LAYER M3 ;
      RECT 19.1875 39.79 19.6875 40.0 ;
      LAYER M4 ;
      RECT 19.1875 39.79 19.6875 40.0 ;
      END
    END wd_in[60]
  PIN wd_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 18.015625 39.79 18.515625 40.0 ;
      LAYER M2 ;
      RECT 18.015625 39.79 18.515625 40.0 ;
      LAYER M3 ;
      RECT 18.015625 39.79 18.515625 40.0 ;
      LAYER M4 ;
      RECT 18.015625 39.79 18.515625 40.0 ;
      END
    END wd_in[61]
  PIN wd_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 16.84375 39.79 17.34375 40.0 ;
      LAYER M2 ;
      RECT 16.84375 39.79 17.34375 40.0 ;
      LAYER M3 ;
      RECT 16.84375 39.79 17.34375 40.0 ;
      LAYER M4 ;
      RECT 16.84375 39.79 17.34375 40.0 ;
      END
    END wd_in[62]
  PIN wd_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 15.671875 39.79 16.171875 40.0 ;
      LAYER M2 ;
      RECT 15.671875 39.79 16.171875 40.0 ;
      LAYER M3 ;
      RECT 15.671875 39.79 16.171875 40.0 ;
      LAYER M4 ;
      RECT 15.671875 39.79 16.171875 40.0 ;
      END
    END wd_in[63]
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE RING ;
    PORT
      LAYER M3 ;
      RECT 3.5 3.5 5.5 96.5 ;
      END
    PORT
      LAYER M4 ;
      RECT 3.5 3.5 5.5 96.5 ;
      END
    END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE RING ;
    PORT
      LAYER M3 ;
      RECT 0.0 0.0 98.0 2.0 ;
      END
    PORT
      LAYER M4 ;
      RECT 0.0 0.0 98.0 2.0 ;
      END
    END VDD
  OBS
    #core
    LAYER VIA1 ;
    RECT 8.5 8.5 91.5 91.5 ;
    LAYER VIA2 ;
    RECT 8.5 8.5 91.5 91.5 ;
    LAYER VIA3 ;
    RECT 8.5 8.5 91.5 91.5 ;
    LAYER OVERLAP ;
    RECT 8.5 8.5 91.5 91.5 ;
    END
  END nangate45_64x512_1P_BM

END LIBRARY
